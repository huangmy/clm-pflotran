netcdf ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "fractional area burned" ;
		FAREA_BURNED:units = "proportion/sec" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 09/25/14 13:24:15" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:natpft_not_vegetated = 1 ;
		:natpft_needleleaf_evergreen_temperate_tree = 2 ;
		:natpft_needleleaf_evergreen_boreal_tree = 3 ;
		:natpft_needleleaf_deciduous_boreal_tree = 4 ;
		:natpft_broadleaf_evergreen_tropical_tree = 5 ;
		:natpft_broadleaf_evergreen_temperate_tree = 6 ;
		:natpft_broadleaf_deciduous_tropical_tree = 7 ;
		:natpft_broadleaf_deciduous_temperate_tree = 8 ;
		:natpft_broadleaf_deciduous_boreal_tree = 9 ;
		:natpft_broadleaf_evergreen_shrub = 10 ;
		:natpft_broadleaf_deciduous_temperate_shrub = 11 ;
		:natpft_broadleaf_deciduous_boreal_shrub = 12 ;
		:natpft_c3_arctic_grass = 13 ;
		:natpft_c3_non-arctic_grass = 14 ;
		:natpft_c4_grass = 15 ;
		:natpft_c3_crop = 16 ;
		:natpft_c3_irrigated = 17 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "09/25/14" ;

 time_written =
  "13:24:15" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.044949e-14, 5.058576e-14, 5.055929e-14, 5.066909e-14, 5.060821e-14, 
    5.068008e-14, 5.047715e-14, 5.059115e-14, 5.051839e-14, 5.046179e-14, 
    5.088186e-14, 5.067399e-14, 5.109757e-14, 5.096525e-14, 5.129742e-14, 
    5.107696e-14, 5.134183e-14, 5.129111e-14, 5.144381e-14, 5.140008e-14, 
    5.159509e-14, 5.146398e-14, 5.169611e-14, 5.156382e-14, 5.158451e-14, 
    5.145965e-14, 5.071589e-14, 5.085598e-14, 5.070758e-14, 5.072757e-14, 
    5.07186e-14, 5.060945e-14, 5.055439e-14, 5.04391e-14, 5.046004e-14, 
    5.054473e-14, 5.073656e-14, 5.06715e-14, 5.083547e-14, 5.083177e-14, 
    5.101405e-14, 5.093189e-14, 5.123788e-14, 5.1151e-14, 5.140191e-14, 
    5.133885e-14, 5.139894e-14, 5.138073e-14, 5.139918e-14, 5.130669e-14, 
    5.134632e-14, 5.126492e-14, 5.094728e-14, 5.10407e-14, 5.076183e-14, 
    5.059379e-14, 5.048214e-14, 5.040283e-14, 5.041405e-14, 5.043541e-14, 
    5.054522e-14, 5.064841e-14, 5.072698e-14, 5.07795e-14, 5.083124e-14, 
    5.09876e-14, 5.107037e-14, 5.125542e-14, 5.122208e-14, 5.127858e-14, 
    5.133258e-14, 5.142314e-14, 5.140825e-14, 5.144812e-14, 5.127711e-14, 
    5.139078e-14, 5.120307e-14, 5.125444e-14, 5.084517e-14, 5.068906e-14, 
    5.062253e-14, 5.056437e-14, 5.042267e-14, 5.052053e-14, 5.048196e-14, 
    5.057374e-14, 5.063201e-14, 5.06032e-14, 5.078094e-14, 5.071186e-14, 
    5.107527e-14, 5.091887e-14, 5.132628e-14, 5.122893e-14, 5.134961e-14, 
    5.128805e-14, 5.13935e-14, 5.12986e-14, 5.146297e-14, 5.149871e-14, 
    5.147428e-14, 5.156814e-14, 5.129333e-14, 5.139893e-14, 5.060239e-14, 
    5.060708e-14, 5.062899e-14, 5.053268e-14, 5.05268e-14, 5.043851e-14, 
    5.051708e-14, 5.055051e-14, 5.06354e-14, 5.068555e-14, 5.073322e-14, 
    5.083796e-14, 5.095482e-14, 5.111807e-14, 5.123524e-14, 5.131371e-14, 
    5.126561e-14, 5.130807e-14, 5.126059e-14, 5.123834e-14, 5.148531e-14, 
    5.134668e-14, 5.155464e-14, 5.154315e-14, 5.144906e-14, 5.154445e-14, 
    5.061038e-14, 5.058334e-14, 5.048937e-14, 5.056292e-14, 5.04289e-14, 
    5.050392e-14, 5.054702e-14, 5.071328e-14, 5.074981e-14, 5.078363e-14, 
    5.085044e-14, 5.09361e-14, 5.108622e-14, 5.121671e-14, 5.133573e-14, 
    5.132702e-14, 5.133008e-14, 5.135664e-14, 5.129082e-14, 5.136744e-14, 
    5.138028e-14, 5.134668e-14, 5.154161e-14, 5.148596e-14, 5.154291e-14, 
    5.150668e-14, 5.059214e-14, 5.063764e-14, 5.061305e-14, 5.065928e-14, 
    5.06267e-14, 5.077144e-14, 5.08148e-14, 5.101754e-14, 5.093441e-14, 
    5.106672e-14, 5.094787e-14, 5.096893e-14, 5.107098e-14, 5.09543e-14, 
    5.120949e-14, 5.103649e-14, 5.135767e-14, 5.118507e-14, 5.136848e-14, 
    5.133521e-14, 5.139029e-14, 5.143959e-14, 5.15016e-14, 5.161589e-14, 
    5.158944e-14, 5.168497e-14, 5.070545e-14, 5.07644e-14, 5.075924e-14, 
    5.082092e-14, 5.086651e-14, 5.09653e-14, 5.112355e-14, 5.106407e-14, 
    5.117327e-14, 5.119517e-14, 5.102928e-14, 5.113113e-14, 5.080386e-14, 
    5.085677e-14, 5.082528e-14, 5.071009e-14, 5.107774e-14, 5.088918e-14, 
    5.123717e-14, 5.11352e-14, 5.143256e-14, 5.128474e-14, 5.157487e-14, 
    5.169861e-14, 5.181506e-14, 5.195085e-14, 5.079659e-14, 5.075655e-14, 
    5.082826e-14, 5.092736e-14, 5.101932e-14, 5.114141e-14, 5.115391e-14, 
    5.117676e-14, 5.123596e-14, 5.12857e-14, 5.118396e-14, 5.129817e-14, 
    5.086898e-14, 5.109411e-14, 5.074138e-14, 5.084767e-14, 5.092153e-14, 
    5.088916e-14, 5.105728e-14, 5.109686e-14, 5.125756e-14, 5.117453e-14, 
    5.166806e-14, 5.144996e-14, 5.205423e-14, 5.188567e-14, 5.074255e-14, 
    5.079646e-14, 5.09839e-14, 5.089475e-14, 5.114957e-14, 5.12122e-14, 
    5.126311e-14, 5.132812e-14, 5.133515e-14, 5.137365e-14, 5.131056e-14, 
    5.137117e-14, 5.114167e-14, 5.124429e-14, 5.096252e-14, 5.103114e-14, 
    5.099959e-14, 5.096494e-14, 5.107183e-14, 5.118556e-14, 5.118803e-14, 
    5.122447e-14, 5.132701e-14, 5.115061e-14, 5.16961e-14, 5.135945e-14, 
    5.085523e-14, 5.095891e-14, 5.097376e-14, 5.093361e-14, 5.120592e-14, 
    5.110732e-14, 5.137272e-14, 5.130106e-14, 5.141846e-14, 5.136013e-14, 
    5.135155e-14, 5.12766e-14, 5.122989e-14, 5.111183e-14, 5.10157e-14, 
    5.093944e-14, 5.095718e-14, 5.104094e-14, 5.119252e-14, 5.133577e-14, 
    5.13044e-14, 5.140955e-14, 5.113111e-14, 5.124792e-14, 5.120278e-14, 
    5.132047e-14, 5.106248e-14, 5.128208e-14, 5.100627e-14, 5.103049e-14, 
    5.110536e-14, 5.125581e-14, 5.128914e-14, 5.132463e-14, 5.130274e-14, 
    5.119638e-14, 5.117896e-14, 5.110355e-14, 5.10827e-14, 5.102522e-14, 
    5.097758e-14, 5.102109e-14, 5.106677e-14, 5.119644e-14, 5.131315e-14, 
    5.144028e-14, 5.147139e-14, 5.161961e-14, 5.149891e-14, 5.169796e-14, 
    5.152867e-14, 5.182161e-14, 5.129486e-14, 5.152377e-14, 5.110878e-14, 
    5.115357e-14, 5.123449e-14, 5.141997e-14, 5.131992e-14, 5.143694e-14, 
    5.117828e-14, 5.104381e-14, 5.100904e-14, 5.094406e-14, 5.101053e-14, 
    5.100512e-14, 5.106868e-14, 5.104827e-14, 5.120074e-14, 5.111886e-14, 
    5.135132e-14, 5.143602e-14, 5.167495e-14, 5.182114e-14, 5.196983e-14, 
    5.203539e-14, 5.205534e-14, 5.206367e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.177466e-15, -7.166129e-15, -7.168332e-15, -7.1592e-15, -7.164266e-15, 
    -7.158286e-15, -7.175168e-15, -7.165679e-15, -7.171736e-15, 
    -7.176447e-15, -7.141511e-15, -7.158793e-15, -7.123634e-15, 
    -7.134613e-15, -7.107082e-15, -7.125339e-15, -7.103409e-15, 
    -7.107613e-15, -7.094982e-15, -7.098598e-15, -7.082464e-15, 
    -7.093314e-15, -7.074127e-15, -7.085056e-15, -7.083343e-15, 
    -7.093672e-15, -7.155315e-15, -7.143658e-15, -7.156005e-15, 
    -7.154342e-15, -7.15509e-15, -7.16416e-15, -7.168733e-15, -7.178337e-15, 
    -7.176593e-15, -7.169541e-15, -7.153594e-15, -7.159006e-15, 
    -7.145386e-15, -7.145694e-15, -7.130566e-15, -7.137382e-15, 
    -7.112019e-15, -7.119217e-15, -7.098447e-15, -7.103662e-15, 
    -7.098691e-15, -7.100199e-15, -7.098671e-15, -7.106323e-15, 
    -7.103043e-15, -7.109782e-15, -7.136104e-15, -7.128353e-15, 
    -7.151497e-15, -7.165452e-15, -7.17475e-15, -7.181355e-15, -7.18042e-15, 
    -7.178639e-15, -7.169499e-15, -7.160924e-15, -7.154396e-15, 
    -7.150033e-15, -7.145738e-15, -7.132744e-15, -7.125889e-15, 
    -7.110563e-15, -7.113329e-15, -7.108646e-15, -7.104182e-15, 
    -7.096689e-15, -7.097922e-15, -7.094622e-15, -7.108772e-15, 
    -7.099363e-15, -7.114905e-15, -7.110649e-15, -7.144555e-15, 
    -7.157546e-15, -7.163063e-15, -7.167909e-15, -7.179702e-15, 
    -7.171554e-15, -7.174765e-15, -7.167134e-15, -7.162288e-15, 
    -7.164684e-15, -7.149914e-15, -7.155651e-15, -7.125483e-15, 
    -7.138458e-15, -7.104702e-15, -7.112762e-15, -7.102773e-15, 
    -7.107869e-15, -7.099139e-15, -7.106995e-15, -7.093396e-15, 
    -7.090437e-15, -7.092459e-15, -7.084704e-15, -7.107431e-15, -7.09869e-15, 
    -7.164751e-15, -7.16436e-15, -7.16254e-15, -7.170543e-15, -7.171034e-15, 
    -7.178383e-15, -7.171845e-15, -7.169062e-15, -7.162008e-15, 
    -7.157838e-15, -7.153876e-15, -7.145177e-15, -7.135475e-15, -7.12194e-15, 
    -7.112239e-15, -7.105745e-15, -7.109727e-15, -7.106211e-15, 
    -7.110141e-15, -7.111984e-15, -7.091545e-15, -7.103011e-15, 
    -7.085819e-15, -7.086769e-15, -7.094543e-15, -7.086662e-15, 
    -7.164085e-15, -7.166336e-15, -7.17415e-15, -7.168034e-15, -7.179184e-15, 
    -7.172938e-15, -7.169349e-15, -7.155528e-15, -7.1525e-15, -7.149688e-15, 
    -7.144143e-15, -7.137033e-15, -7.12458e-15, -7.11377e-15, -7.103923e-15, 
    -7.104644e-15, -7.10439e-15, -7.10219e-15, -7.107638e-15, -7.101297e-15, 
    -7.100232e-15, -7.103015e-15, -7.086896e-15, -7.091497e-15, 
    -7.086789e-15, -7.089784e-15, -7.165605e-15, -7.16182e-15, -7.163864e-15, 
    -7.160019e-15, -7.162727e-15, -7.150694e-15, -7.147092e-15, -7.13027e-15, 
    -7.137172e-15, -7.126196e-15, -7.136057e-15, -7.134307e-15, 
    -7.125831e-15, -7.135524e-15, -7.114363e-15, -7.128695e-15, 
    -7.102105e-15, -7.116379e-15, -7.101212e-15, -7.103965e-15, 
    -7.099408e-15, -7.095329e-15, -7.090203e-15, -7.080754e-15, 
    -7.082941e-15, -7.075051e-15, -7.156184e-15, -7.151282e-15, 
    -7.151717e-15, -7.146593e-15, -7.142807e-15, -7.134612e-15, 
    -7.121489e-15, -7.126421e-15, -7.117373e-15, -7.115558e-15, 
    -7.129307e-15, -7.120858e-15, -7.148007e-15, -7.143608e-15, 
    -7.146229e-15, -7.155795e-15, -7.12528e-15, -7.140918e-15, -7.112078e-15, 
    -7.120525e-15, -7.09591e-15, -7.108134e-15, -7.084145e-15, -7.073914e-15, 
    -7.064317e-15, -7.053107e-15, -7.148612e-15, -7.15194e-15, -7.145986e-15, 
    -7.137751e-15, -7.130129e-15, -7.120009e-15, -7.118976e-15, 
    -7.117082e-15, -7.112181e-15, -7.108062e-15, -7.116479e-15, 
    -7.107031e-15, -7.142583e-15, -7.123926e-15, -7.153197e-15, 
    -7.144363e-15, -7.138237e-15, -7.140927e-15, -7.126986e-15, 
    -7.123704e-15, -7.110388e-15, -7.117269e-15, -7.076435e-15, 
    -7.094463e-15, -7.044598e-15, -7.058484e-15, -7.153103e-15, 
    -7.148625e-15, -7.133064e-15, -7.140463e-15, -7.119336e-15, 
    -7.114146e-15, -7.109934e-15, -7.104548e-15, -7.103969e-15, 
    -7.100782e-15, -7.106006e-15, -7.100989e-15, -7.119987e-15, -7.11149e-15, 
    -7.134844e-15, -7.129149e-15, -7.131769e-15, -7.134642e-15, 
    -7.125779e-15, -7.116346e-15, -7.11615e-15, -7.113128e-15, -7.104613e-15, 
    -7.11925e-15, -7.074103e-15, -7.101932e-15, -7.143746e-15, -7.135132e-15, 
    -7.133908e-15, -7.137242e-15, -7.114666e-15, -7.122835e-15, -7.10086e-15, 
    -7.106791e-15, -7.097078e-15, -7.101902e-15, -7.102612e-15, 
    -7.108816e-15, -7.112681e-15, -7.122459e-15, -7.130428e-15, 
    -7.136759e-15, -7.135287e-15, -7.128335e-15, -7.115771e-15, 
    -7.103915e-15, -7.106509e-15, -7.097815e-15, -7.120865e-15, 
    -7.111185e-15, -7.114923e-15, -7.105184e-15, -7.126552e-15, 
    -7.108336e-15, -7.131215e-15, -7.129206e-15, -7.122997e-15, 
    -7.110526e-15, -7.107778e-15, -7.104837e-15, -7.106652e-15, 
    -7.115454e-15, -7.116899e-15, -7.123149e-15, -7.124874e-15, 
    -7.129644e-15, -7.133594e-15, -7.129984e-15, -7.126193e-15, 
    -7.115452e-15, -7.105786e-15, -7.09527e-15, -7.092701e-15, -7.080432e-15, 
    -7.090411e-15, -7.073948e-15, -7.087931e-15, -7.063753e-15, 
    -7.107289e-15, -7.088353e-15, -7.122716e-15, -7.119005e-15, 
    -7.112293e-15, -7.096942e-15, -7.10523e-15, -7.095541e-15, -7.116955e-15, 
    -7.128093e-15, -7.130985e-15, -7.136373e-15, -7.130861e-15, 
    -7.131309e-15, -7.12604e-15, -7.127733e-15, -7.115095e-15, -7.12188e-15, 
    -7.102628e-15, -7.095618e-15, -7.075876e-15, -7.063806e-15, 
    -7.051555e-15, -7.046153e-15, -7.04451e-15, -7.043823e-15 ;

 CH4_SURF_DIFF_UNSAT =
  1.481542e-14, 1.438706e-14, 1.447035e-14, 1.412482e-14, 1.431651e-14, 
    1.409024e-14, 1.47286e-14, 1.437003e-14, 1.459895e-14, 1.477689e-14, 
    1.345416e-14, 1.410941e-14, 1.277366e-14, 1.319159e-14, 1.21417e-14, 
    1.283866e-14, 1.200116e-14, 1.216187e-14, 1.167828e-14, 1.181683e-14, 
    1.119805e-14, 1.161433e-14, 1.087731e-14, 1.129751e-14, 1.123176e-14, 
    1.162805e-14, 1.39776e-14, 1.353572e-14, 1.400377e-14, 1.394076e-14, 
    1.396904e-14, 1.431253e-14, 1.448559e-14, 1.484819e-14, 1.478237e-14, 
    1.451607e-14, 1.391243e-14, 1.411738e-14, 1.360095e-14, 1.361262e-14, 
    1.303759e-14, 1.329687e-14, 1.233029e-14, 1.260505e-14, 1.181105e-14, 
    1.201074e-14, 1.182042e-14, 1.187814e-14, 1.181967e-14, 1.211254e-14, 
    1.198706e-14, 1.224478e-14, 1.32483e-14, 1.295338e-14, 1.383288e-14, 
    1.436157e-14, 1.471286e-14, 1.49621e-14, 1.492686e-14, 1.485968e-14, 
    1.451451e-14, 1.419003e-14, 1.394273e-14, 1.37773e-14, 1.361429e-14, 
    1.312072e-14, 1.285958e-14, 1.22747e-14, 1.238031e-14, 1.220144e-14, 
    1.203061e-14, 1.174372e-14, 1.179095e-14, 1.166453e-14, 1.220619e-14, 
    1.18462e-14, 1.244045e-14, 1.227792e-14, 1.356979e-14, 1.40621e-14, 
    1.427118e-14, 1.445433e-14, 1.489977e-14, 1.459215e-14, 1.471341e-14, 
    1.442496e-14, 1.424165e-14, 1.433232e-14, 1.377277e-14, 1.399031e-14, 
    1.28441e-14, 1.333785e-14, 1.205054e-14, 1.235864e-14, 1.197669e-14, 
    1.217161e-14, 1.183761e-14, 1.213821e-14, 1.16175e-14, 1.150408e-14, 
    1.158158e-14, 1.128391e-14, 1.215486e-14, 1.18204e-14, 1.433485e-14, 
    1.432006e-14, 1.425118e-14, 1.455395e-14, 1.457248e-14, 1.484999e-14, 
    1.460308e-14, 1.449792e-14, 1.423104e-14, 1.407314e-14, 1.392305e-14, 
    1.359304e-14, 1.322443e-14, 1.270899e-14, 1.233866e-14, 1.209039e-14, 
    1.224265e-14, 1.210823e-14, 1.225848e-14, 1.232891e-14, 1.154656e-14, 
    1.198588e-14, 1.132672e-14, 1.136321e-14, 1.166152e-14, 1.13591e-14, 
    1.430968e-14, 1.439478e-14, 1.469018e-14, 1.4459e-14, 1.488021e-14, 
    1.464442e-14, 1.450882e-14, 1.398572e-14, 1.387083e-14, 1.376424e-14, 
    1.355376e-14, 1.32836e-14, 1.280962e-14, 1.23972e-14, 1.202068e-14, 
    1.204827e-14, 1.203856e-14, 1.195442e-14, 1.21628e-14, 1.192021e-14, 
    1.187948e-14, 1.198595e-14, 1.13681e-14, 1.154463e-14, 1.136399e-14, 
    1.147894e-14, 1.436712e-14, 1.422394e-14, 1.430131e-14, 1.415581e-14, 
    1.42583e-14, 1.380252e-14, 1.366586e-14, 1.302641e-14, 1.32889e-14, 
    1.287119e-14, 1.324649e-14, 1.317998e-14, 1.285749e-14, 1.322622e-14, 
    1.24199e-14, 1.296651e-14, 1.195115e-14, 1.2497e-14, 1.191694e-14, 
    1.202231e-14, 1.184786e-14, 1.169159e-14, 1.149502e-14, 1.11322e-14, 
    1.121623e-14, 1.091281e-14, 1.40105e-14, 1.382476e-14, 1.384115e-14, 
    1.364679e-14, 1.350304e-14, 1.319151e-14, 1.269175e-14, 1.28797e-14, 
    1.253469e-14, 1.246541e-14, 1.298959e-14, 1.266772e-14, 1.370048e-14, 
    1.35336e-14, 1.363299e-14, 1.399583e-14, 1.283634e-14, 1.34314e-14, 
    1.233254e-14, 1.265497e-14, 1.171387e-14, 1.21819e-14, 1.126248e-14, 
    1.086922e-14, 1.049919e-14, 1.006647e-14, 1.372343e-14, 1.384963e-14, 
    1.362369e-14, 1.331101e-14, 1.302097e-14, 1.263529e-14, 1.259585e-14, 
    1.252358e-14, 1.233642e-14, 1.217903e-14, 1.25007e-14, 1.213958e-14, 
    1.349483e-14, 1.27847e-14, 1.389731e-14, 1.356226e-14, 1.332946e-14, 
    1.343162e-14, 1.290119e-14, 1.277615e-14, 1.226798e-14, 1.25307e-14, 
    1.096625e-14, 1.165853e-14, 9.737039e-15, 1.02742e-14, 1.389372e-14, 
    1.372388e-14, 1.31327e-14, 1.3414e-14, 1.260957e-14, 1.241151e-14, 
    1.225053e-14, 1.204467e-14, 1.202248e-14, 1.19005e-14, 1.210037e-14, 
    1.190841e-14, 1.263447e-14, 1.231004e-14, 1.320032e-14, 1.298363e-14, 
    1.308333e-14, 1.319266e-14, 1.285522e-14, 1.249562e-14, 1.2488e-14, 
    1.237267e-14, 1.204757e-14, 1.260631e-14, 1.087677e-14, 1.194494e-14, 
    1.353867e-14, 1.321143e-14, 1.316476e-14, 1.329152e-14, 1.243137e-14, 
    1.274305e-14, 1.190348e-14, 1.213043e-14, 1.175859e-14, 1.194336e-14, 
    1.197054e-14, 1.220785e-14, 1.235557e-14, 1.272875e-14, 1.303237e-14, 
    1.327314e-14, 1.321716e-14, 1.295267e-14, 1.247364e-14, 1.202044e-14, 
    1.211971e-14, 1.178685e-14, 1.26679e-14, 1.229846e-14, 1.244124e-14, 
    1.206895e-14, 1.288468e-14, 1.218988e-14, 1.306223e-14, 1.298577e-14, 
    1.274923e-14, 1.227336e-14, 1.216816e-14, 1.205572e-14, 1.212511e-14, 
    1.246149e-14, 1.251662e-14, 1.2755e-14, 1.282078e-14, 1.300242e-14, 
    1.315277e-14, 1.301539e-14, 1.28711e-14, 1.246137e-14, 1.209205e-14, 
    1.168936e-14, 1.159082e-14, 1.112006e-14, 1.150321e-14, 1.087081e-14, 
    1.140836e-14, 1.04778e-14, 1.21497e-14, 1.142428e-14, 1.273849e-14, 
    1.259695e-14, 1.234087e-14, 1.175356e-14, 1.207071e-14, 1.169983e-14, 
    1.251878e-14, 1.294352e-14, 1.305347e-14, 1.325849e-14, 1.304878e-14, 
    1.306584e-14, 1.286516e-14, 1.292966e-14, 1.244777e-14, 1.270663e-14, 
    1.197121e-14, 1.170277e-14, 1.094459e-14, 1.047961e-14, 1.000627e-14, 
    9.797218e-15, 9.733591e-15, 9.706988e-15 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.93195e-23, 1.931952e-23, 1.931949e-23, 1.93195e-23, 1.931947e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931945e-23, 
    1.931946e-23, 1.931951e-23, 1.93195e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931951e-23, 1.931952e-23, 1.93195e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.93195e-23, 1.931949e-23, 1.931951e-23, 
    1.931952e-23, 1.931953e-23, 1.931954e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.93195e-23, 
    1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.93195e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931947e-23, 1.931946e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931945e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931946e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.93195e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931948e-23, 1.931951e-23, 
    1.93195e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 
    1.931944e-23, 1.931943e-23, 1.931942e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.93195e-23, 1.931949e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 
    1.931944e-23, 1.931946e-23, 1.931942e-23, 1.931943e-23, 1.931951e-23, 
    1.931951e-23, 1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931948e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931944e-23, 1.931947e-23, 
    1.93195e-23, 1.93195e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931944e-23, 
    1.931945e-23, 1.931943e-23, 1.931947e-23, 1.931946e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 
    1.931948e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931946e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975384e-24, 1.975386e-24, 1.975381e-24, 1.975383e-24, 1.975379e-24, 
    1.975382e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975376e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 1.975377e-24, 
    1.975378e-24, 1.975385e-24, 1.975384e-24, 1.975385e-24, 1.975385e-24, 
    1.975385e-24, 1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975385e-24, 1.975386e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975383e-24, 1.97538e-24, 1.975381e-24, 1.975378e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 1.975385e-24, 
    1.975387e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 
    1.975383e-24, 1.975382e-24, 1.97538e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 1.97538e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975384e-24, 1.975386e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975382e-24, 1.975383e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 
    1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975379e-24, 1.975386e-24, 
    1.975386e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975377e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975385e-24, 1.975384e-24, 1.975382e-24, 1.975383e-24, 
    1.975382e-24, 1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975383e-24, 
    1.97538e-24, 1.975382e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975376e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975384e-24, 1.975383e-24, 1.975381e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975382e-24, 1.975381e-24, 1.975384e-24, 
    1.975384e-24, 1.975384e-24, 1.975385e-24, 1.975382e-24, 1.975384e-24, 
    1.97538e-24, 1.975381e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 
    1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975384e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975384e-24, 1.975381e-24, 1.975385e-24, 1.975384e-24, 1.975383e-24, 
    1.975384e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.975376e-24, 1.975378e-24, 1.975372e-24, 1.975373e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975375e-24, 1.975379e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975383e-24, 1.97538e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 1.975382e-24, 
    1.975383e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975382e-24, 1.97538e-24, 1.975382e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975382e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975378e-24, 1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975375e-24, 
    1.975377e-24, 1.975374e-24, 1.975379e-24, 1.975377e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 
    1.975381e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975381e-24, 
    1.975379e-24, 1.975378e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24 ;

 CONC_CH4_SAT =
  3.291541e-08, 3.289345e-08, 3.289773e-08, 3.288e-08, 3.288985e-08, 
    3.287823e-08, 3.291098e-08, 3.289256e-08, 3.290432e-08, 3.291346e-08, 
    3.284558e-08, 3.287921e-08, 3.281087e-08, 3.283225e-08, 3.277863e-08, 
    3.281417e-08, 3.277147e-08, 3.277969e-08, 3.275506e-08, 3.276212e-08, 
    3.273056e-08, 3.275181e-08, 3.271429e-08, 3.273566e-08, 3.27323e-08, 
    3.27525e-08, 3.287248e-08, 3.284975e-08, 3.287382e-08, 3.287058e-08, 
    3.287204e-08, 3.288963e-08, 3.289847e-08, 3.291712e-08, 3.291374e-08, 
    3.290006e-08, 3.286912e-08, 3.287965e-08, 3.285321e-08, 3.285381e-08, 
    3.282438e-08, 3.283765e-08, 3.278828e-08, 3.280231e-08, 3.276183e-08, 
    3.277199e-08, 3.27623e-08, 3.276524e-08, 3.276226e-08, 3.277717e-08, 
    3.277078e-08, 3.278392e-08, 3.283516e-08, 3.282008e-08, 3.286506e-08, 
    3.289209e-08, 3.291016e-08, 3.292296e-08, 3.292115e-08, 3.291769e-08, 
    3.289998e-08, 3.288337e-08, 3.287071e-08, 3.286224e-08, 3.285389e-08, 
    3.282856e-08, 3.281526e-08, 3.278542e-08, 3.279084e-08, 3.278169e-08, 
    3.277301e-08, 3.275839e-08, 3.27608e-08, 3.275435e-08, 3.278196e-08, 
    3.276359e-08, 3.279392e-08, 3.278561e-08, 3.285149e-08, 3.287681e-08, 
    3.288747e-08, 3.28969e-08, 3.291976e-08, 3.290396e-08, 3.291018e-08, 
    3.289541e-08, 3.288601e-08, 3.289067e-08, 3.2862e-08, 3.287314e-08, 
    3.281447e-08, 3.283972e-08, 3.277402e-08, 3.278973e-08, 3.277026e-08, 
    3.27802e-08, 3.276316e-08, 3.27785e-08, 3.275196e-08, 3.274617e-08, 
    3.275013e-08, 3.273499e-08, 3.277934e-08, 3.276228e-08, 3.289079e-08, 
    3.289003e-08, 3.288651e-08, 3.2902e-08, 3.290296e-08, 3.291721e-08, 
    3.290454e-08, 3.289913e-08, 3.288548e-08, 3.287738e-08, 3.286969e-08, 
    3.28528e-08, 3.283392e-08, 3.280759e-08, 3.278871e-08, 3.277606e-08, 
    3.278383e-08, 3.277697e-08, 3.278463e-08, 3.278823e-08, 3.274833e-08, 
    3.277071e-08, 3.273717e-08, 3.273903e-08, 3.275419e-08, 3.273882e-08, 
    3.28895e-08, 3.289387e-08, 3.2909e-08, 3.289716e-08, 3.291876e-08, 
    3.290665e-08, 3.289968e-08, 3.287287e-08, 3.286702e-08, 3.286155e-08, 
    3.285079e-08, 3.283697e-08, 3.281273e-08, 3.279168e-08, 3.277251e-08, 
    3.277392e-08, 3.277342e-08, 3.276912e-08, 3.277975e-08, 3.276738e-08, 
    3.276529e-08, 3.277073e-08, 3.273928e-08, 3.274826e-08, 3.273907e-08, 
    3.274492e-08, 3.289245e-08, 3.288511e-08, 3.288907e-08, 3.28816e-08, 
    3.288686e-08, 3.286349e-08, 3.285648e-08, 3.282378e-08, 3.283723e-08, 
    3.281587e-08, 3.283507e-08, 3.283166e-08, 3.281511e-08, 3.283404e-08, 
    3.279282e-08, 3.28207e-08, 3.276896e-08, 3.279672e-08, 3.276721e-08, 
    3.277259e-08, 3.27637e-08, 3.275573e-08, 3.274573e-08, 3.272725e-08, 
    3.273153e-08, 3.271612e-08, 3.287417e-08, 3.286464e-08, 3.28655e-08, 
    3.285555e-08, 3.284819e-08, 3.283226e-08, 3.280672e-08, 3.281633e-08, 
    3.279872e-08, 3.279518e-08, 3.282195e-08, 3.280548e-08, 3.285828e-08, 
    3.284972e-08, 3.285484e-08, 3.287341e-08, 3.281408e-08, 3.284449e-08, 
    3.278839e-08, 3.280485e-08, 3.275687e-08, 3.278069e-08, 3.273389e-08, 
    3.271384e-08, 3.269511e-08, 3.26731e-08, 3.285947e-08, 3.286594e-08, 
    3.285438e-08, 3.283834e-08, 3.282354e-08, 3.280384e-08, 3.280184e-08, 
    3.279814e-08, 3.278861e-08, 3.278058e-08, 3.279695e-08, 3.277857e-08, 
    3.284768e-08, 3.281146e-08, 3.286836e-08, 3.285118e-08, 3.283929e-08, 
    3.284453e-08, 3.281744e-08, 3.281105e-08, 3.278509e-08, 3.279852e-08, 
    3.271877e-08, 3.275401e-08, 3.265644e-08, 3.268365e-08, 3.28682e-08, 
    3.28595e-08, 3.282923e-08, 3.284363e-08, 3.280254e-08, 3.279242e-08, 
    3.278423e-08, 3.277371e-08, 3.277259e-08, 3.276637e-08, 3.277657e-08, 
    3.276678e-08, 3.28038e-08, 3.278725e-08, 3.283272e-08, 3.282163e-08, 
    3.282674e-08, 3.283233e-08, 3.281509e-08, 3.279669e-08, 3.279634e-08, 
    3.279043e-08, 3.277373e-08, 3.280238e-08, 3.271414e-08, 3.276852e-08, 
    3.285002e-08, 3.283324e-08, 3.283089e-08, 3.283738e-08, 3.279344e-08, 
    3.280935e-08, 3.276653e-08, 3.27781e-08, 3.275915e-08, 3.276856e-08, 
    3.276995e-08, 3.278205e-08, 3.278958e-08, 3.280861e-08, 3.282412e-08, 
    3.283645e-08, 3.283358e-08, 3.282004e-08, 3.279557e-08, 3.277248e-08, 
    3.277752e-08, 3.276059e-08, 3.280552e-08, 3.278664e-08, 3.279392e-08, 
    3.277496e-08, 3.281658e-08, 3.2781e-08, 3.282566e-08, 3.282176e-08, 
    3.280966e-08, 3.278534e-08, 3.278002e-08, 3.277427e-08, 3.277783e-08, 
    3.279496e-08, 3.279779e-08, 3.280996e-08, 3.281331e-08, 3.282261e-08, 
    3.283029e-08, 3.282326e-08, 3.281587e-08, 3.279497e-08, 3.277612e-08, 
    3.275561e-08, 3.275061e-08, 3.272657e-08, 3.274608e-08, 3.271383e-08, 
    3.274116e-08, 3.269392e-08, 3.277901e-08, 3.274205e-08, 3.280913e-08, 
    3.28019e-08, 3.278879e-08, 3.275884e-08, 3.277505e-08, 3.275612e-08, 
    3.27979e-08, 3.281955e-08, 3.282521e-08, 3.283569e-08, 3.282497e-08, 
    3.282585e-08, 3.28156e-08, 3.281889e-08, 3.279428e-08, 3.28075e-08, 
    3.276997e-08, 3.275628e-08, 3.271771e-08, 3.269408e-08, 3.26701e-08, 
    3.265951e-08, 3.265629e-08, 3.265494e-08,
  5.414219e-11, 5.416548e-11, 5.4161e-11, 5.417967e-11, 5.416937e-11, 
    5.418155e-11, 5.414699e-11, 5.416634e-11, 5.415403e-11, 5.414439e-11, 
    5.421563e-11, 5.418052e-11, 5.425267e-11, 5.423025e-11, 5.428671e-11, 
    5.424908e-11, 5.429431e-11, 5.428579e-11, 5.431182e-11, 5.430438e-11, 
    5.433726e-11, 5.431525e-11, 5.435455e-11, 5.43321e-11, 5.433555e-11, 
    5.43145e-11, 5.418775e-11, 5.421121e-11, 5.418632e-11, 5.418968e-11, 
    5.418821e-11, 5.416953e-11, 5.416e-11, 5.414052e-11, 5.414409e-11, 
    5.415846e-11, 5.419119e-11, 5.41802e-11, 5.42082e-11, 5.420758e-11, 
    5.423858e-11, 5.422461e-11, 5.427672e-11, 5.426197e-11, 5.430469e-11, 
    5.429394e-11, 5.430416e-11, 5.430108e-11, 5.43042e-11, 5.428843e-11, 
    5.429518e-11, 5.428135e-11, 5.42272e-11, 5.424308e-11, 5.419555e-11, 
    5.416664e-11, 5.414781e-11, 5.41343e-11, 5.413621e-11, 5.413982e-11, 
    5.415854e-11, 5.417625e-11, 5.418969e-11, 5.419864e-11, 5.420748e-11, 
    5.423378e-11, 5.424804e-11, 5.427963e-11, 5.427407e-11, 5.428359e-11, 
    5.429287e-11, 5.430826e-11, 5.430575e-11, 5.431249e-11, 5.428344e-11, 
    5.43027e-11, 5.427087e-11, 5.427957e-11, 5.420933e-11, 5.418319e-11, 
    5.417158e-11, 5.416184e-11, 5.413767e-11, 5.415433e-11, 5.414776e-11, 
    5.416352e-11, 5.417345e-11, 5.416856e-11, 5.419889e-11, 5.418709e-11, 
    5.424888e-11, 5.42223e-11, 5.429179e-11, 5.427522e-11, 5.429578e-11, 
    5.428532e-11, 5.430319e-11, 5.428711e-11, 5.431504e-11, 5.432105e-11, 
    5.431693e-11, 5.433293e-11, 5.42862e-11, 5.430411e-11, 5.41684e-11, 
    5.416919e-11, 5.417295e-11, 5.41564e-11, 5.415542e-11, 5.414039e-11, 
    5.415381e-11, 5.415948e-11, 5.417406e-11, 5.418258e-11, 5.419071e-11, 
    5.420858e-11, 5.422841e-11, 5.425624e-11, 5.427629e-11, 5.428968e-11, 
    5.428151e-11, 5.428872e-11, 5.428064e-11, 5.427687e-11, 5.431876e-11, 
    5.429521e-11, 5.433063e-11, 5.432869e-11, 5.431263e-11, 5.432892e-11, 
    5.416976e-11, 5.416517e-11, 5.414906e-11, 5.416167e-11, 5.413876e-11, 
    5.415152e-11, 5.415881e-11, 5.418721e-11, 5.419358e-11, 5.41993e-11, 
    5.421073e-11, 5.422532e-11, 5.425084e-11, 5.427308e-11, 5.429344e-11, 
    5.429196e-11, 5.429247e-11, 5.429696e-11, 5.428577e-11, 5.42988e-11, 
    5.430093e-11, 5.429527e-11, 5.432843e-11, 5.431898e-11, 5.432865e-11, 
    5.432251e-11, 5.416667e-11, 5.417441e-11, 5.417022e-11, 5.417808e-11, 
    5.41725e-11, 5.419711e-11, 5.420447e-11, 5.423904e-11, 5.4225e-11, 
    5.424749e-11, 5.422733e-11, 5.423087e-11, 5.424799e-11, 5.422846e-11, 
    5.427175e-11, 5.424221e-11, 5.429714e-11, 5.426747e-11, 5.429898e-11, 
    5.429335e-11, 5.430272e-11, 5.431105e-11, 5.432162e-11, 5.434095e-11, 
    5.43365e-11, 5.435273e-11, 5.4186e-11, 5.419597e-11, 5.419519e-11, 
    5.42057e-11, 5.421344e-11, 5.423032e-11, 5.425724e-11, 5.424716e-11, 
    5.426578e-11, 5.426947e-11, 5.424125e-11, 5.425849e-11, 5.420272e-11, 
    5.421164e-11, 5.42064e-11, 5.418672e-11, 5.424934e-11, 5.421718e-11, 
    5.42766e-11, 5.425925e-11, 5.430985e-11, 5.42846e-11, 5.433402e-11, 
    5.435482e-11, 5.438006e-11, 5.44091e-11, 5.420152e-11, 5.419474e-11, 
    5.420698e-11, 5.42237e-11, 5.423949e-11, 5.426029e-11, 5.426247e-11, 
    5.426633e-11, 5.427646e-11, 5.428491e-11, 5.426745e-11, 5.428704e-11, 
    5.421349e-11, 5.425218e-11, 5.419207e-11, 5.421006e-11, 5.422276e-11, 
    5.42173e-11, 5.424603e-11, 5.425276e-11, 5.428002e-11, 5.426599e-11, 
    5.43496e-11, 5.431266e-11, 5.443151e-11, 5.439511e-11, 5.419234e-11, 
    5.420155e-11, 5.423339e-11, 5.421827e-11, 5.426173e-11, 5.427236e-11, 
    5.428109e-11, 5.429206e-11, 5.429332e-11, 5.429983e-11, 5.428915e-11, 
    5.429945e-11, 5.426033e-11, 5.427784e-11, 5.422988e-11, 5.424151e-11, 
    5.42362e-11, 5.423029e-11, 5.42485e-11, 5.42677e-11, 5.426828e-11, 
    5.42744e-11, 5.429134e-11, 5.426191e-11, 5.435405e-11, 5.429694e-11, 
    5.421157e-11, 5.422904e-11, 5.423174e-11, 5.422494e-11, 5.427129e-11, 
    5.425449e-11, 5.42997e-11, 5.428753e-11, 5.43075e-11, 5.429757e-11, 
    5.42961e-11, 5.428336e-11, 5.427539e-11, 5.425523e-11, 5.423886e-11, 
    5.422595e-11, 5.422896e-11, 5.424315e-11, 5.426891e-11, 5.429336e-11, 
    5.428799e-11, 5.430599e-11, 5.425858e-11, 5.427839e-11, 5.427068e-11, 
    5.429081e-11, 5.424685e-11, 5.428379e-11, 5.423734e-11, 5.424145e-11, 
    5.425416e-11, 5.427962e-11, 5.42855e-11, 5.429147e-11, 5.428782e-11, 
    5.42696e-11, 5.426668e-11, 5.425389e-11, 5.425027e-11, 5.424057e-11, 
    5.423244e-11, 5.423982e-11, 5.424753e-11, 5.426968e-11, 5.42895e-11, 
    5.431115e-11, 5.43165e-11, 5.434131e-11, 5.432089e-11, 5.435433e-11, 
    5.432555e-11, 5.438101e-11, 5.428617e-11, 5.432505e-11, 5.42548e-11, 
    5.426242e-11, 5.427603e-11, 5.430754e-11, 5.429071e-11, 5.431047e-11, 
    5.426658e-11, 5.424355e-11, 5.423779e-11, 5.42267e-11, 5.423805e-11, 
    5.423713e-11, 5.424797e-11, 5.42445e-11, 5.427041e-11, 5.425651e-11, 
    5.429602e-11, 5.431035e-11, 5.435097e-11, 5.438119e-11, 5.441342e-11, 
    5.442752e-11, 5.443183e-11, 5.443362e-11,
  2.421313e-14, 2.425105e-14, 2.42437e-14, 2.427424e-14, 2.425734e-14, 
    2.42773e-14, 2.422086e-14, 2.425251e-14, 2.423234e-14, 2.421661e-14, 
    2.433339e-14, 2.427561e-14, 2.439397e-14, 2.435699e-14, 2.445007e-14, 
    2.438814e-14, 2.446259e-14, 2.44484e-14, 2.449139e-14, 2.447908e-14, 
    2.453385e-14, 2.449708e-14, 2.456244e-14, 2.452513e-14, 2.453092e-14, 
    2.449585e-14, 2.428735e-14, 2.432616e-14, 2.428502e-14, 2.429056e-14, 
    2.42881e-14, 2.425765e-14, 2.424223e-14, 2.421031e-14, 2.421612e-14, 
    2.423961e-14, 2.429306e-14, 2.427499e-14, 2.432077e-14, 2.431974e-14, 
    2.437066e-14, 2.434769e-14, 2.443345e-14, 2.440909e-14, 2.44796e-14, 
    2.446184e-14, 2.447874e-14, 2.447363e-14, 2.447881e-14, 2.445278e-14, 
    2.446392e-14, 2.444106e-14, 2.435197e-14, 2.43781e-14, 2.430014e-14, 
    2.425314e-14, 2.422223e-14, 2.420022e-14, 2.420333e-14, 2.420924e-14, 
    2.423975e-14, 2.426855e-14, 2.429048e-14, 2.430513e-14, 2.431958e-14, 
    2.436306e-14, 2.438634e-14, 2.443832e-14, 2.442903e-14, 2.444484e-14, 
    2.446008e-14, 2.448554e-14, 2.448137e-14, 2.449256e-14, 2.444449e-14, 
    2.44764e-14, 2.442372e-14, 2.443811e-14, 2.432312e-14, 2.427988e-14, 
    2.426117e-14, 2.42451e-14, 2.420572e-14, 2.423289e-14, 2.422217e-14, 
    2.424776e-14, 2.426398e-14, 2.425597e-14, 2.430553e-14, 2.428624e-14, 
    2.438773e-14, 2.434399e-14, 2.44583e-14, 2.443095e-14, 2.446487e-14, 
    2.444758e-14, 2.447718e-14, 2.445054e-14, 2.449677e-14, 2.450679e-14, 
    2.449993e-14, 2.452641e-14, 2.444905e-14, 2.44787e-14, 2.425573e-14, 
    2.425703e-14, 2.426315e-14, 2.423626e-14, 2.423464e-14, 2.421013e-14, 
    2.423197e-14, 2.424124e-14, 2.426495e-14, 2.42789e-14, 2.429219e-14, 
    2.432143e-14, 2.435403e-14, 2.439977e-14, 2.443271e-14, 2.445479e-14, 
    2.444128e-14, 2.44532e-14, 2.443986e-14, 2.443362e-14, 2.450301e-14, 
    2.4464e-14, 2.45226e-14, 2.451937e-14, 2.449281e-14, 2.451974e-14, 
    2.425795e-14, 2.425044e-14, 2.422425e-14, 2.424475e-14, 2.420747e-14, 
    2.422828e-14, 2.424023e-14, 2.428656e-14, 2.429684e-14, 2.430625e-14, 
    2.432493e-14, 2.434887e-14, 2.439086e-14, 2.442748e-14, 2.446098e-14, 
    2.445854e-14, 2.445939e-14, 2.446684e-14, 2.444834e-14, 2.446988e-14, 
    2.447346e-14, 2.446405e-14, 2.451894e-14, 2.450326e-14, 2.45193e-14, 
    2.45091e-14, 2.42529e-14, 2.426555e-14, 2.425871e-14, 2.427155e-14, 
    2.426247e-14, 2.430276e-14, 2.431485e-14, 2.437155e-14, 2.434837e-14, 
    2.438537e-14, 2.435216e-14, 2.435802e-14, 2.438641e-14, 2.435398e-14, 
    2.442538e-14, 2.437682e-14, 2.446713e-14, 2.441844e-14, 2.447017e-14, 
    2.446084e-14, 2.447633e-14, 2.449017e-14, 2.450766e-14, 2.453982e-14, 
    2.453238e-14, 2.455935e-14, 2.428446e-14, 2.430085e-14, 2.429948e-14, 
    2.431668e-14, 2.43294e-14, 2.435705e-14, 2.440135e-14, 2.438471e-14, 
    2.441534e-14, 2.442147e-14, 2.437498e-14, 2.440345e-14, 2.431187e-14, 
    2.432658e-14, 2.431788e-14, 2.428571e-14, 2.438844e-14, 2.433565e-14, 
    2.443324e-14, 2.440464e-14, 2.448819e-14, 2.444654e-14, 2.452828e-14, 
    2.456305e-14, 2.45992e-14, 2.464115e-14, 2.430987e-14, 2.429873e-14, 
    2.431875e-14, 2.434633e-14, 2.437215e-14, 2.440636e-14, 2.440991e-14, 
    2.44163e-14, 2.443295e-14, 2.444691e-14, 2.441825e-14, 2.445042e-14, 
    2.432984e-14, 2.439306e-14, 2.429444e-14, 2.432402e-14, 2.434474e-14, 
    2.433573e-14, 2.438283e-14, 2.439391e-14, 2.443893e-14, 2.44157e-14, 
    2.45544e-14, 2.449299e-14, 2.467336e-14, 2.462097e-14, 2.429482e-14, 
    2.430987e-14, 2.436219e-14, 2.43373e-14, 2.440869e-14, 2.442624e-14, 
    2.444058e-14, 2.445879e-14, 2.446081e-14, 2.447161e-14, 2.44539e-14, 
    2.447094e-14, 2.440644e-14, 2.443527e-14, 2.43563e-14, 2.437546e-14, 
    2.436667e-14, 2.435697e-14, 2.43869e-14, 2.441868e-14, 2.441948e-14, 
    2.442965e-14, 2.445811e-14, 2.440898e-14, 2.45621e-14, 2.446729e-14, 
    2.432628e-14, 2.435513e-14, 2.43594e-14, 2.43482e-14, 2.442448e-14, 
    2.439681e-14, 2.447137e-14, 2.445123e-14, 2.448425e-14, 2.446783e-14, 
    2.446541e-14, 2.444436e-14, 2.443122e-14, 2.439806e-14, 2.437113e-14, 
    2.434984e-14, 2.43548e-14, 2.437819e-14, 2.442065e-14, 2.446094e-14, 
    2.445209e-14, 2.448175e-14, 2.440351e-14, 2.443624e-14, 2.442355e-14, 
    2.445667e-14, 2.438424e-14, 2.444555e-14, 2.436854e-14, 2.437532e-14, 
    2.439626e-14, 2.443838e-14, 2.444788e-14, 2.445781e-14, 2.445171e-14, 
    2.442175e-14, 2.44169e-14, 2.439579e-14, 2.43899e-14, 2.437385e-14, 
    2.436051e-14, 2.437267e-14, 2.438541e-14, 2.442182e-14, 2.445457e-14, 
    2.449035e-14, 2.449916e-14, 2.454068e-14, 2.450671e-14, 2.45626e-14, 
    2.451482e-14, 2.460092e-14, 2.444928e-14, 2.451367e-14, 2.439726e-14, 
    2.440982e-14, 2.443241e-14, 2.448453e-14, 2.445652e-14, 2.448934e-14, 
    2.441672e-14, 2.437893e-14, 2.436931e-14, 2.435111e-14, 2.436973e-14, 
    2.436822e-14, 2.438603e-14, 2.438031e-14, 2.442303e-14, 2.440008e-14, 
    2.446532e-14, 2.448911e-14, 2.455648e-14, 2.460096e-14, 2.46472e-14, 
    2.466755e-14, 2.467376e-14, 2.467634e-14,
  3.249557e-18, 3.257782e-18, 3.256186e-18, 3.263073e-18, 3.259152e-18, 
    3.263785e-18, 3.251232e-18, 3.258101e-18, 3.25372e-18, 3.250309e-18, 
    3.276824e-18, 3.263392e-18, 3.290908e-18, 3.282294e-18, 3.303993e-18, 
    3.289555e-18, 3.306914e-18, 3.303597e-18, 3.313639e-18, 3.310761e-18, 
    3.323586e-18, 3.314968e-18, 3.330283e-18, 3.321538e-18, 3.322897e-18, 
    3.314681e-18, 3.266111e-18, 3.275143e-18, 3.265572e-18, 3.26686e-18, 
    3.266286e-18, 3.259225e-18, 3.255872e-18, 3.248943e-18, 3.250204e-18, 
    3.255301e-18, 3.267439e-18, 3.263242e-18, 3.273868e-18, 3.273628e-18, 
    3.285475e-18, 3.280129e-18, 3.300106e-18, 3.294423e-18, 3.310881e-18, 
    3.306733e-18, 3.310683e-18, 3.309488e-18, 3.310699e-18, 3.304618e-18, 
    3.307221e-18, 3.301881e-18, 3.281126e-18, 3.287209e-18, 3.269082e-18, 
    3.258243e-18, 3.25153e-18, 3.246758e-18, 3.247432e-18, 3.248714e-18, 
    3.255331e-18, 3.26175e-18, 3.266834e-18, 3.270236e-18, 3.273593e-18, 
    3.283719e-18, 3.289133e-18, 3.301246e-18, 3.299075e-18, 3.302767e-18, 
    3.306322e-18, 3.312273e-18, 3.311296e-18, 3.313916e-18, 3.302682e-18, 
    3.310138e-18, 3.297834e-18, 3.301194e-18, 3.274437e-18, 3.264377e-18, 
    3.260049e-18, 3.256491e-18, 3.247949e-18, 3.253842e-18, 3.251516e-18, 
    3.257066e-18, 3.260689e-18, 3.258848e-18, 3.270329e-18, 3.265853e-18, 
    3.289454e-18, 3.279273e-18, 3.305907e-18, 3.299522e-18, 3.307442e-18, 
    3.303402e-18, 3.31032e-18, 3.304094e-18, 3.314897e-18, 3.317244e-18, 
    3.315639e-18, 3.321835e-18, 3.303747e-18, 3.310676e-18, 3.258796e-18, 
    3.25908e-18, 3.260497e-18, 3.254574e-18, 3.254221e-18, 3.248905e-18, 
    3.253641e-18, 3.255654e-18, 3.260913e-18, 3.26415e-18, 3.267234e-18, 
    3.274023e-18, 3.281608e-18, 3.292257e-18, 3.299934e-18, 3.305085e-18, 
    3.301931e-18, 3.304715e-18, 3.3016e-18, 3.300144e-18, 3.31636e-18, 
    3.307241e-18, 3.320943e-18, 3.320186e-18, 3.313975e-18, 3.320272e-18, 
    3.259293e-18, 3.257648e-18, 3.251968e-18, 3.256412e-18, 3.248328e-18, 
    3.252842e-18, 3.255435e-18, 3.265932e-18, 3.268312e-18, 3.270498e-18, 
    3.274837e-18, 3.280402e-18, 3.290179e-18, 3.298715e-18, 3.306532e-18, 
    3.30596e-18, 3.306161e-18, 3.307901e-18, 3.303581e-18, 3.308612e-18, 
    3.30945e-18, 3.307248e-18, 3.320084e-18, 3.316414e-18, 3.32017e-18, 
    3.317782e-18, 3.25818e-18, 3.261054e-18, 3.259467e-18, 3.262448e-18, 
    3.260342e-18, 3.269695e-18, 3.272503e-18, 3.285687e-18, 3.280289e-18, 
    3.288903e-18, 3.281168e-18, 3.282534e-18, 3.289155e-18, 3.281591e-18, 
    3.29823e-18, 3.286916e-18, 3.307969e-18, 3.296617e-18, 3.30868e-18, 
    3.306498e-18, 3.310118e-18, 3.313355e-18, 3.317444e-18, 3.324978e-18, 
    3.323235e-18, 3.329554e-18, 3.265439e-18, 3.269246e-18, 3.268924e-18, 
    3.272921e-18, 3.275876e-18, 3.282305e-18, 3.292622e-18, 3.288744e-18, 
    3.295881e-18, 3.297311e-18, 3.286477e-18, 3.293113e-18, 3.271806e-18, 
    3.275228e-18, 3.2732e-18, 3.265732e-18, 3.289619e-18, 3.277335e-18, 
    3.300059e-18, 3.293387e-18, 3.312892e-18, 3.303167e-18, 3.322273e-18, 
    3.330431e-18, 3.338487e-18, 3.347855e-18, 3.27134e-18, 3.26875e-18, 
    3.2734e-18, 3.279818e-18, 3.28582e-18, 3.293791e-18, 3.294614e-18, 
    3.296106e-18, 3.299987e-18, 3.303247e-18, 3.296565e-18, 3.304066e-18, 
    3.275995e-18, 3.290693e-18, 3.267759e-18, 3.274634e-18, 3.279446e-18, 
    3.277347e-18, 3.288304e-18, 3.290886e-18, 3.301389e-18, 3.295964e-18, 
    3.328405e-18, 3.314021e-18, 3.355043e-18, 3.343348e-18, 3.267842e-18, 
    3.271337e-18, 3.283504e-18, 3.277713e-18, 3.29433e-18, 3.298425e-18, 
    3.301768e-18, 3.306023e-18, 3.306492e-18, 3.309017e-18, 3.304879e-18, 
    3.308859e-18, 3.293808e-18, 3.300529e-18, 3.282128e-18, 3.286591e-18, 
    3.284542e-18, 3.282285e-18, 3.289252e-18, 3.296666e-18, 3.296846e-18, 
    3.299222e-18, 3.305889e-18, 3.294398e-18, 3.330225e-18, 3.308028e-18, 
    3.27515e-18, 3.281868e-18, 3.282853e-18, 3.280245e-18, 3.298013e-18, 
    3.291564e-18, 3.308959e-18, 3.304255e-18, 3.31197e-18, 3.308133e-18, 
    3.307567e-18, 3.30265e-18, 3.299585e-18, 3.291855e-18, 3.285583e-18, 
    3.280626e-18, 3.28178e-18, 3.287227e-18, 3.297125e-18, 3.306525e-18, 
    3.304461e-18, 3.311383e-18, 3.293122e-18, 3.300759e-18, 3.297799e-18, 
    3.305526e-18, 3.288636e-18, 3.302951e-18, 3.284978e-18, 3.286555e-18, 
    3.291436e-18, 3.301264e-18, 3.303472e-18, 3.305794e-18, 3.304365e-18, 
    3.297381e-18, 3.296247e-18, 3.291323e-18, 3.289954e-18, 3.286213e-18, 
    3.283109e-18, 3.28594e-18, 3.28891e-18, 3.297392e-18, 3.305039e-18, 
    3.313398e-18, 3.315455e-18, 3.325193e-18, 3.317235e-18, 3.330345e-18, 
    3.319152e-18, 3.338887e-18, 3.303813e-18, 3.318867e-18, 3.291666e-18, 
    3.294593e-18, 3.29987e-18, 3.312044e-18, 3.30549e-18, 3.313166e-18, 
    3.296204e-18, 3.287404e-18, 3.285157e-18, 3.280923e-18, 3.285253e-18, 
    3.284902e-18, 3.289048e-18, 3.287717e-18, 3.297675e-18, 3.292324e-18, 
    3.307548e-18, 3.313111e-18, 3.328884e-18, 3.338886e-18, 3.349196e-18, 
    3.353743e-18, 3.355129e-18, 3.355707e-18,
  1.373188e-22, 1.378299e-22, 1.377306e-22, 1.381604e-22, 1.379149e-22, 
    1.382049e-22, 1.374227e-22, 1.378498e-22, 1.375773e-22, 1.373653e-22, 
    1.39022e-22, 1.381803e-22, 1.399152e-22, 1.393642e-22, 1.407688e-22, 
    1.398272e-22, 1.409594e-22, 1.407425e-22, 1.413986e-22, 1.412104e-22, 
    1.420501e-22, 1.414855e-22, 1.424886e-22, 1.419157e-22, 1.420048e-22, 
    1.414667e-22, 1.383502e-22, 1.389167e-22, 1.383165e-22, 1.383972e-22, 
    1.383612e-22, 1.379197e-22, 1.377114e-22, 1.372805e-22, 1.373588e-22, 
    1.376757e-22, 1.384335e-22, 1.381707e-22, 1.388358e-22, 1.388208e-22, 
    1.395637e-22, 1.392283e-22, 1.405146e-22, 1.401439e-22, 1.412183e-22, 
    1.409473e-22, 1.412054e-22, 1.411272e-22, 1.412064e-22, 1.408092e-22, 
    1.409792e-22, 1.406304e-22, 1.392908e-22, 1.396739e-22, 1.385362e-22, 
    1.378589e-22, 1.374412e-22, 1.371448e-22, 1.371867e-22, 1.372664e-22, 
    1.376775e-22, 1.380774e-22, 1.383954e-22, 1.386084e-22, 1.388186e-22, 
    1.394541e-22, 1.397995e-22, 1.405893e-22, 1.404473e-22, 1.406885e-22, 
    1.409204e-22, 1.413094e-22, 1.412454e-22, 1.414168e-22, 1.406827e-22, 
    1.4117e-22, 1.403663e-22, 1.405856e-22, 1.388725e-22, 1.382417e-22, 
    1.379715e-22, 1.377496e-22, 1.372188e-22, 1.37585e-22, 1.374404e-22, 
    1.377852e-22, 1.380111e-22, 1.378959e-22, 1.386142e-22, 1.383341e-22, 
    1.398204e-22, 1.391747e-22, 1.408934e-22, 1.404765e-22, 1.409936e-22, 
    1.407297e-22, 1.411818e-22, 1.407749e-22, 1.414809e-22, 1.416346e-22, 
    1.415295e-22, 1.419349e-22, 1.407522e-22, 1.412051e-22, 1.378927e-22, 
    1.379104e-22, 1.37999e-22, 1.376305e-22, 1.376085e-22, 1.372782e-22, 
    1.375724e-22, 1.376976e-22, 1.380249e-22, 1.382275e-22, 1.384205e-22, 
    1.388456e-22, 1.393212e-22, 1.400029e-22, 1.405034e-22, 1.408396e-22, 
    1.406336e-22, 1.408154e-22, 1.406121e-22, 1.40517e-22, 1.415768e-22, 
    1.409806e-22, 1.418765e-22, 1.418269e-22, 1.414208e-22, 1.418325e-22, 
    1.379238e-22, 1.378213e-22, 1.374684e-22, 1.377445e-22, 1.372423e-22, 
    1.375228e-22, 1.376841e-22, 1.383392e-22, 1.384879e-22, 1.386249e-22, 
    1.388965e-22, 1.392454e-22, 1.398674e-22, 1.40424e-22, 1.409341e-22, 
    1.408967e-22, 1.409098e-22, 1.410236e-22, 1.407414e-22, 1.4107e-22, 
    1.411249e-22, 1.409809e-22, 1.418203e-22, 1.415801e-22, 1.418259e-22, 
    1.416695e-22, 1.378544e-22, 1.380338e-22, 1.379346e-22, 1.381211e-22, 
    1.379894e-22, 1.385748e-22, 1.387507e-22, 1.395772e-22, 1.392384e-22, 
    1.397844e-22, 1.392934e-22, 1.393792e-22, 1.398013e-22, 1.393199e-22, 
    1.403926e-22, 1.396552e-22, 1.410281e-22, 1.402877e-22, 1.410745e-22, 
    1.409319e-22, 1.411684e-22, 1.413801e-22, 1.416475e-22, 1.421409e-22, 
    1.420267e-22, 1.424407e-22, 1.383081e-22, 1.385466e-22, 1.385262e-22, 
    1.387765e-22, 1.389617e-22, 1.393647e-22, 1.400266e-22, 1.397737e-22, 
    1.402389e-22, 1.403322e-22, 1.396264e-22, 1.400587e-22, 1.387068e-22, 
    1.389214e-22, 1.387941e-22, 1.383266e-22, 1.398311e-22, 1.390534e-22, 
    1.405116e-22, 1.400763e-22, 1.413499e-22, 1.407147e-22, 1.419637e-22, 
    1.424987e-22, 1.430151e-22, 1.436173e-22, 1.386775e-22, 1.385153e-22, 
    1.388065e-22, 1.392091e-22, 1.395853e-22, 1.401027e-22, 1.401563e-22, 
    1.402536e-22, 1.405068e-22, 1.407196e-22, 1.402838e-22, 1.40773e-22, 
    1.389699e-22, 1.39901e-22, 1.384534e-22, 1.388842e-22, 1.391856e-22, 
    1.39054e-22, 1.39745e-22, 1.399133e-22, 1.405985e-22, 1.402443e-22, 
    1.423659e-22, 1.41424e-22, 1.440792e-22, 1.433277e-22, 1.384585e-22, 
    1.386773e-22, 1.394401e-22, 1.390768e-22, 1.401378e-22, 1.404049e-22, 
    1.40623e-22, 1.40901e-22, 1.409315e-22, 1.410966e-22, 1.408261e-22, 
    1.410861e-22, 1.401038e-22, 1.405422e-22, 1.393535e-22, 1.396337e-22, 
    1.395049e-22, 1.393634e-22, 1.398068e-22, 1.402905e-22, 1.403019e-22, 
    1.404571e-22, 1.408935e-22, 1.401422e-22, 1.42486e-22, 1.410331e-22, 
    1.389161e-22, 1.393376e-22, 1.393991e-22, 1.392355e-22, 1.403781e-22, 
    1.399576e-22, 1.410927e-22, 1.407854e-22, 1.412895e-22, 1.410387e-22, 
    1.410018e-22, 1.406806e-22, 1.404806e-22, 1.399766e-22, 1.395704e-22, 
    1.392593e-22, 1.393317e-22, 1.39675e-22, 1.403204e-22, 1.409338e-22, 
    1.407991e-22, 1.412511e-22, 1.400591e-22, 1.405574e-22, 1.403643e-22, 
    1.408684e-22, 1.397668e-22, 1.407014e-22, 1.395323e-22, 1.396313e-22, 
    1.399492e-22, 1.405906e-22, 1.407343e-22, 1.408861e-22, 1.407926e-22, 
    1.40337e-22, 1.402629e-22, 1.399417e-22, 1.398527e-22, 1.396098e-22, 
    1.39415e-22, 1.395927e-22, 1.397847e-22, 1.403376e-22, 1.408368e-22, 
    1.41383e-22, 1.415173e-22, 1.421557e-22, 1.416345e-22, 1.424939e-22, 
    1.417609e-22, 1.430418e-22, 1.407572e-22, 1.417414e-22, 1.39964e-22, 
    1.401549e-22, 1.404996e-22, 1.412948e-22, 1.408661e-22, 1.413681e-22, 
    1.402601e-22, 1.396868e-22, 1.395435e-22, 1.39278e-22, 1.395496e-22, 
    1.395276e-22, 1.397935e-22, 1.397067e-22, 1.40356e-22, 1.40007e-22, 
    1.410006e-22, 1.413644e-22, 1.423969e-22, 1.430412e-22, 1.43703e-22, 
    1.439954e-22, 1.440846e-22, 1.441218e-22,
  1.884578e-27, 1.894281e-27, 1.892394e-27, 1.900461e-27, 1.895894e-27, 
    1.901288e-27, 1.886547e-27, 1.894662e-27, 1.889481e-27, 1.885457e-27, 
    1.916515e-27, 1.90083e-27, 1.933211e-27, 1.922885e-27, 1.949276e-27, 
    1.931558e-27, 1.952868e-27, 1.948777e-27, 1.961147e-27, 1.957597e-27, 
    1.973463e-27, 1.962787e-27, 1.981753e-27, 1.970917e-27, 1.972603e-27, 
    1.962434e-27, 1.903991e-27, 1.914552e-27, 1.903363e-27, 1.904867e-27, 
    1.904195e-27, 1.895983e-27, 1.892034e-27, 1.883847e-27, 1.885333e-27, 
    1.891353e-27, 1.905543e-27, 1.90065e-27, 1.913031e-27, 1.912751e-27, 
    1.926608e-27, 1.920349e-27, 1.944485e-27, 1.937505e-27, 1.957746e-27, 
    1.952636e-27, 1.957503e-27, 1.956028e-27, 1.957522e-27, 1.950034e-27, 
    1.953239e-27, 1.946665e-27, 1.921517e-27, 1.928672e-27, 1.907454e-27, 
    1.89484e-27, 1.8869e-27, 1.881292e-27, 1.882069e-27, 1.883581e-27, 
    1.891388e-27, 1.898914e-27, 1.90483e-27, 1.908795e-27, 1.91271e-27, 
    1.924571e-27, 1.931035e-27, 1.945892e-27, 1.943216e-27, 1.947761e-27, 
    1.952129e-27, 1.959465e-27, 1.958258e-27, 1.961493e-27, 1.94765e-27, 
    1.956836e-27, 1.941689e-27, 1.945821e-27, 1.91373e-27, 1.901971e-27, 
    1.896953e-27, 1.892755e-27, 1.882679e-27, 1.889629e-27, 1.886885e-27, 
    1.893429e-27, 1.897681e-27, 1.895534e-27, 1.908903e-27, 1.903689e-27, 
    1.931428e-27, 1.919353e-27, 1.951619e-27, 1.943766e-27, 1.953508e-27, 
    1.948534e-27, 1.957059e-27, 1.949385e-27, 1.962702e-27, 1.965607e-27, 
    1.963621e-27, 1.971276e-27, 1.948959e-27, 1.957498e-27, 1.895474e-27, 
    1.89581e-27, 1.897455e-27, 1.890494e-27, 1.890076e-27, 1.883804e-27, 
    1.889388e-27, 1.891767e-27, 1.897938e-27, 1.901706e-27, 1.905298e-27, 
    1.913216e-27, 1.922086e-27, 1.934857e-27, 1.944273e-27, 1.950605e-27, 
    1.946724e-27, 1.95015e-27, 1.946318e-27, 1.944527e-27, 1.964515e-27, 
    1.953266e-27, 1.970174e-27, 1.969236e-27, 1.961568e-27, 1.969342e-27, 
    1.896058e-27, 1.894116e-27, 1.887415e-27, 1.892657e-27, 1.883123e-27, 
    1.888448e-27, 1.891513e-27, 1.903788e-27, 1.906552e-27, 1.909104e-27, 
    1.914163e-27, 1.920669e-27, 1.93231e-27, 1.942779e-27, 1.952385e-27, 
    1.951681e-27, 1.951929e-27, 1.954075e-27, 1.948756e-27, 1.95495e-27, 
    1.955987e-27, 1.95327e-27, 1.969111e-27, 1.964574e-27, 1.969217e-27, 
    1.966263e-27, 1.894744e-27, 1.898104e-27, 1.896259e-27, 1.899728e-27, 
    1.89728e-27, 1.908174e-27, 1.911451e-27, 1.926866e-27, 1.920538e-27, 
    1.930749e-27, 1.921565e-27, 1.923166e-27, 1.931074e-27, 1.922057e-27, 
    1.942191e-27, 1.928325e-27, 1.954158e-27, 1.940219e-27, 1.955034e-27, 
    1.952344e-27, 1.956804e-27, 1.960801e-27, 1.965848e-27, 1.975175e-27, 
    1.973014e-27, 1.980844e-27, 1.903206e-27, 1.907647e-27, 1.907264e-27, 
    1.911927e-27, 1.91538e-27, 1.922894e-27, 1.935301e-27, 1.930545e-27, 
    1.939293e-27, 1.94105e-27, 1.927777e-27, 1.935905e-27, 1.910631e-27, 
    1.914631e-27, 1.912255e-27, 1.903551e-27, 1.931628e-27, 1.917092e-27, 
    1.944428e-27, 1.936236e-27, 1.960229e-27, 1.948256e-27, 1.971823e-27, 
    1.981948e-27, 1.991684e-27, 2.00333e-27, 1.910084e-27, 1.907061e-27, 
    1.912485e-27, 1.919995e-27, 1.927012e-27, 1.936733e-27, 1.937739e-27, 
    1.939571e-27, 1.944335e-27, 1.948344e-27, 1.940142e-27, 1.94935e-27, 
    1.915543e-27, 1.93294e-27, 1.905911e-27, 1.91394e-27, 1.919555e-27, 
    1.917099e-27, 1.930004e-27, 1.933168e-27, 1.946066e-27, 1.939395e-27, 
    1.979437e-27, 1.961633e-27, 2.012266e-27, 1.997727e-27, 1.906004e-27, 
    1.910078e-27, 1.924304e-27, 1.917525e-27, 1.937391e-27, 1.942419e-27, 
    1.946523e-27, 1.951765e-27, 1.952338e-27, 1.955451e-27, 1.950351e-27, 
    1.955253e-27, 1.936754e-27, 1.945003e-27, 1.922684e-27, 1.927915e-27, 
    1.92551e-27, 1.922868e-27, 1.931166e-27, 1.940269e-27, 1.940478e-27, 
    1.943403e-27, 1.951639e-27, 1.937474e-27, 1.981718e-27, 1.954268e-27, 
    1.914528e-27, 1.922394e-27, 1.923537e-27, 1.920482e-27, 1.941914e-27, 
    1.934002e-27, 1.955378e-27, 1.949583e-27, 1.959088e-27, 1.954359e-27, 
    1.953663e-27, 1.947609e-27, 1.943844e-27, 1.934361e-27, 1.926735e-27, 
    1.920927e-27, 1.922277e-27, 1.928693e-27, 1.94083e-27, 1.952383e-27, 
    1.949846e-27, 1.958365e-27, 1.93591e-27, 1.945291e-27, 1.941656e-27, 
    1.951149e-27, 1.930416e-27, 1.948017e-27, 1.92602e-27, 1.927869e-27, 
    1.933846e-27, 1.94592e-27, 1.948621e-27, 1.951483e-27, 1.949719e-27, 
    1.941142e-27, 1.939746e-27, 1.933703e-27, 1.932031e-27, 1.927467e-27, 
    1.923832e-27, 1.92715e-27, 1.930755e-27, 1.941152e-27, 1.950554e-27, 
    1.960856e-27, 1.963389e-27, 1.975461e-27, 1.96561e-27, 1.981869e-27, 
    1.968008e-27, 1.992214e-27, 1.949062e-27, 1.967631e-27, 1.934123e-27, 
    1.937712e-27, 1.944204e-27, 1.959196e-27, 1.951105e-27, 1.960577e-27, 
    1.939693e-27, 1.928916e-27, 1.926231e-27, 1.921277e-27, 1.926344e-27, 
    1.925932e-27, 1.930916e-27, 1.929285e-27, 1.941498e-27, 1.93493e-27, 
    1.953642e-27, 1.960505e-27, 1.980017e-27, 1.992192e-27, 2.004981e-27, 
    2.01064e-27, 2.012367e-27, 2.013088e-27,
  8.306839e-33, 8.364191e-33, 8.353025e-33, 8.400282e-33, 8.373716e-33, 
    8.405094e-33, 8.318461e-33, 8.366452e-33, 8.3358e-33, 8.312022e-33, 
    8.494805e-33, 8.402431e-33, 8.594389e-33, 8.532886e-33, 8.689637e-33, 
    8.584615e-33, 8.710969e-33, 8.686652e-33, 8.760185e-33, 8.739064e-33, 
    8.83362e-33, 8.76995e-33, 8.883112e-33, 8.818409e-33, 8.828478e-33, 
    8.767847e-33, 8.420812e-33, 8.48306e-33, 8.417163e-33, 8.425919e-33, 
    8.422003e-33, 8.374243e-33, 8.350915e-33, 8.302511e-33, 8.311289e-33, 
    8.346872e-33, 8.429861e-33, 8.401366e-33, 8.473895e-33, 8.472221e-33, 
    8.5552e-33, 8.517689e-33, 8.66118e-33, 8.619795e-33, 8.739946e-33, 
    8.709573e-33, 8.738506e-33, 8.729732e-33, 8.738621e-33, 8.694119e-33, 
    8.713156e-33, 8.674113e-33, 8.524691e-33, 8.567524e-33, 8.440984e-33, 
    8.367525e-33, 8.32055e-33, 8.287453e-33, 8.292016e-33, 8.30095e-33, 
    8.34708e-33, 8.39127e-33, 8.425692e-33, 8.448784e-33, 8.471978e-33, 
    8.543025e-33, 8.581514e-33, 8.669541e-33, 8.653645e-33, 8.680631e-33, 
    8.70656e-33, 8.750184e-33, 8.742997e-33, 8.762255e-33, 8.679955e-33, 
    8.734552e-33, 8.64459e-33, 8.669102e-33, 8.478147e-33, 8.409054e-33, 
    8.3799e-33, 8.355163e-33, 8.295619e-33, 8.336684e-33, 8.320467e-33, 
    8.35914e-33, 8.384102e-33, 8.37159e-33, 8.449417e-33, 8.419052e-33, 
    8.583836e-33, 8.511736e-33, 8.703532e-33, 8.65691e-33, 8.714749e-33, 
    8.6852e-33, 8.735871e-33, 8.690256e-33, 8.769449e-33, 8.786758e-33, 
    8.774921e-33, 8.820542e-33, 8.687728e-33, 8.738486e-33, 8.37124e-33, 
    8.373227e-33, 8.382788e-33, 8.341796e-33, 8.339323e-33, 8.302261e-33, 
    8.335249e-33, 8.349319e-33, 8.385592e-33, 8.407515e-33, 8.428419e-33, 
    8.475009e-33, 8.528109e-33, 8.604127e-33, 8.659922e-33, 8.697503e-33, 
    8.674455e-33, 8.694799e-33, 8.672052e-33, 8.661418e-33, 8.780254e-33, 
    8.713322e-33, 8.813966e-33, 8.808376e-33, 8.762705e-33, 8.809006e-33, 
    8.374668e-33, 8.363198e-33, 8.32359e-33, 8.354572e-33, 8.298237e-33, 
    8.329699e-33, 8.347828e-33, 8.419641e-33, 8.435718e-33, 8.450589e-33, 
    8.48067e-33, 8.519604e-33, 8.589043e-33, 8.651065e-33, 8.708079e-33, 
    8.703894e-33, 8.705365e-33, 8.718124e-33, 8.686522e-33, 8.723325e-33, 
    8.729496e-33, 8.713339e-33, 8.807627e-33, 8.780595e-33, 8.808257e-33, 
    8.790652e-33, 8.366915e-33, 8.386563e-33, 8.375834e-33, 8.39601e-33, 
    8.381775e-33, 8.445189e-33, 8.464481e-33, 8.556762e-33, 8.518824e-33, 
    8.579808e-33, 8.524969e-33, 8.534567e-33, 8.581761e-33, 8.527912e-33, 
    8.647595e-33, 8.565492e-33, 8.718621e-33, 8.63592e-33, 8.723823e-33, 
    8.707831e-33, 8.734345e-33, 8.758131e-33, 8.78818e-33, 8.843819e-33, 
    8.830914e-33, 8.877665e-33, 8.416241e-33, 8.442109e-33, 8.439867e-33, 
    8.467298e-33, 8.487951e-33, 8.532928e-33, 8.606743e-33, 8.578588e-33, 
    8.630385e-33, 8.640806e-33, 8.562197e-33, 8.610332e-33, 8.459562e-33, 
    8.483494e-33, 8.469265e-33, 8.418257e-33, 8.585015e-33, 8.498215e-33, 
    8.66084e-33, 8.612279e-33, 8.754731e-33, 8.683573e-33, 8.823809e-33, 
    8.884297e-33, 8.942317e-33, 9.012262e-33, 8.456301e-33, 8.438684e-33, 
    8.470628e-33, 8.515587e-33, 8.557615e-33, 8.615226e-33, 8.62118e-33, 
    8.632041e-33, 8.660281e-33, 8.684073e-33, 8.63544e-33, 8.690051e-33, 
    8.488976e-33, 8.592776e-33, 8.431997e-33, 8.479362e-33, 8.512948e-33, 
    8.498238e-33, 8.575386e-33, 8.594108e-33, 8.67057e-33, 8.630987e-33, 
    8.869297e-33, 8.763108e-33, 9.06672e-33, 8.978599e-33, 8.432527e-33, 
    8.456258e-33, 8.541395e-33, 8.500784e-33, 8.619117e-33, 8.648925e-33, 
    8.673262e-33, 8.704402e-33, 8.707798e-33, 8.72631e-33, 8.695991e-33, 
    8.725126e-33, 8.615349e-33, 8.664251e-33, 8.531666e-33, 8.563035e-33, 
    8.548604e-33, 8.532772e-33, 8.582261e-33, 8.636194e-33, 8.637412e-33, 
    8.654764e-33, 8.703725e-33, 8.619608e-33, 8.882973e-33, 8.719342e-33, 
    8.482848e-33, 8.529962e-33, 8.536786e-33, 8.518479e-33, 8.645931e-33, 
    8.599052e-33, 8.725867e-33, 8.691436e-33, 8.747935e-33, 8.71981e-33, 
    8.715677e-33, 8.679711e-33, 8.657372e-33, 8.601185e-33, 8.555957e-33, 
    8.521139e-33, 8.529228e-33, 8.567641e-33, 8.639518e-33, 8.708078e-33, 
    8.693008e-33, 8.74363e-33, 8.610347e-33, 8.665969e-33, 8.644411e-33, 
    8.70074e-33, 8.577827e-33, 8.682202e-33, 8.551663e-33, 8.562748e-33, 
    8.598125e-33, 8.669712e-33, 8.685719e-33, 8.702727e-33, 8.692241e-33, 
    8.641361e-33, 8.63308e-33, 8.597278e-33, 8.587387e-33, 8.560339e-33, 
    8.538546e-33, 8.558439e-33, 8.579839e-33, 8.641409e-33, 8.697212e-33, 
    8.758461e-33, 8.773535e-33, 8.845564e-33, 8.786801e-33, 8.883879e-33, 
    8.80115e-33, 8.94556e-33, 8.688378e-33, 8.798856e-33, 8.599759e-33, 
    8.621019e-33, 8.65953e-33, 8.748603e-33, 8.700476e-33, 8.756815e-33, 
    8.632761e-33, 8.568973e-33, 8.552927e-33, 8.523241e-33, 8.553607e-33, 
    8.551136e-33, 8.580777e-33, 8.571128e-33, 8.643461e-33, 8.604539e-33, 
    8.715557e-33, 8.756385e-33, 8.872732e-33, 8.945393e-33, 9.022153e-33, 
    9.056702e-33, 9.067332e-33, 9.071776e-33,
  1.197076e-38, 1.208709e-38, 1.20644e-38, 1.21598e-38, 1.210643e-38, 
    1.216947e-38, 1.199428e-38, 1.20917e-38, 1.202943e-38, 1.198123e-38, 
    1.235082e-38, 1.216412e-38, 1.255302e-38, 1.24282e-38, 1.275007e-38, 
    1.253329e-38, 1.279456e-38, 1.27438e-38, 1.289748e-38, 1.285324e-38, 
    1.305196e-38, 1.291796e-38, 1.315653e-38, 1.301986e-38, 1.30411e-38, 
    1.291355e-38, 1.220107e-38, 1.232697e-38, 1.219373e-38, 1.221137e-38, 
    1.220347e-38, 1.21075e-38, 1.206015e-38, 1.196197e-38, 1.197975e-38, 
    1.205191e-38, 1.221931e-38, 1.216195e-38, 1.230825e-38, 1.230486e-38, 
    1.24737e-38, 1.239725e-38, 1.269078e-38, 1.260485e-38, 1.285509e-38, 
    1.279161e-38, 1.285208e-38, 1.283372e-38, 1.285232e-38, 1.275937e-38, 
    1.27991e-38, 1.271768e-38, 1.241151e-38, 1.249876e-38, 1.224172e-38, 
    1.209392e-38, 1.199852e-38, 1.193144e-38, 1.194075e-38, 1.195883e-38, 
    1.205234e-38, 1.214166e-38, 1.221089e-38, 1.225743e-38, 1.230437e-38, 
    1.244893e-38, 1.252701e-38, 1.27082e-38, 1.267511e-38, 1.273128e-38, 
    1.278532e-38, 1.287653e-38, 1.286148e-38, 1.290183e-38, 1.272985e-38, 
    1.284383e-38, 1.265628e-38, 1.270725e-38, 1.231701e-38, 1.217741e-38, 
    1.211889e-38, 1.206874e-38, 1.194804e-38, 1.203123e-38, 1.199835e-38, 
    1.20768e-38, 1.212727e-38, 1.210211e-38, 1.22587e-38, 1.219752e-38, 
    1.25317e-38, 1.238516e-38, 1.2779e-38, 1.26819e-38, 1.280241e-38, 
    1.274077e-38, 1.284658e-38, 1.27513e-38, 1.291691e-38, 1.295327e-38, 
    1.292841e-38, 1.302433e-38, 1.274604e-38, 1.285205e-38, 1.21014e-38, 
    1.210545e-38, 1.212463e-38, 1.204161e-38, 1.203659e-38, 1.196147e-38, 
    1.202831e-38, 1.205687e-38, 1.213025e-38, 1.217432e-38, 1.221639e-38, 
    1.231053e-38, 1.241849e-38, 1.257268e-38, 1.268816e-38, 1.276641e-38, 
    1.271838e-38, 1.276077e-38, 1.271339e-38, 1.269126e-38, 1.293962e-38, 
    1.279945e-38, 1.301048e-38, 1.299871e-38, 1.290278e-38, 1.300003e-38, 
    1.210834e-38, 1.208505e-38, 1.200467e-38, 1.206752e-38, 1.195333e-38, 
    1.201706e-38, 1.205386e-38, 1.219874e-38, 1.223109e-38, 1.226108e-38, 
    1.232201e-38, 1.240115e-38, 1.254219e-38, 1.266976e-38, 1.278848e-38, 
    1.277974e-38, 1.278282e-38, 1.280947e-38, 1.274353e-38, 1.282033e-38, 
    1.283325e-38, 1.279947e-38, 1.299713e-38, 1.29403e-38, 1.299846e-38, 
    1.296143e-38, 1.20926e-38, 1.213221e-38, 1.211067e-38, 1.215119e-38, 
    1.212261e-38, 1.225021e-38, 1.228921e-38, 1.247692e-38, 1.239957e-38, 
    1.252355e-38, 1.241207e-38, 1.243163e-38, 1.252755e-38, 1.241805e-38, 
    1.266258e-38, 1.24947e-38, 1.281051e-38, 1.263837e-38, 1.282137e-38, 
    1.278796e-38, 1.284336e-38, 1.289319e-38, 1.295624e-38, 1.307344e-38, 
    1.30462e-38, 1.314498e-38, 1.219187e-38, 1.224399e-38, 1.223944e-38, 
    1.229488e-38, 1.23368e-38, 1.242827e-38, 1.257796e-38, 1.252106e-38, 
    1.262681e-38, 1.264844e-38, 1.248796e-38, 1.258527e-38, 1.227921e-38, 
    1.232778e-38, 1.229888e-38, 1.219594e-38, 1.253407e-38, 1.235768e-38, 
    1.269007e-38, 1.258928e-38, 1.288606e-38, 1.273742e-38, 1.303122e-38, 
    1.315908e-38, 1.328167e-38, 1.343035e-38, 1.22726e-38, 1.223706e-38, 
    1.230163e-38, 1.2393e-38, 1.247862e-38, 1.259539e-38, 1.260772e-38, 
    1.263025e-38, 1.26889e-38, 1.273842e-38, 1.263733e-38, 1.275087e-38, 
    1.233897e-38, 1.254973e-38, 1.22236e-38, 1.23194e-38, 1.238762e-38, 
    1.23577e-38, 1.251459e-38, 1.25524e-38, 1.271033e-38, 1.262805e-38, 
    1.312734e-38, 1.290366e-38, 1.354838e-38, 1.335797e-38, 1.222465e-38, 
    1.22725e-38, 1.244555e-38, 1.236287e-38, 1.260344e-38, 1.266531e-38, 
    1.27159e-38, 1.278083e-38, 1.27879e-38, 1.282658e-38, 1.276326e-38, 
    1.282409e-38, 1.259565e-38, 1.269716e-38, 1.242569e-38, 1.248969e-38, 
    1.246022e-38, 1.242795e-38, 1.252847e-38, 1.26389e-38, 1.264139e-38, 
    1.267745e-38, 1.277956e-38, 1.260446e-38, 1.315637e-38, 1.281214e-38, 
    1.232642e-38, 1.242227e-38, 1.243614e-38, 1.239884e-38, 1.265909e-38, 
    1.25624e-38, 1.282565e-38, 1.275376e-38, 1.287181e-38, 1.281299e-38, 
    1.280435e-38, 1.272933e-38, 1.268286e-38, 1.256672e-38, 1.247524e-38, 
    1.240426e-38, 1.242073e-38, 1.249899e-38, 1.264579e-38, 1.27885e-38, 
    1.275707e-38, 1.28628e-38, 1.258527e-38, 1.270075e-38, 1.265595e-38, 
    1.277317e-38, 1.251953e-38, 1.273466e-38, 1.246646e-38, 1.248909e-38, 
    1.256053e-38, 1.270857e-38, 1.274185e-38, 1.277733e-38, 1.275544e-38, 
    1.264961e-38, 1.263241e-38, 1.255881e-38, 1.253884e-38, 1.248417e-38, 
    1.243971e-38, 1.24803e-38, 1.252361e-38, 1.264969e-38, 1.276583e-38, 
    1.289388e-38, 1.292548e-38, 1.30772e-38, 1.295342e-38, 1.31583e-38, 
    1.298368e-38, 1.32886e-38, 1.274747e-38, 1.297877e-38, 1.256382e-38, 
    1.260738e-38, 1.268738e-38, 1.287327e-38, 1.277262e-38, 1.289046e-38, 
    1.263175e-38, 1.25017e-38, 1.246904e-38, 1.240854e-38, 1.247043e-38, 
    1.246539e-38, 1.252547e-38, 1.2506e-38, 1.265395e-38, 1.257348e-38, 
    1.280411e-38, 1.288955e-38, 1.313455e-38, 1.328818e-38, 1.345166e-38, 
    1.352658e-38, 1.354968e-38, 1.355935e-38,
  7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  8.734524e-06, 8.571744e-06, 8.603407e-06, 8.472e-06, 8.544916e-06, 
    8.458845e-06, 8.701544e-06, 8.565271e-06, 8.652284e-06, 8.719888e-06, 
    8.216618e-06, 8.466137e-06, 7.957028e-06, 8.116502e-06, 7.715558e-06, 
    7.981846e-06, 7.661804e-06, 7.723266e-06, 7.538236e-06, 7.591272e-06, 
    7.354279e-06, 7.513751e-06, 7.231284e-06, 7.392392e-06, 7.367194e-06, 
    7.519006e-06, 8.415975e-06, 8.247702e-06, 8.425935e-06, 8.401954e-06, 
    8.412719e-06, 8.543404e-06, 8.609205e-06, 8.74697e-06, 8.721971e-06, 
    8.620789e-06, 8.39117e-06, 8.469168e-06, 8.272545e-06, 8.276988e-06, 
    8.057758e-06, 8.156647e-06, 7.787655e-06, 7.892636e-06, 7.589059e-06, 
    7.665469e-06, 7.592646e-06, 7.614734e-06, 7.592358e-06, 7.704404e-06, 
    7.656409e-06, 7.754966e-06, 8.138129e-06, 8.025627e-06, 8.360882e-06, 
    8.562058e-06, 8.695567e-06, 8.790221e-06, 8.776843e-06, 8.751334e-06, 
    8.620197e-06, 8.496809e-06, 8.402701e-06, 8.339714e-06, 8.277627e-06, 
    8.089478e-06, 7.989829e-06, 7.766408e-06, 7.806771e-06, 7.738398e-06, 
    7.673068e-06, 7.56329e-06, 7.581368e-06, 7.532976e-06, 7.740214e-06, 
    7.602514e-06, 7.829753e-06, 7.767639e-06, 8.260684e-06, 8.448133e-06, 
    8.527682e-06, 8.597319e-06, 8.766556e-06, 8.649702e-06, 8.695776e-06, 
    8.586151e-06, 8.516442e-06, 8.550925e-06, 8.337992e-06, 8.42081e-06, 
    7.98392e-06, 8.172274e-06, 7.68069e-06, 7.79849e-06, 7.652441e-06, 
    7.72699e-06, 7.599224e-06, 7.714218e-06, 7.514966e-06, 7.471532e-06, 
    7.501214e-06, 7.387178e-06, 7.720588e-06, 7.59264e-06, 8.55189e-06, 
    8.546265e-06, 8.520069e-06, 8.635185e-06, 8.642227e-06, 8.747653e-06, 
    8.653854e-06, 8.613888e-06, 8.512405e-06, 8.452334e-06, 8.39521e-06, 
    8.269532e-06, 8.12903e-06, 7.932334e-06, 7.790855e-06, 7.695933e-06, 
    7.754151e-06, 7.702753e-06, 7.760205e-06, 7.787127e-06, 7.487804e-06, 
    7.655957e-06, 7.403587e-06, 7.417566e-06, 7.531823e-06, 7.415991e-06, 
    8.542317e-06, 8.574676e-06, 8.686948e-06, 8.599092e-06, 8.75913e-06, 
    8.669563e-06, 8.618033e-06, 8.419067e-06, 8.375329e-06, 8.334742e-06, 
    8.254562e-06, 8.151587e-06, 7.970754e-06, 7.813226e-06, 7.669269e-06, 
    7.679823e-06, 7.676107e-06, 7.643922e-06, 7.723624e-06, 7.630833e-06, 
    7.615247e-06, 7.655985e-06, 7.419438e-06, 7.487063e-06, 7.417863e-06, 
    7.461901e-06, 8.56416e-06, 8.509706e-06, 8.539133e-06, 8.48379e-06, 
    8.522777e-06, 8.349322e-06, 8.297277e-06, 8.053496e-06, 8.153612e-06, 
    7.99426e-06, 8.137438e-06, 8.112075e-06, 7.989033e-06, 8.129708e-06, 
    7.821905e-06, 8.03064e-06, 7.64267e-06, 7.851369e-06, 7.62958e-06, 
    7.669892e-06, 7.603148e-06, 7.543335e-06, 7.468061e-06, 7.329033e-06, 
    7.361242e-06, 7.244898e-06, 8.428496e-06, 8.357791e-06, 8.364029e-06, 
    8.290009e-06, 8.23524e-06, 8.11647e-06, 7.92575e-06, 7.997503e-06, 
    7.865758e-06, 7.83929e-06, 8.039439e-06, 7.916575e-06, 8.310461e-06, 
    8.246887e-06, 8.28475e-06, 8.422913e-06, 7.980956e-06, 8.207939e-06, 
    7.788514e-06, 7.911702e-06, 7.551864e-06, 7.730929e-06, 7.378967e-06, 
    7.22818e-06, 7.086158e-06, 6.919917e-06, 8.3192e-06, 8.367258e-06, 
    8.281208e-06, 8.162043e-06, 8.051417e-06, 7.904189e-06, 7.889123e-06, 
    7.861517e-06, 7.789997e-06, 7.729828e-06, 7.852776e-06, 7.714742e-06, 
    8.232117e-06, 7.961242e-06, 8.385413e-06, 8.257807e-06, 8.169075e-06, 
    8.208018e-06, 8.005705e-06, 7.957974e-06, 7.763837e-06, 7.864236e-06, 
    7.265402e-06, 7.530682e-06, 6.793232e-06, 6.999745e-06, 8.384043e-06, 
    8.319371e-06, 8.094041e-06, 8.2013e-06, 7.894361e-06, 7.818697e-06, 
    7.757165e-06, 7.678448e-06, 7.669956e-06, 7.623293e-06, 7.699748e-06, 
    7.626318e-06, 7.903875e-06, 7.779914e-06, 8.119829e-06, 8.037167e-06, 
    8.075205e-06, 8.116907e-06, 7.988158e-06, 7.850837e-06, 7.847921e-06, 
    7.803855e-06, 7.679567e-06, 7.893116e-06, 7.231087e-06, 7.640305e-06, 
    8.248815e-06, 8.124074e-06, 8.10627e-06, 8.154607e-06, 7.826284e-06, 
    7.945337e-06, 7.624433e-06, 7.711243e-06, 7.568982e-06, 7.639691e-06, 
    7.65009e-06, 7.740848e-06, 7.797316e-06, 7.939877e-06, 8.055764e-06, 
    8.147599e-06, 8.126252e-06, 8.025355e-06, 7.842438e-06, 7.669178e-06, 
    7.707148e-06, 7.579799e-06, 7.916639e-06, 7.77549e-06, 7.830056e-06, 
    7.687734e-06, 7.999405e-06, 7.733988e-06, 8.067158e-06, 8.037983e-06, 
    7.947699e-06, 7.765898e-06, 7.725672e-06, 7.682672e-06, 7.709211e-06, 
    7.837794e-06, 7.858857e-06, 7.949899e-06, 7.975015e-06, 8.044337e-06, 
    8.101694e-06, 8.049285e-06, 7.994222e-06, 7.837748e-06, 7.69657e-06, 
    7.542481e-06, 7.504752e-06, 7.324381e-06, 7.471204e-06, 7.2288e-06, 
    7.434878e-06, 7.077953e-06, 7.71862e-06, 7.440972e-06, 7.943595e-06, 
    7.889543e-06, 7.791701e-06, 7.567061e-06, 7.688403e-06, 7.546492e-06, 
    7.859684e-06, 8.021862e-06, 8.063815e-06, 8.142015e-06, 8.062027e-06, 
    8.068535e-06, 7.991954e-06, 8.016569e-06, 7.83255e-06, 7.931429e-06, 
    7.650347e-06, 7.547618e-06, 7.257089e-06, 7.078644e-06, 6.896769e-06, 
    6.816381e-06, 6.791905e-06, 6.78167e-06,
  3.492803e-06, 3.360878e-06, 3.386376e-06, 3.281086e-06, 3.339341e-06, 
    3.270622e-06, 3.465909e-06, 3.355673e-06, 3.425893e-06, 3.48086e-06, 
    3.080487e-06, 3.276421e-06, 2.882245e-06, 3.003364e-06, 2.703089e-06, 
    2.900945e-06, 2.663914e-06, 2.708735e-06, 2.574853e-06, 2.612911e-06, 
    2.444837e-06, 2.55737e-06, 2.359677e-06, 2.471521e-06, 2.453866e-06, 
    2.561116e-06, 3.236627e-06, 3.104611e-06, 3.244512e-06, 3.225536e-06, 
    3.23405e-06, 3.338126e-06, 3.391046e-06, 3.502981e-06, 3.48256e-06, 
    3.400405e-06, 3.217018e-06, 3.278838e-06, 3.123976e-06, 3.12744e-06, 
    2.958497e-06, 3.034198e-06, 2.756047e-06, 2.833977e-06, 2.611319e-06, 
    2.666582e-06, 2.6139e-06, 2.62983e-06, 2.613693e-06, 2.694945e-06, 
    2.660001e-06, 2.731982e-06, 3.019957e-06, 2.934079e-06, 3.193152e-06, 
    3.353083e-06, 3.461041e-06, 3.538426e-06, 3.527446e-06, 3.506547e-06, 
    3.399926e-06, 3.300862e-06, 3.226133e-06, 3.17652e-06, 3.127938e-06, 
    2.982673e-06, 2.906976e-06, 2.74039e-06, 2.770166e-06, 2.719817e-06, 
    2.672108e-06, 2.592798e-06, 2.605784e-06, 2.57109e-06, 2.721154e-06, 
    2.621008e-06, 2.787184e-06, 2.7413e-06, 3.114708e-06, 3.262118e-06, 
    3.325521e-06, 3.381467e-06, 3.519012e-06, 3.423796e-06, 3.46121e-06, 
    3.372475e-06, 3.316544e-06, 3.344164e-06, 3.175168e-06, 3.240455e-06, 
    2.902515e-06, 3.046232e-06, 2.677654e-06, 2.764045e-06, 2.657123e-06, 
    2.711463e-06, 2.618637e-06, 2.702118e-06, 2.558234e-06, 2.527347e-06, 
    2.548436e-06, 2.467868e-06, 2.706776e-06, 2.613893e-06, 3.344936e-06, 
    3.340424e-06, 3.319445e-06, 3.412043e-06, 3.417744e-06, 3.503538e-06, 
    3.427165e-06, 3.394833e-06, 3.313319e-06, 3.265454e-06, 3.220213e-06, 
    3.121625e-06, 3.012967e-06, 2.863693e-06, 2.758409e-06, 2.688765e-06, 
    2.731385e-06, 2.693742e-06, 2.735834e-06, 2.755661e-06, 2.538897e-06, 
    2.659672e-06, 2.479386e-06, 2.489221e-06, 2.570265e-06, 2.488112e-06, 
    3.337259e-06, 3.363241e-06, 3.454031e-06, 3.382901e-06, 3.512931e-06, 
    3.439905e-06, 3.398176e-06, 3.239069e-06, 3.204532e-06, 3.172615e-06, 
    3.109971e-06, 3.030304e-06, 2.892588e-06, 2.774937e-06, 2.669346e-06, 
    2.677025e-06, 2.67432e-06, 2.650944e-06, 2.708998e-06, 2.641466e-06, 
    2.630197e-06, 2.659695e-06, 2.490539e-06, 2.538375e-06, 2.48943e-06, 
    2.520527e-06, 3.354789e-06, 3.311161e-06, 3.334707e-06, 3.29048e-06, 
    3.321608e-06, 3.184058e-06, 3.143267e-06, 2.955247e-06, 3.03186e-06, 
    2.910328e-06, 3.019428e-06, 2.999973e-06, 2.906368e-06, 3.013495e-06, 
    2.781357e-06, 2.937874e-06, 2.650038e-06, 2.803214e-06, 2.64056e-06, 
    2.669799e-06, 2.62147e-06, 2.578499e-06, 2.52489e-06, 2.427246e-06, 
    2.449709e-06, 2.369036e-06, 3.246543e-06, 3.190719e-06, 3.195633e-06, 
    3.1376e-06, 3.094952e-06, 3.003343e-06, 2.858756e-06, 2.912786e-06, 
    2.813933e-06, 2.794255e-06, 2.94457e-06, 2.851878e-06, 3.153585e-06, 
    3.103993e-06, 3.133492e-06, 3.242117e-06, 2.900279e-06, 3.073782e-06, 
    2.756681e-06, 2.848232e-06, 2.584606e-06, 2.714341e-06, 2.462111e-06, 
    2.35754e-06, 2.261031e-06, 2.150497e-06, 3.16043e-06, 3.198175e-06, 
    3.130731e-06, 3.038346e-06, 2.953672e-06, 2.84261e-06, 2.831354e-06, 
    2.810774e-06, 2.757778e-06, 2.713542e-06, 2.804267e-06, 2.702501e-06, 
    3.092509e-06, 2.885421e-06, 3.212479e-06, 3.112485e-06, 3.043767e-06, 
    3.073849e-06, 2.918991e-06, 2.882967e-06, 2.7385e-06, 2.812801e-06, 
    2.383151e-06, 2.569444e-06, 2.06808e-06, 2.20324e-06, 3.211402e-06, 
    3.160567e-06, 2.986171e-06, 3.068652e-06, 2.835266e-06, 2.778988e-06, 
    2.7336e-06, 2.676021e-06, 2.669845e-06, 2.636011e-06, 2.691549e-06, 
    2.638201e-06, 2.842375e-06, 2.750341e-06, 3.005919e-06, 2.942841e-06, 
    2.971796e-06, 3.003679e-06, 2.905725e-06, 2.802826e-06, 2.800666e-06, 
    2.768007e-06, 2.67681e-06, 2.834336e-06, 2.359521e-06, 2.6483e-06, 
    3.105502e-06, 3.009163e-06, 2.99553e-06, 3.03263e-06, 2.784608e-06, 
    2.873461e-06, 2.636837e-06, 2.699943e-06, 2.596885e-06, 2.64788e-06, 
    2.655417e-06, 2.721619e-06, 2.763179e-06, 2.869357e-06, 2.956979e-06, 
    3.02724e-06, 3.010845e-06, 2.933874e-06, 2.796587e-06, 2.669276e-06, 
    2.696946e-06, 2.604657e-06, 2.851931e-06, 2.747078e-06, 2.787401e-06, 
    2.682786e-06, 2.914222e-06, 2.716566e-06, 2.965661e-06, 2.943463e-06, 
    2.875236e-06, 2.740012e-06, 2.710497e-06, 2.679096e-06, 2.698459e-06, 
    2.793142e-06, 2.808795e-06, 2.876892e-06, 2.895802e-06, 2.948292e-06, 
    2.992031e-06, 2.952052e-06, 2.910301e-06, 2.793111e-06, 2.689225e-06, 
    2.577887e-06, 2.550957e-06, 2.423999e-06, 2.527106e-06, 2.357949e-06, 
    2.501393e-06, 2.255495e-06, 2.705323e-06, 2.50571e-06, 2.872155e-06, 
    2.831668e-06, 2.759027e-06, 2.595496e-06, 2.683274e-06, 2.580753e-06, 
    2.80941e-06, 2.931221e-06, 2.963113e-06, 3.022946e-06, 2.961751e-06, 
    2.96671e-06, 2.908593e-06, 2.927218e-06, 2.789254e-06, 2.863019e-06, 
    2.655601e-06, 2.581561e-06, 2.377428e-06, 2.25597e-06, 2.135329e-06, 
    2.083025e-06, 2.067227e-06, 2.060638e-06,
  1.618293e-06, 1.550218e-06, 1.563347e-06, 1.509219e-06, 1.539138e-06, 
    1.503852e-06, 1.604386e-06, 1.547539e-06, 1.583721e-06, 1.612116e-06, 
    1.406746e-06, 1.506826e-06, 1.306349e-06, 1.367583e-06, 1.216395e-06, 
    1.315781e-06, 1.196827e-06, 1.219218e-06, 1.15248e-06, 1.171407e-06, 
    1.088095e-06, 1.143797e-06, 1.046158e-06, 1.101274e-06, 1.092552e-06, 
    1.145657e-06, 1.486433e-06, 1.419023e-06, 1.490471e-06, 1.480755e-06, 
    1.485114e-06, 1.538514e-06, 1.565753e-06, 1.62356e-06, 1.612995e-06, 
    1.570577e-06, 1.476397e-06, 1.508066e-06, 1.428887e-06, 1.430653e-06, 
    1.344861e-06, 1.383225e-06, 1.242906e-06, 1.282039e-06, 1.170614e-06, 
    1.198159e-06, 1.171899e-06, 1.179832e-06, 1.171796e-06, 1.212324e-06, 
    1.194874e-06, 1.230851e-06, 1.375998e-06, 1.332514e-06, 1.464192e-06, 
    1.546206e-06, 1.601871e-06, 1.641918e-06, 1.636228e-06, 1.625406e-06, 
    1.57033e-06, 1.519368e-06, 1.481061e-06, 1.455694e-06, 1.430907e-06, 
    1.357099e-06, 1.318825e-06, 1.235061e-06, 1.249986e-06, 1.224762e-06, 
    1.200917e-06, 1.1614e-06, 1.16786e-06, 1.150611e-06, 1.225431e-06, 
    1.175438e-06, 1.258525e-06, 1.235517e-06, 1.424166e-06, 1.499492e-06, 
    1.532034e-06, 1.560818e-06, 1.631859e-06, 1.58264e-06, 1.601958e-06, 
    1.556187e-06, 1.527421e-06, 1.541619e-06, 1.455004e-06, 1.488394e-06, 
    1.316573e-06, 1.389335e-06, 1.203686e-06, 1.246916e-06, 1.193439e-06, 
    1.220582e-06, 1.174258e-06, 1.215909e-06, 1.144227e-06, 1.128905e-06, 
    1.139363e-06, 1.099469e-06, 1.218239e-06, 1.171896e-06, 1.542015e-06, 
    1.539695e-06, 1.528912e-06, 1.576577e-06, 1.579517e-06, 1.623848e-06, 
    1.584378e-06, 1.567705e-06, 1.525765e-06, 1.501203e-06, 1.478031e-06, 
    1.42769e-06, 1.372452e-06, 1.296999e-06, 1.24409e-06, 1.209236e-06, 
    1.230552e-06, 1.211723e-06, 1.23278e-06, 1.242713e-06, 1.134632e-06, 
    1.19471e-06, 1.105162e-06, 1.110026e-06, 1.150201e-06, 1.109478e-06, 
    1.538068e-06, 1.551434e-06, 1.598249e-06, 1.561557e-06, 1.628711e-06, 
    1.590954e-06, 1.569428e-06, 1.487684e-06, 1.47001e-06, 1.4537e-06, 
    1.421753e-06, 1.381248e-06, 1.311564e-06, 1.252379e-06, 1.199538e-06, 
    1.203372e-06, 1.202021e-06, 1.190357e-06, 1.21935e-06, 1.185631e-06, 
    1.180015e-06, 1.194721e-06, 1.110678e-06, 1.134373e-06, 1.11013e-06, 
    1.125525e-06, 1.547084e-06, 1.524656e-06, 1.536756e-06, 1.514038e-06, 
    1.530023e-06, 1.459545e-06, 1.438723e-06, 1.343216e-06, 1.382038e-06, 
    1.320517e-06, 1.375729e-06, 1.365864e-06, 1.318518e-06, 1.37272e-06, 
    1.2556e-06, 1.334432e-06, 1.189905e-06, 1.266574e-06, 1.185179e-06, 
    1.199764e-06, 1.175668e-06, 1.154292e-06, 1.127687e-06, 1.079417e-06, 
    1.0905e-06, 1.050758e-06, 1.491512e-06, 1.462949e-06, 1.46546e-06, 
    1.435833e-06, 1.414106e-06, 1.367572e-06, 1.294512e-06, 1.321758e-06, 
    1.271961e-06, 1.262075e-06, 1.337816e-06, 1.291049e-06, 1.443986e-06, 
    1.418709e-06, 1.433738e-06, 1.489245e-06, 1.315445e-06, 1.403336e-06, 
    1.243224e-06, 1.289213e-06, 1.157327e-06, 1.222022e-06, 1.096624e-06, 
    1.045108e-06, 9.97818e-07, 9.439672e-07, 1.44748e-06, 1.46676e-06, 
    1.43233e-06, 1.38533e-06, 1.34242e-06, 1.286383e-06, 1.28072e-06, 
    1.270373e-06, 1.243774e-06, 1.221622e-06, 1.267104e-06, 1.216101e-06, 
    1.412863e-06, 1.30795e-06, 1.474075e-06, 1.423033e-06, 1.388083e-06, 
    1.40337e-06, 1.324891e-06, 1.306713e-06, 1.234114e-06, 1.271391e-06, 
    1.057699e-06, 1.149793e-06, 9.04036e-07, 9.696207e-07, 1.473524e-06, 
    1.447549e-06, 1.358871e-06, 1.400728e-06, 1.282688e-06, 1.254411e-06, 
    1.231661e-06, 1.20287e-06, 1.199787e-06, 1.182912e-06, 1.210627e-06, 
    1.184003e-06, 1.286265e-06, 1.240046e-06, 1.368878e-06, 1.336943e-06, 
    1.351591e-06, 1.367743e-06, 1.318193e-06, 1.26638e-06, 1.265294e-06, 
    1.248903e-06, 1.203265e-06, 1.28222e-06, 1.046081e-06, 1.189038e-06, 
    1.419477e-06, 1.370523e-06, 1.363612e-06, 1.382429e-06, 1.257232e-06, 
    1.30192e-06, 1.183324e-06, 1.214822e-06, 1.163432e-06, 1.188828e-06, 
    1.192588e-06, 1.225664e-06, 1.246481e-06, 1.299852e-06, 1.344093e-06, 
    1.379693e-06, 1.371376e-06, 1.33241e-06, 1.263246e-06, 1.199503e-06, 
    1.213324e-06, 1.167299e-06, 1.291075e-06, 1.238411e-06, 1.258634e-06, 
    1.206249e-06, 1.322483e-06, 1.223135e-06, 1.348485e-06, 1.337257e-06, 
    1.302815e-06, 1.234872e-06, 1.2201e-06, 1.204406e-06, 1.21408e-06, 
    1.261516e-06, 1.269378e-06, 1.30365e-06, 1.313186e-06, 1.339699e-06, 
    1.361839e-06, 1.341601e-06, 1.320503e-06, 1.2615e-06, 1.209466e-06, 
    1.153987e-06, 1.140615e-06, 1.077816e-06, 1.128786e-06, 1.045309e-06, 
    1.11605e-06, 9.951134e-07, 1.217512e-06, 1.118187e-06, 1.301262e-06, 
    1.280878e-06, 1.2444e-06, 1.162742e-06, 1.206493e-06, 1.155412e-06, 
    1.269687e-06, 1.33107e-06, 1.347196e-06, 1.377514e-06, 1.346507e-06, 
    1.349016e-06, 1.319641e-06, 1.329047e-06, 1.259564e-06, 1.296659e-06, 
    1.192679e-06, 1.155813e-06, 1.054884e-06, 9.953453e-07, 9.366034e-07, 
    9.112628e-07, 9.036237e-07, 9.004399e-07,
  4.082445e-07, 3.877676e-07, 3.917013e-07, 3.75533e-07, 3.84454e-07, 
    3.739371e-07, 4.040451e-07, 3.869661e-07, 3.978203e-07, 4.06378e-07, 
    3.452849e-07, 3.748214e-07, 3.161218e-07, 3.338516e-07, 2.904082e-07, 
    3.188412e-07, 2.848683e-07, 2.912089e-07, 2.723862e-07, 2.77701e-07, 
    2.544486e-07, 2.699543e-07, 2.428851e-07, 2.581021e-07, 2.556832e-07, 
    2.70475e-07, 3.687657e-07, 3.488835e-07, 3.699633e-07, 3.670832e-07, 
    3.683746e-07, 3.842674e-07, 3.924231e-07, 4.09837e-07, 4.066436e-07, 
    3.938705e-07, 3.657925e-07, 3.751899e-07, 3.517794e-07, 3.522984e-07, 
    3.272516e-07, 3.384091e-07, 2.979446e-07, 3.091332e-07, 2.774779e-07, 
    2.852446e-07, 2.778394e-07, 2.800727e-07, 2.778104e-07, 2.892539e-07, 
    2.843165e-07, 2.945131e-07, 3.36302e-07, 3.236755e-07, 3.62183e-07, 
    3.865676e-07, 4.032865e-07, 4.153973e-07, 4.136726e-07, 4.103955e-07, 
    3.937964e-07, 3.785546e-07, 3.671736e-07, 3.596735e-07, 3.52373e-07, 
    3.308035e-07, 3.197196e-07, 2.957108e-07, 2.99963e-07, 2.927828e-07, 
    2.860245e-07, 2.748886e-07, 2.767034e-07, 2.718623e-07, 2.929727e-07, 
    2.788354e-07, 3.024008e-07, 2.958404e-07, 3.50393e-07, 3.726414e-07, 
    3.823325e-07, 3.909429e-07, 4.123491e-07, 3.974952e-07, 4.033128e-07, 
    3.895551e-07, 3.809556e-07, 3.851952e-07, 3.594697e-07, 3.69347e-07, 
    3.190697e-07, 3.401927e-07, 2.868078e-07, 2.990874e-07, 2.83911e-07, 
    2.915961e-07, 2.785031e-07, 2.902703e-07, 2.700745e-07, 2.657927e-07, 
    2.687141e-07, 2.576011e-07, 2.90931e-07, 2.778386e-07, 3.853139e-07, 
    3.846204e-07, 3.814004e-07, 3.956726e-07, 3.965563e-07, 4.099242e-07, 
    3.980178e-07, 3.930084e-07, 3.804614e-07, 3.731495e-07, 3.662763e-07, 
    3.514276e-07, 3.352693e-07, 3.134303e-07, 2.982819e-07, 2.883789e-07, 
    2.94428e-07, 2.890835e-07, 2.950616e-07, 2.978894e-07, 2.673916e-07, 
    2.842702e-07, 2.591818e-07, 2.605336e-07, 2.717475e-07, 2.603811e-07, 
    3.84134e-07, 3.881316e-07, 4.021945e-07, 3.911643e-07, 4.113957e-07, 
    3.999968e-07, 3.935257e-07, 3.691367e-07, 3.639027e-07, 3.590852e-07, 
    3.49684e-07, 3.378326e-07, 3.176248e-07, 3.00646e-07, 2.856346e-07, 
    2.867189e-07, 2.863368e-07, 2.830408e-07, 2.912462e-07, 2.817073e-07, 
    2.801243e-07, 2.842733e-07, 2.607149e-07, 2.673192e-07, 2.605624e-07, 
    2.648497e-07, 3.868298e-07, 3.801309e-07, 3.837421e-07, 3.769674e-07, 
    3.81732e-07, 3.608104e-07, 3.546722e-07, 3.267751e-07, 3.38063e-07, 
    3.20208e-07, 3.362238e-07, 3.333514e-07, 3.196311e-07, 3.353471e-07, 
    3.015658e-07, 3.242308e-07, 2.829132e-07, 3.047028e-07, 2.815799e-07, 
    2.856985e-07, 2.789e-07, 2.728942e-07, 2.654529e-07, 2.520478e-07, 
    2.551145e-07, 2.441487e-07, 3.70272e-07, 3.618156e-07, 3.625576e-07, 
    3.538215e-07, 3.474408e-07, 3.338484e-07, 3.127153e-07, 3.205662e-07, 
    3.062443e-07, 3.034156e-07, 3.252104e-07, 3.117198e-07, 3.562217e-07, 
    3.487908e-07, 3.532055e-07, 3.695995e-07, 3.187442e-07, 3.442861e-07, 
    2.98035e-07, 3.111925e-07, 2.737455e-07, 2.920048e-07, 2.56812e-07, 
    2.42597e-07, 2.296778e-07, 2.151225e-07, 3.57251e-07, 3.629417e-07, 
    3.527915e-07, 3.390237e-07, 3.26544e-07, 3.103798e-07, 3.087546e-07, 
    3.057897e-07, 2.981916e-07, 2.918912e-07, 3.04854e-07, 2.903247e-07, 
    3.470767e-07, 3.165831e-07, 3.651051e-07, 3.500602e-07, 3.398271e-07, 
    3.442959e-07, 3.214714e-07, 3.162264e-07, 2.954414e-07, 3.060812e-07, 
    2.460579e-07, 2.716334e-07, 2.044398e-07, 2.220354e-07, 3.64942e-07, 
    3.572714e-07, 3.313181e-07, 3.435227e-07, 3.093192e-07, 3.012261e-07, 
    2.947434e-07, 2.865771e-07, 2.85705e-07, 2.809408e-07, 2.88773e-07, 
    2.812484e-07, 3.10346e-07, 2.971298e-07, 3.342284e-07, 3.249574e-07, 
    3.292038e-07, 3.33898e-07, 3.19537e-07, 3.046469e-07, 3.043363e-07, 
    2.996541e-07, 2.866892e-07, 3.09185e-07, 2.428646e-07, 2.826692e-07, 
    3.490161e-07, 3.347075e-07, 3.326964e-07, 3.381768e-07, 3.020316e-07, 
    3.148464e-07, 2.810568e-07, 2.89962e-07, 2.754594e-07, 2.826094e-07, 
    2.836707e-07, 2.930389e-07, 2.989636e-07, 3.142513e-07, 3.270289e-07, 
    3.373791e-07, 3.349556e-07, 3.236455e-07, 3.037505e-07, 2.856248e-07, 
    2.895375e-07, 2.765458e-07, 3.117274e-07, 2.966643e-07, 3.024322e-07, 
    2.875332e-07, 3.207757e-07, 2.923213e-07, 3.283027e-07, 3.250484e-07, 
    3.15104e-07, 2.956569e-07, 2.91459e-07, 2.870116e-07, 2.897516e-07, 
    3.032558e-07, 3.055049e-07, 3.153443e-07, 3.180924e-07, 3.257555e-07, 
    3.321808e-07, 3.263065e-07, 3.20204e-07, 3.032513e-07, 2.884441e-07, 
    2.728089e-07, 2.690639e-07, 2.516056e-07, 2.657596e-07, 2.426526e-07, 
    2.622102e-07, 2.289431e-07, 2.907252e-07, 2.628049e-07, 3.146569e-07, 
    3.088e-07, 2.983703e-07, 2.752656e-07, 2.876022e-07, 2.732084e-07, 
    3.055935e-07, 3.232578e-07, 3.279287e-07, 3.367438e-07, 3.277289e-07, 
    3.284568e-07, 3.199549e-07, 3.226727e-07, 3.026979e-07, 3.133326e-07, 
    2.836966e-07, 2.73321e-07, 2.452831e-07, 2.290059e-07, 2.131452e-07, 
    2.06366e-07, 2.043299e-07, 2.034824e-07,
  3.720525e-08, 3.489912e-08, 3.533964e-08, 3.353666e-08, 3.452895e-08, 
    3.33598e-08, 3.672969e-08, 3.48095e-08, 3.602726e-08, 3.699371e-08, 
    3.021941e-08, 3.345777e-08, 2.709295e-08, 2.898504e-08, 2.4398e-08, 
    2.738142e-08, 2.382525e-08, 2.4481e-08, 2.254531e-08, 2.308849e-08, 
    2.073229e-08, 2.229767e-08, 1.958046e-08, 2.109899e-08, 2.085605e-08, 
    2.235065e-08, 3.278808e-08, 3.061017e-08, 3.292029e-08, 3.260255e-08, 
    3.274494e-08, 3.450813e-08, 3.542062e-08, 3.738591e-08, 3.702378e-08, 
    3.558308e-08, 3.246037e-08, 3.34986e-08, 3.092533e-08, 3.098189e-08, 
    2.827753e-08, 2.947574e-08, 2.518167e-08, 2.635463e-08, 2.306564e-08, 
    2.386405e-08, 2.310267e-08, 2.333175e-08, 2.30997e-08, 2.427841e-08, 
    2.376835e-08, 2.482419e-08, 2.924866e-08, 2.789576e-08, 3.206345e-08, 
    3.4765e-08, 3.664393e-08, 3.801824e-08, 3.782186e-08, 3.744933e-08, 
    3.557476e-08, 3.387204e-08, 3.261249e-08, 3.178811e-08, 3.099003e-08, 
    2.865787e-08, 2.747471e-08, 2.494886e-08, 2.539243e-08, 2.464436e-08, 
    2.394453e-08, 2.280073e-08, 2.298634e-08, 2.249192e-08, 2.466407e-08, 
    2.320478e-08, 2.564749e-08, 2.496234e-08, 3.077441e-08, 3.321634e-08, 
    3.429243e-08, 3.525462e-08, 3.767131e-08, 3.599066e-08, 3.664691e-08, 
    3.509912e-08, 3.413907e-08, 3.461166e-08, 3.176578e-08, 3.285224e-08, 
    2.740567e-08, 2.966827e-08, 2.402543e-08, 2.530096e-08, 2.372655e-08, 
    2.452115e-08, 2.317071e-08, 2.438369e-08, 2.23099e-08, 2.187523e-08, 
    2.21716e-08, 2.10486e-08, 2.445218e-08, 2.310259e-08, 3.462492e-08, 
    3.454751e-08, 3.418857e-08, 3.57856e-08, 3.588498e-08, 3.739581e-08, 
    3.60495e-08, 3.548628e-08, 3.408406e-08, 3.327258e-08, 3.251364e-08, 
    3.0887e-08, 2.91375e-08, 2.68081e-08, 2.521687e-08, 2.418785e-08, 
    2.481534e-08, 2.426076e-08, 2.488126e-08, 2.51759e-08, 2.203734e-08, 
    2.376358e-08, 2.12076e-08, 2.134376e-08, 2.248022e-08, 2.132839e-08, 
    3.449324e-08, 3.493981e-08, 3.652055e-08, 3.527942e-08, 3.756293e-08, 
    3.627254e-08, 3.554437e-08, 3.282904e-08, 3.225241e-08, 3.172365e-08, 
    3.069717e-08, 2.941357e-08, 2.725229e-08, 2.546385e-08, 2.390429e-08, 
    2.401624e-08, 2.397678e-08, 2.363693e-08, 2.448486e-08, 2.349972e-08, 
    2.333706e-08, 2.376389e-08, 2.136204e-08, 2.202998e-08, 2.134666e-08, 
    2.177972e-08, 3.479425e-08, 3.40473e-08, 3.444952e-08, 3.369577e-08, 
    3.422551e-08, 3.19128e-08, 3.124093e-08, 2.822662e-08, 2.943842e-08, 
    2.752661e-08, 2.924023e-08, 2.893129e-08, 2.746533e-08, 2.914585e-08, 
    2.556009e-08, 2.795499e-08, 2.362379e-08, 2.588886e-08, 2.348662e-08, 
    2.391088e-08, 2.32114e-08, 2.259712e-08, 2.184079e-08, 2.049201e-08, 
    2.0799e-08, 1.970565e-08, 3.295438e-08, 3.202312e-08, 3.210458e-08, 
    3.114803e-08, 3.045333e-08, 2.898468e-08, 2.673252e-08, 2.756468e-08, 
    2.605069e-08, 2.575382e-08, 2.805947e-08, 2.66274e-08, 3.141024e-08, 
    3.060006e-08, 3.108082e-08, 3.288013e-08, 2.737109e-08, 3.011111e-08, 
    2.519111e-08, 2.657174e-08, 2.268398e-08, 2.456359e-08, 2.096934e-08, 
    1.955195e-08, 1.828176e-08, 1.68721e-08, 3.152281e-08, 3.214678e-08, 
    3.103566e-08, 2.954206e-08, 2.820191e-08, 2.648602e-08, 2.631476e-08, 
    2.600294e-08, 2.520744e-08, 2.455178e-08, 2.590471e-08, 2.438932e-08, 
    3.041384e-08, 2.714183e-08, 3.238469e-08, 3.073814e-08, 2.962879e-08, 
    3.011216e-08, 2.766097e-08, 2.710402e-08, 2.49208e-08, 2.603356e-08, 
    1.989516e-08, 2.246862e-08, 1.585238e-08, 1.753874e-08, 3.236673e-08, 
    3.152504e-08, 2.871303e-08, 3.00284e-08, 2.637422e-08, 2.552453e-08, 
    2.484815e-08, 2.40016e-08, 2.391155e-08, 2.342093e-08, 2.422862e-08, 
    2.345253e-08, 2.648244e-08, 2.50967e-08, 2.902553e-08, 2.803248e-08, 
    2.848641e-08, 2.899002e-08, 2.745528e-08, 2.588297e-08, 2.585037e-08, 
    2.536016e-08, 2.401324e-08, 2.636009e-08, 1.957847e-08, 2.359873e-08, 
    3.062452e-08, 2.907708e-08, 2.886093e-08, 2.945069e-08, 2.560883e-08, 
    2.695788e-08, 2.343284e-08, 2.435175e-08, 2.285907e-08, 2.359252e-08, 
    2.370179e-08, 2.467094e-08, 2.528803e-08, 2.689491e-08, 2.825373e-08, 
    2.936468e-08, 2.910373e-08, 2.789255e-08, 2.578895e-08, 2.390329e-08, 
    2.430778e-08, 2.29702e-08, 2.662819e-08, 2.504818e-08, 2.565079e-08, 
    2.410039e-08, 2.758697e-08, 2.459648e-08, 2.838995e-08, 2.804218e-08, 
    2.698515e-08, 2.494326e-08, 2.450694e-08, 2.404649e-08, 2.432995e-08, 
    2.573709e-08, 2.597303e-08, 2.701058e-08, 2.73019e-08, 2.811767e-08, 
    2.880557e-08, 2.817653e-08, 2.752618e-08, 2.57366e-08, 2.419461e-08, 
    2.258842e-08, 2.220715e-08, 2.044785e-08, 2.187189e-08, 1.955749e-08, 
    2.151296e-08, 1.821009e-08, 2.443087e-08, 2.157299e-08, 2.693782e-08, 
    2.631953e-08, 2.522611e-08, 2.283928e-08, 2.410752e-08, 2.262918e-08, 
    2.598233e-08, 2.785124e-08, 2.834994e-08, 2.929623e-08, 2.832856e-08, 
    2.840644e-08, 2.749969e-08, 2.778887e-08, 2.567861e-08, 2.679775e-08, 
    2.370447e-08, 2.264067e-08, 1.98182e-08, 1.82162e-08, 1.668237e-08, 
    1.603528e-08, 1.584196e-08, 1.576162e-08,
  1.074225e-09, 9.912241e-10, 1.00697e-09, 9.428566e-10, 9.780327e-10, 
    9.366153e-10, 1.056995e-09, 9.880277e-10, 1.031652e-09, 1.066553e-09, 
    8.272728e-10, 9.400712e-10, 7.213313e-10, 7.850844e-10, 6.325266e-10, 
    7.309783e-10, 6.139706e-10, 6.352246e-10, 5.729226e-10, 5.902703e-10, 
    5.158114e-10, 5.650492e-10, 4.801855e-10, 5.27262e-10, 5.196701e-10, 
    5.667316e-10, 9.16499e-10, 8.407229e-10, 9.211428e-10, 9.09991e-10, 
    9.149845e-10, 9.772924e-10, 1.009871e-09, 1.080785e-09, 1.067643e-09, 
    1.015694e-09, 9.050101e-10, 9.41512e-10, 8.516012e-10, 8.535571e-10, 
    7.611139e-10, 8.017997e-10, 6.580989e-10, 6.967619e-10, 5.895384e-10, 
    6.152234e-10, 5.907249e-10, 5.98074e-10, 5.906295e-10, 6.286423e-10, 
    6.12133e-10, 6.464075e-10, 7.940552e-10, 7.482439e-10, 8.911351e-10, 
    9.864416e-10, 1.053894e-09, 1.103815e-09, 1.096651e-09, 1.08309e-09, 
    1.015396e-09, 9.54715e-10, 9.10339e-10, 8.815365e-10, 8.538385e-10, 
    7.739818e-10, 7.341037e-10, 6.504802e-10, 6.650122e-10, 6.40543e-10, 
    6.178251e-10, 5.810669e-10, 5.869997e-10, 5.712233e-10, 6.411847e-10, 
    5.939986e-10, 6.733981e-10, 6.509206e-10, 8.463895e-10, 9.315586e-10, 
    9.696249e-10, 1.003927e-09, 1.091167e-09, 1.030336e-09, 1.054002e-09, 
    9.983665e-10, 9.641793e-10, 9.80977e-10, 8.807587e-10, 9.187517e-10, 
    7.317901e-10, 8.083783e-10, 6.204426e-10, 6.620101e-10, 6.107839e-10, 
    6.365307e-10, 5.929057e-10, 6.320608e-10, 5.654376e-10, 5.516708e-10, 
    5.610499e-10, 5.256853e-10, 6.34287e-10, 5.907224e-10, 9.81449e-10, 
    9.786932e-10, 9.659359e-10, 1.022964e-09, 1.026535e-09, 1.081145e-09, 
    1.032453e-09, 1.012224e-09, 9.62228e-10, 9.335399e-10, 9.068751e-10, 
    8.502767e-10, 7.902703e-10, 7.118311e-10, 6.592525e-10, 6.257041e-10, 
    6.461184e-10, 6.280693e-10, 6.482709e-10, 6.579097e-10, 5.56797e-10, 
    6.11979e-10, 5.306634e-10, 5.34934e-10, 5.708512e-10, 5.344516e-10, 
    9.767623e-10, 9.926759e-10, 1.049436e-09, 1.004814e-09, 1.087222e-09, 
    1.040487e-09, 1.014306e-09, 9.179373e-10, 8.977346e-10, 8.792926e-10, 
    8.437215e-10, 7.996778e-10, 7.266561e-10, 6.673583e-10, 6.165237e-10, 
    6.20145e-10, 6.188681e-10, 6.078938e-10, 6.353502e-10, 6.034748e-10, 
    5.982448e-10, 6.11989e-10, 5.355079e-10, 5.565637e-10, 5.350251e-10, 
    5.48655e-10, 9.874828e-10, 9.609245e-10, 9.75207e-10, 9.484785e-10, 
    9.672475e-10, 8.858813e-10, 8.625273e-10, 7.593953e-10, 8.005258e-10, 
    7.358434e-10, 7.937678e-10, 7.832579e-10, 7.337897e-10, 7.90554e-10, 
    6.705226e-10, 7.502382e-10, 6.074704e-10, 6.813555e-10, 6.030532e-10, 
    6.16737e-10, 5.942106e-10, 5.745727e-10, 5.505829e-10, 5.083363e-10, 
    5.178904e-10, 4.840318e-10, 9.223406e-10, 8.89728e-10, 8.925703e-10, 
    8.593076e-10, 8.353169e-10, 7.85072e-10, 7.093147e-10, 7.371199e-10, 
    6.866995e-10, 6.769009e-10, 7.537568e-10, 7.058185e-10, 8.683995e-10, 
    8.403727e-10, 8.569806e-10, 9.197316e-10, 7.306321e-10, 8.235517e-10, 
    6.584082e-10, 7.039681e-10, 5.773411e-10, 6.379124e-10, 5.232073e-10, 
    4.793109e-10, 4.406613e-10, 3.985726e-10, 8.723087e-10, 8.940439e-10, 
    8.554171e-10, 8.04065e-10, 7.585608e-10, 7.011212e-10, 6.954401e-10, 
    6.851215e-10, 6.589433e-10, 6.375275e-10, 6.818781e-10, 6.322439e-10, 
    8.339591e-10, 7.229635e-10, 9.02361e-10, 8.451359e-10, 8.070282e-10, 
    8.235873e-10, 7.403513e-10, 7.217e-10, 6.495631e-10, 6.861333e-10, 
    4.898671e-10, 5.704823e-10, 3.68679e-10, 4.183686e-10, 9.017323e-10, 
    8.723859e-10, 7.758504e-10, 8.207127e-10, 6.974115e-10, 6.693527e-10, 
    6.471895e-10, 6.196714e-10, 6.167588e-10, 6.009402e-10, 6.270265e-10, 
    6.019565e-10, 7.010026e-10, 6.553159e-10, 7.864606e-10, 7.528474e-10, 
    7.681742e-10, 7.852531e-10, 7.334517e-10, 6.811607e-10, 6.800843e-10, 
    6.639528e-10, 6.200499e-10, 6.969427e-10, 4.801257e-10, 6.066646e-10, 
    8.412153e-10, 7.882144e-10, 7.808683e-10, 8.009441e-10, 6.721259e-10, 
    7.168227e-10, 6.013232e-10, 6.310231e-10, 5.829301e-10, 6.064629e-10, 
    6.099852e-10, 6.414087e-10, 6.615856e-10, 7.147233e-10, 7.603101e-10, 
    7.980097e-10, 7.891204e-10, 7.481358e-10, 6.780592e-10, 6.164917e-10, 
    6.295959e-10, 5.864833e-10, 7.058442e-10, 6.537283e-10, 6.735073e-10, 
    6.228696e-10, 7.378678e-10, 6.389847e-10, 7.649119e-10, 7.531742e-10, 
    7.177323e-10, 6.502973e-10, 6.360683e-10, 6.211242e-10, 6.303152e-10, 
    6.763496e-10, 6.841336e-10, 7.185806e-10, 7.283155e-10, 7.557188e-10, 
    7.789889e-10, 7.577043e-10, 7.35829e-10, 6.763333e-10, 6.259236e-10, 
    5.742956e-10, 5.621767e-10, 5.069658e-10, 5.515658e-10, 4.794819e-10, 
    5.402528e-10, 4.385019e-10, 6.335952e-10, 5.421406e-10, 7.161535e-10, 
    6.955982e-10, 6.595557e-10, 5.822987e-10, 6.231008e-10, 5.755947e-10, 
    6.844407e-10, 7.467465e-10, 7.635598e-10, 7.956761e-10, 7.628372e-10, 
    7.654694e-10, 7.349401e-10, 7.446483e-10, 6.744232e-10, 7.114861e-10, 
    6.100718e-10, 5.759607e-10, 4.874955e-10, 4.386852e-10, 3.929742e-10, 
    3.740055e-10, 3.683757e-10, 3.660416e-10,
  8.656255e-12, 7.785162e-12, 7.948839e-12, 7.287171e-12, 7.64862e-12, 
    7.223447e-12, 8.473755e-12, 7.752031e-12, 8.206907e-12, 8.574884e-12, 
    6.127883e-12, 7.258717e-12, 5.106666e-12, 5.71621e-12, 4.284566e-12, 
    5.197904e-12, 4.117021e-12, 4.309048e-12, 3.751928e-12, 3.905274e-12, 
    3.257365e-12, 3.682799e-12, 2.957273e-12, 3.35522e-12, 3.290265e-12, 
    3.697546e-12, 7.018902e-12, 6.260457e-12, 7.066004e-12, 6.953013e-12, 
    7.003557e-12, 7.640975e-12, 7.979086e-12, 8.725957e-12, 8.586435e-12, 
    8.039852e-12, 6.902677e-12, 7.273428e-12, 6.368123e-12, 6.387528e-12, 
    5.485216e-12, 5.87854e-12, 4.517917e-12, 4.875965e-12, 3.898776e-12, 
    4.128281e-12, 3.909312e-12, 3.974711e-12, 3.908466e-12, 4.249364e-12, 
    4.100509e-12, 4.410879e-12, 5.803203e-12, 5.362086e-12, 6.762886e-12, 
    7.735608e-12, 8.441005e-12, 8.971635e-12, 8.895058e-12, 8.750487e-12, 
    8.036734e-12, 7.408584e-12, 6.956529e-12, 6.666552e-12, 6.390321e-12, 
    5.608963e-12, 5.227537e-12, 4.448103e-12, 4.581481e-12, 4.357412e-12, 
    4.151693e-12, 3.823746e-12, 3.876257e-12, 3.736986e-12, 4.363253e-12, 
    3.938416e-12, 4.658856e-12, 4.452128e-12, 6.316501e-12, 7.171903e-12, 
    7.561885e-12, 7.917153e-12, 8.836525e-12, 8.193097e-12, 8.442145e-12, 
    7.859309e-12, 7.505806e-12, 7.679047e-12, 6.658761e-12, 7.041742e-12, 
    5.205596e-12, 5.942711e-12, 4.17528e-12, 4.553853e-12, 4.088398e-12, 
    4.320912e-12, 3.928695e-12, 4.280336e-12, 3.686204e-12, 3.566021e-12, 
    3.6478e-12, 3.341703e-12, 4.300534e-12, 3.909292e-12, 7.683929e-12, 
    7.655443e-12, 7.52388e-12, 8.11586e-12, 8.153258e-12, 8.729788e-12, 
    8.215306e-12, 8.003617e-12, 7.485736e-12, 7.192088e-12, 6.921512e-12, 
    6.354992e-12, 5.766467e-12, 5.017176e-12, 4.52851e-12, 4.222782e-12, 
    4.408239e-12, 4.244176e-12, 4.427899e-12, 4.516178e-12, 3.610666e-12, 
    4.099128e-12, 3.384415e-12, 3.421155e-12, 3.733715e-12, 3.417e-12, 
    7.635498e-12, 7.800217e-12, 8.393968e-12, 7.926383e-12, 8.794475e-12, 
    8.299721e-12, 8.025358e-12, 7.033488e-12, 6.829293e-12, 6.644079e-12, 
    6.29008e-12, 5.857878e-12, 5.156977e-12, 4.603101e-12, 4.139978e-12, 
    4.172596e-12, 4.161087e-12, 4.062483e-12, 4.310187e-12, 4.02293e-12, 
    3.976236e-12, 4.099216e-12, 3.426099e-12, 3.608629e-12, 3.42194e-12, 
    3.539814e-12, 7.746378e-12, 7.472338e-12, 7.619441e-12, 7.344674e-12, 
    7.537387e-12, 6.710126e-12, 6.476702e-12, 5.468742e-12, 5.866134e-12, 
    5.244047e-12, 5.800411e-12, 5.698534e-12, 5.224563e-12, 5.769213e-12, 
    4.632298e-12, 5.381131e-12, 4.058689e-12, 4.732559e-12, 4.019161e-12, 
    4.141897e-12, 3.940299e-12, 3.766455e-12, 3.556561e-12, 3.193841e-12, 
    3.275078e-12, 2.989344e-12, 7.078164e-12, 6.748746e-12, 6.777313e-12, 
    6.444657e-12, 6.207077e-12, 5.716087e-12, 4.99353e-12, 5.256166e-12, 
    4.782185e-12, 4.691264e-12, 5.414749e-12, 4.960725e-12, 6.535217e-12, 
    6.256985e-12, 6.421528e-12, 7.051685e-12, 5.194619e-12, 6.091306e-12, 
    4.520756e-12, 4.943379e-12, 3.790853e-12, 4.333477e-12, 3.32049e-12, 
    2.949994e-12, 2.63247e-12, 2.296663e-12, 6.574236e-12, 6.792136e-12, 
    6.405995e-12, 5.900624e-12, 5.460739e-12, 4.916722e-12, 4.863622e-12, 
    4.767518e-12, 4.525668e-12, 4.329973e-12, 4.737401e-12, 4.281996e-12, 
    6.193706e-12, 5.122074e-12, 6.875937e-12, 6.304082e-12, 5.929529e-12, 
    6.091649e-12, 5.286884e-12, 5.11014e-12, 4.439715e-12, 4.77692e-12, 
    3.03816e-12, 3.730476e-12, 2.064915e-12, 2.453265e-12, 6.869591e-12, 
    6.575006e-12, 5.626974e-12, 6.063435e-12, 4.882033e-12, 4.621495e-12, 
    4.418018e-12, 4.168329e-12, 4.142093e-12, 4.000286e-12, 4.23474e-12, 
    4.009361e-12, 4.915612e-12, 4.492383e-12, 5.729532e-12, 5.406055e-12, 
    5.553027e-12, 5.71784e-12, 5.221344e-12, 4.730747e-12, 4.720759e-12, 
    4.571731e-12, 4.171757e-12, 4.877653e-12, 2.956786e-12, 4.051486e-12, 
    6.265303e-12, 5.746535e-12, 5.675425e-12, 5.870205e-12, 4.6471e-12, 
    5.064147e-12, 4.003704e-12, 4.270928e-12, 3.840219e-12, 4.049666e-12, 
    4.081233e-12, 4.365292e-12, 4.549951e-12, 5.04438e-12, 5.477508e-12, 
    5.841642e-12, 5.755309e-12, 5.361054e-12, 4.701994e-12, 4.139692e-12, 
    4.258e-12, 3.871679e-12, 4.960962e-12, 4.477836e-12, 4.65987e-12, 
    4.197177e-12, 5.263273e-12, 4.343241e-12, 5.521669e-12, 5.409179e-12, 
    5.072718e-12, 4.446432e-12, 4.31671e-12, 4.181429e-12, 4.264513e-12, 
    4.686162e-12, 4.75834e-12, 5.080713e-12, 5.172677e-12, 5.43352e-12, 
    5.657264e-12, 5.452533e-12, 5.243909e-12, 4.68601e-12, 4.224769e-12, 
    3.764015e-12, 3.657653e-12, 3.182233e-12, 3.565114e-12, 2.951426e-12, 
    3.467058e-12, 2.614991e-12, 4.294264e-12, 3.48337e-12, 5.057843e-12, 
    4.865098e-12, 4.531299e-12, 3.83464e-12, 4.199264e-12, 3.775462e-12, 
    4.761192e-12, 5.347803e-12, 5.508685e-12, 5.818952e-12, 5.501749e-12, 
    5.527025e-12, 5.235466e-12, 5.327794e-12, 4.668336e-12, 5.013929e-12, 
    4.08201e-12, 3.778685e-12, 3.018295e-12, 2.616469e-12, 2.252816e-12, 
    2.105776e-12, 2.062593e-12, 2.044751e-12,
  1.093206e-14, 9.020758e-15, 9.371128e-15, 7.981011e-15, 8.731677e-15, 
    7.850901e-15, 1.052231e-14, 8.950353e-15, 9.93193e-15, 1.074876e-14, 
    5.726269e-15, 7.922829e-15, 3.958056e-15, 4.986867e-15, 2.709109e-15, 
    4.106791e-15, 2.476152e-15, 2.743782e-15, 1.996288e-15, 2.193069e-15, 
    1.411913e-15, 1.90991e-15, 1.097729e-15, 1.521173e-15, 1.448282e-15, 
    1.928214e-15, 7.437918e-15, 5.971557e-15, 7.532382e-15, 7.306431e-15, 
    7.407226e-15, 8.71559e-15, 9.436355e-15, 1.10898e-14, 1.077472e-14, 
    9.567756e-15, 7.206488e-15, 7.952877e-15, 6.173195e-15, 6.209781e-15, 
    4.587397e-15, 5.274295e-15, 3.046199e-15, 3.590657e-15, 2.184588e-15, 
    2.491554e-15, 2.198347e-15, 2.28447e-15, 2.197241e-15, 2.659512e-15, 
    2.45361e-15, 2.889778e-15, 5.140226e-15, 4.379176e-15, 6.931265e-15, 
    8.915536e-15, 1.044929e-14, 1.165128e-14, 1.147537e-14, 1.114549e-14, 
    9.561003e-15, 8.230765e-15, 7.313413e-15, 6.743631e-15, 6.215053e-15, 
    4.800012e-15, 4.155499e-15, 2.943842e-15, 3.140495e-15, 2.812781e-15, 
    2.523712e-15, 2.087572e-15, 2.155295e-15, 1.977496e-15, 2.821149e-15, 
    2.236523e-15, 3.256672e-15, 2.949701e-15, 6.076274e-15, 7.746149e-15, 
    8.549635e-15, 9.302977e-15, 1.134146e-14, 9.901674e-15, 1.045183e-14, 
    9.178949e-15, 8.432522e-15, 8.795832e-15, 6.728529e-15, 7.483672e-15, 
    4.119408e-15, 5.389419e-15, 2.556264e-15, 3.099382e-15, 2.437127e-15, 
    2.760645e-15, 2.223744e-15, 2.703118e-15, 1.914131e-15, 1.767379e-15, 
    1.866745e-15, 1.505881e-15, 2.731699e-15, 2.198324e-15, 8.806144e-15, 
    8.746054e-15, 8.470197e-15, 9.732933e-15, 9.814521e-15, 1.109849e-14, 
    9.950349e-15, 9.489319e-15, 8.390742e-15, 7.787113e-15, 7.243823e-15, 
    6.148483e-15, 5.075279e-15, 3.814046e-15, 3.06184e-15, 2.622288e-15, 
    2.885955e-15, 2.652228e-15, 2.914447e-15, 3.043629e-15, 1.821365e-15, 
    2.45173e-15, 1.554394e-15, 1.59661e-15, 1.973393e-15, 1.591813e-15, 
    8.704054e-15, 9.052795e-15, 1.034469e-14, 9.322802e-15, 1.124554e-14, 
    1.013608e-14, 9.536366e-15, 7.46714e-15, 7.061564e-15, 6.700109e-15, 
    6.026777e-15, 5.237408e-15, 4.039823e-15, 3.17281e-15, 2.507599e-15, 
    2.552549e-15, 2.536656e-15, 2.402005e-15, 2.745398e-15, 2.348766e-15, 
    2.286497e-15, 2.451845e-15, 1.602325e-15, 1.818882e-15, 1.597516e-15, 
    1.735978e-15, 8.938332e-15, 8.362894e-15, 8.670287e-15, 8.09899e-15, 
    8.498397e-15, 6.828309e-15, 6.378847e-15, 4.559359e-15, 5.252141e-15, 
    4.182722e-15, 5.135275e-15, 4.955899e-15, 4.150616e-15, 5.080111e-15, 
    3.21664e-15, 4.411179e-15, 2.396879e-15, 3.368771e-15, 2.343716e-15, 
    2.510236e-15, 2.238996e-15, 2.014628e-15, 1.756016e-15, 1.342733e-15, 
    1.43144e-15, 1.129748e-15, 7.556824e-15, 6.903623e-15, 6.959496e-15, 
    6.317909e-15, 5.872336e-15, 4.986646e-15, 3.776305e-15, 4.202736e-15, 
    3.444967e-15, 3.305788e-15, 4.467815e-15, 3.724174e-15, 6.490564e-15, 
    5.965057e-15, 6.274065e-15, 7.503627e-15, 4.101393e-15, 5.659166e-15, 
    3.050389e-15, 3.696705e-15, 2.045572e-15, 2.778561e-15, 1.482019e-15, 
    1.09052e-15, 7.955706e-16, 5.284482e-16, 6.565416e-15, 6.988554e-15, 
    6.244664e-15, 5.313831e-15, 4.545739e-15, 3.654644e-15, 3.57136e-15, 
    3.422379e-15, 3.057639e-15, 2.773552e-15, 3.376168e-15, 2.705462e-15, 
    5.84762e-15, 3.983029e-15, 7.153567e-15, 6.052983e-15, 5.365705e-15, 
    5.659782e-15, 4.253641e-15, 3.963665e-15, 2.931627e-15, 3.436852e-15, 
    1.17923e-15, 1.969338e-15, 3.733147e-16, 6.470179e-16, 7.141021e-15, 
    6.566891e-15, 4.831204e-15, 5.608224e-15, 3.600158e-15, 3.200389e-15, 
    2.900114e-15, 2.546659e-15, 2.510507e-15, 2.31849e-15, 2.639008e-15, 
    2.330604e-15, 3.652897e-15, 3.008612e-15, 5.010242e-15, 4.453144e-15, 
    4.703476e-15, 4.989718e-15, 4.145283e-15, 3.365987e-15, 3.350712e-15, 
    3.125968e-15, 2.551431e-15, 3.593301e-15, 1.097266e-15, 2.38719e-15, 
    5.980532e-15, 5.040161e-15, 4.915508e-15, 5.259401e-15, 3.238929e-15, 
    3.889389e-15, 2.32305e-15, 2.689844e-15, 2.108726e-15, 2.384703e-15, 
    2.427398e-15, 2.824075e-15, 3.09359e-15, 3.857618e-15, 4.574265e-15, 
    5.208478e-15, 5.055591e-15, 4.377443e-15, 3.322116e-15, 2.507212e-15, 
    2.67165e-15, 2.149357e-15, 3.724543e-15, 2.987279e-15, 3.258216e-15, 
    2.586623e-15, 4.214499e-15, 2.792529e-15, 4.64967e-15, 4.45841e-15, 
    3.903194e-15, 2.941413e-15, 2.754667e-15, 2.564778e-15, 2.680805e-15, 
    3.298047e-15, 3.408272e-15, 3.916083e-15, 4.065458e-15, 4.49956e-15, 
    4.883842e-15, 4.531799e-15, 4.182489e-15, 3.297809e-15, 2.625069e-15, 
    2.011546e-15, 1.878856e-15, 1.330256e-15, 1.766298e-15, 1.091954e-15, 
    1.650016e-15, 7.805094e-16, 2.722836e-15, 1.66913e-15, 3.87924e-15, 
    3.573665e-15, 3.065975e-15, 2.101565e-15, 2.589524e-15, 2.026038e-15, 
    3.412652e-15, 4.355245e-15, 4.627454e-15, 5.16815e-15, 4.615602e-15, 
    4.658846e-15, 4.168549e-15, 4.32177e-15, 3.271017e-15, 3.808845e-15, 
    2.428456e-15, 2.030122e-15, 1.158985e-15, 7.817703e-16, 4.97194e-16, 
    3.988428e-16, 3.718863e-16, 3.610095e-16,
  3.698125e-20, 3.058219e-20, 3.175642e-20, 2.709416e-20, 2.961295e-20, 
    2.665729e-20, 3.561066e-20, 3.034617e-20, 3.363474e-20, 3.636822e-20, 
    1.950962e-20, 2.689881e-20, 1.353641e-20, 1.701502e-20, 9.299156e-21, 
    1.403992e-20, 8.506522e-21, 9.41706e-21, 6.870922e-21, 7.542145e-21, 
    4.872744e-21, 6.576046e-21, 3.794725e-21, 5.246964e-21, 4.997347e-21, 
    6.638544e-21, 2.527004e-20, 2.033628e-20, 2.558743e-20, 2.482816e-20, 
    2.51669e-20, 2.9559e-20, 3.197496e-20, 3.750869e-20, 3.645505e-20, 
    3.241515e-20, 2.449222e-20, 2.69997e-20, 2.101553e-20, 2.113874e-20, 
    1.566546e-20, 1.798524e-20, 1.044469e-20, 1.229178e-20, 7.513231e-21, 
    8.558954e-21, 7.560138e-21, 7.85367e-21, 7.556367e-21, 9.130473e-21, 
    8.42978e-21, 9.91332e-21, 1.753277e-20, 1.496147e-20, 2.356683e-20, 
    3.022944e-20, 3.536637e-20, 3.938539e-20, 3.879754e-20, 3.769489e-20, 
    3.239253e-20, 2.79325e-20, 2.485163e-20, 2.293567e-20, 2.115649e-20, 
    1.638392e-20, 1.420477e-20, 1.009701e-20, 1.076486e-20, 9.651635e-21, 
    8.668414e-21, 7.182384e-21, 7.413354e-21, 6.806783e-21, 9.68008e-21, 
    7.690271e-21, 1.115916e-20, 1.011692e-20, 2.068907e-20, 2.630551e-20, 
    2.900238e-20, 3.152806e-20, 3.834998e-20, 3.353343e-20, 3.537487e-20, 
    3.111242e-20, 2.86095e-20, 2.982808e-20, 2.288486e-20, 2.542378e-20, 
    1.408263e-20, 1.837367e-20, 8.779201e-21, 1.062528e-20, 8.373659e-21, 
    9.474397e-21, 7.646713e-21, 9.278781e-21, 6.590461e-21, 6.089134e-21, 
    6.428634e-21, 5.194609e-21, 9.375976e-21, 7.560059e-21, 2.986266e-20, 
    2.966116e-20, 2.87359e-20, 3.296839e-20, 3.324161e-20, 3.753775e-20, 
    3.369641e-20, 3.215239e-20, 2.846932e-20, 2.644308e-20, 2.461772e-20, 
    2.093229e-20, 1.731353e-20, 1.304868e-20, 1.04978e-20, 9.003849e-21, 
    9.900328e-21, 9.105698e-21, 9.997143e-21, 1.043596e-20, 6.273612e-21, 
    8.42338e-21, 5.360686e-21, 5.505159e-21, 6.792776e-21, 5.488744e-21, 
    2.952031e-20, 3.068959e-20, 3.501634e-20, 3.15945e-20, 3.802936e-20, 
    3.431819e-20, 3.231e-20, 2.536823e-20, 2.400499e-20, 2.278925e-20, 
    2.052232e-20, 1.786076e-20, 1.381324e-20, 1.087455e-20, 8.613572e-21, 
    8.766558e-21, 8.71247e-21, 8.254058e-21, 9.422557e-21, 8.072728e-21, 
    7.860578e-21, 8.423772e-21, 5.524713e-21, 6.26513e-21, 5.50826e-21, 
    5.981804e-21, 3.030587e-20, 2.837588e-20, 2.940706e-20, 2.749022e-20, 
    2.883049e-20, 2.322053e-20, 2.170801e-20, 1.557069e-20, 1.791048e-20, 
    1.429688e-20, 1.751606e-20, 1.691045e-20, 1.418824e-20, 1.732984e-20, 
    1.102331e-20, 1.50697e-20, 8.2366e-21, 1.153946e-20, 8.055526e-21, 
    8.622547e-21, 7.698698e-21, 6.93351e-21, 6.050297e-21, 4.635632e-21, 
    4.93965e-21, 3.904733e-21, 2.566955e-20, 2.347386e-20, 2.366177e-20, 
    2.150285e-20, 2.000194e-20, 1.701427e-20, 1.292083e-20, 1.436461e-20, 
    1.179787e-20, 1.132581e-20, 1.526121e-20, 1.27442e-20, 2.208408e-20, 
    2.031438e-20, 2.135522e-20, 2.549082e-20, 1.402165e-20, 1.928339e-20, 
    1.045892e-20, 1.265114e-20, 7.039101e-21, 9.535305e-21, 5.112895e-21, 
    3.769953e-21, 2.754694e-21, 1.8317e-21, 2.233601e-20, 2.375949e-20, 
    2.125621e-20, 1.811864e-20, 1.552465e-20, 1.250863e-20, 1.222638e-20, 
    1.172128e-20, 1.048354e-20, 9.518278e-21, 1.156455e-20, 9.286756e-21, 
    1.991864e-20, 1.362097e-20, 2.431432e-20, 2.061061e-20, 1.829366e-20, 
    1.928547e-20, 1.453684e-20, 1.35554e-20, 1.005552e-20, 1.177036e-20, 
    4.074667e-21, 6.778935e-21, 1.293535e-21, 2.241873e-21, 2.427214e-20, 
    2.234097e-20, 1.648929e-20, 1.911163e-20, 1.232398e-20, 1.096815e-20, 
    9.948445e-21, 8.746512e-21, 8.623469e-21, 7.969585e-21, 9.060726e-21, 
    8.010858e-21, 1.25027e-20, 1.031703e-20, 1.709395e-20, 1.52116e-20, 
    1.605776e-20, 1.702465e-20, 1.417019e-20, 1.153002e-20, 1.147821e-20, 
    1.071554e-20, 8.762752e-21, 1.230074e-20, 3.793133e-21, 8.203604e-21, 
    2.036652e-20, 1.719496e-20, 1.677404e-20, 1.793498e-20, 1.109895e-20, 
    1.330388e-20, 7.985122e-21, 9.233638e-21, 7.25454e-21, 8.195134e-21, 
    8.340531e-21, 9.690025e-21, 1.060561e-20, 1.319627e-20, 1.562108e-20, 
    1.776313e-20, 1.724706e-20, 1.495561e-20, 1.13812e-20, 8.612254e-21, 
    9.171759e-21, 7.393106e-21, 1.274546e-20, 1.024458e-20, 1.11644e-20, 
    8.882505e-21, 1.440441e-20, 9.582793e-21, 1.587593e-20, 1.522941e-20, 
    1.335063e-20, 1.008876e-20, 9.454072e-21, 8.808173e-21, 9.202898e-21, 
    1.129954e-20, 1.167343e-20, 1.339428e-20, 1.390002e-20, 1.536854e-20, 
    1.666709e-20, 1.547753e-20, 1.42961e-20, 1.129874e-20, 9.01331e-21, 
    6.922992e-21, 6.469998e-21, 4.592853e-21, 6.085442e-21, 3.774879e-21, 
    5.687863e-21, 2.702751e-21, 9.345836e-21, 5.753239e-21, 1.326951e-20, 
    1.223419e-20, 1.051184e-20, 7.230114e-21, 8.892374e-21, 6.972446e-21, 
    1.168829e-20, 1.488053e-20, 1.580085e-20, 1.762702e-20, 1.57608e-20, 
    1.590695e-20, 1.424893e-20, 1.476731e-20, 1.120783e-20, 1.303106e-20, 
    8.344132e-21, 6.986383e-21, 4.005151e-21, 2.7071e-21, 1.723428e-21, 
    1.38223e-21, 1.288571e-21, 1.25076e-21,
  2.715277e-26, 2.247312e-26, 2.333209e-26, 1.992079e-26, 2.176401e-26, 
    1.960103e-26, 2.615073e-26, 2.230046e-26, 2.470587e-26, 2.67046e-26, 
    1.436607e-26, 1.977781e-26, 9.985117e-27, 1.253728e-26, 6.871883e-27, 
    1.035469e-26, 6.288845e-27, 6.95859e-27, 5.08489e-27, 5.579126e-27, 
    3.612038e-27, 4.867693e-27, 2.816175e-27, 3.888079e-27, 3.703962e-27, 
    4.913731e-27, 1.85855e-26, 1.497188e-26, 1.881787e-26, 1.826198e-26, 
    1.850999e-26, 2.172453e-26, 2.349194e-26, 2.753834e-26, 2.676808e-26, 
    2.381392e-26, 1.801601e-26, 1.985165e-26, 1.546957e-26, 1.555985e-26, 
    1.154745e-26, 1.324868e-26, 7.714095e-27, 9.071235e-27, 5.557841e-27, 
    6.327421e-27, 5.592371e-27, 5.808434e-27, 5.589595e-27, 6.747825e-27, 
    6.232383e-27, 7.323482e-27, 1.291693e-26, 1.103096e-26, 1.733838e-26, 
    2.221506e-26, 2.597211e-26, 2.891011e-26, 2.848045e-26, 2.767445e-26, 
    2.379737e-26, 2.053435e-26, 1.827917e-26, 1.687614e-26, 1.557286e-26, 
    1.207445e-26, 1.047568e-26, 7.458528e-27, 7.94941e-27, 7.13108e-27, 
    6.407949e-27, 5.314255e-27, 5.484312e-27, 5.037651e-27, 7.151996e-27, 
    5.688164e-27, 8.239168e-27, 7.473163e-27, 1.523038e-26, 1.934353e-26, 
    2.131726e-26, 2.316506e-26, 2.815331e-26, 2.463179e-26, 2.597833e-26, 
    2.286101e-26, 2.102977e-26, 2.192141e-26, 1.683893e-26, 1.869806e-26, 
    1.038604e-26, 1.353344e-26, 6.489447e-27, 7.846828e-27, 6.191091e-27, 
    7.000753e-27, 5.656101e-27, 6.856899e-27, 4.878312e-27, 4.508938e-27, 
    4.759095e-27, 3.849466e-27, 6.928377e-27, 5.592313e-27, 2.194671e-26, 
    2.179928e-26, 2.112226e-26, 2.421854e-26, 2.441837e-26, 2.755959e-26, 
    2.475097e-26, 2.362173e-26, 2.092719e-26, 1.944423e-26, 1.810791e-26, 
    1.540859e-26, 1.275618e-26, 9.627065e-27, 7.753135e-27, 6.654693e-27, 
    7.313931e-27, 6.729604e-27, 7.385108e-27, 7.707681e-27, 4.644878e-27, 
    6.227674e-27, 3.971945e-27, 4.078476e-27, 5.027335e-27, 4.066372e-27, 
    2.169622e-26, 2.255169e-26, 2.571618e-26, 2.321365e-26, 2.791895e-26, 
    2.520567e-26, 2.373701e-26, 1.865739e-26, 1.765924e-26, 1.67689e-26, 
    1.51082e-26, 1.315742e-26, 1.018832e-26, 8.030024e-27, 6.367603e-27, 
    6.480147e-27, 6.440359e-27, 6.103088e-27, 6.962631e-27, 5.969651e-27, 
    5.813518e-27, 6.227962e-27, 4.092893e-27, 4.638627e-27, 4.080761e-27, 
    4.429839e-27, 2.227097e-26, 2.085882e-26, 2.161337e-26, 2.021066e-26, 
    2.119149e-26, 1.708477e-26, 1.59769e-26, 1.147792e-26, 1.319387e-26, 
    1.054328e-26, 1.290468e-26, 1.24606e-26, 1.046355e-26, 1.276814e-26, 
    8.139343e-27, 1.111037e-26, 6.090241e-27, 8.51859e-27, 5.956992e-27, 
    6.374206e-27, 5.694367e-27, 5.130986e-27, 4.480318e-27, 3.437075e-27, 
    3.661399e-27, 2.897441e-27, 1.887799e-26, 1.727029e-26, 1.740791e-26, 
    1.58266e-26, 1.472688e-26, 1.253673e-26, 9.533191e-27, 1.059298e-26, 
    8.708436e-27, 8.361617e-27, 1.125088e-26, 9.403505e-27, 1.625239e-26, 
    1.495583e-26, 1.571844e-26, 1.874714e-26, 1.034128e-26, 1.420027e-26, 
    7.724555e-27, 9.335163e-27, 5.208746e-27, 7.045541e-27, 3.789196e-27, 
    2.797874e-27, 2.047166e-27, 1.363264e-27, 1.643692e-26, 1.747947e-26, 
    1.564591e-26, 1.334648e-26, 1.144415e-26, 9.230498e-27, 9.023195e-27, 
    8.652165e-27, 7.742649e-27, 7.033021e-27, 8.537025e-27, 6.862764e-27, 
    1.466583e-26, 1.004719e-26, 1.788575e-26, 1.517289e-26, 1.347479e-26, 
    1.42018e-26, 1.071937e-26, 9.999059e-27, 7.42802e-27, 8.688221e-27, 
    3.022952e-27, 5.01714e-27, 9.635816e-28, 1.6674e-27, 1.785486e-26, 
    1.644056e-26, 1.215173e-26, 1.407438e-26, 9.094884e-27, 8.098812e-27, 
    7.349305e-27, 6.465401e-27, 6.374884e-27, 5.893745e-27, 6.696527e-27, 
    5.92412e-27, 9.226149e-27, 7.620265e-27, 1.259516e-26, 1.121448e-26, 
    1.183522e-26, 1.254434e-26, 1.04503e-26, 8.511654e-27, 8.473589e-27, 
    7.913165e-27, 6.477347e-27, 9.077815e-27, 2.814999e-27, 6.065961e-27, 
    1.499404e-26, 1.266924e-26, 1.236056e-26, 1.321183e-26, 8.194924e-27, 
    9.814418e-27, 5.90518e-27, 6.823699e-27, 5.367384e-27, 6.059728e-27, 
    6.166716e-27, 7.159307e-27, 7.832373e-27, 9.735419e-27, 1.151489e-26, 
    1.308584e-26, 1.270744e-26, 1.102666e-26, 8.402315e-27, 6.366633e-27, 
    6.77819e-27, 5.469405e-27, 9.404424e-27, 7.567001e-27, 8.243016e-27, 
    6.565438e-27, 1.062219e-26, 7.08046e-27, 1.170184e-26, 1.122755e-26, 
    9.84874e-27, 7.452461e-27, 6.985806e-27, 6.51076e-27, 6.801092e-27, 
    8.342318e-27, 8.617018e-27, 9.880783e-27, 1.025201e-26, 1.132962e-26, 
    1.228213e-26, 1.140958e-26, 1.05427e-26, 8.341727e-27, 6.661651e-27, 
    5.123239e-27, 4.789569e-27, 3.405505e-27, 4.506218e-27, 2.801513e-27, 
    4.213175e-27, 2.00872e-27, 6.906212e-27, 4.261368e-27, 9.789184e-27, 
    9.028932e-27, 7.763454e-27, 5.349399e-27, 6.572697e-27, 5.159659e-27, 
    8.627932e-27, 1.097157e-26, 1.164677e-26, 1.298604e-26, 1.161738e-26, 
    1.172459e-26, 1.050809e-26, 1.088849e-26, 8.274931e-27, 9.614128e-27, 
    6.169365e-27, 5.169923e-27, 2.971612e-27, 2.011939e-27, 1.282918e-27, 
    1.029513e-27, 9.598902e-28, 9.317748e-28,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.004414367, 0.004411613, 0.00441215, 0.004409926, 0.004411161, 
    0.004409705, 0.004413811, 0.004411502, 0.004412977, 0.004414122, 
    0.00440561, 0.004409828, 0.004401256, 0.004403939, 0.004397211, 
    0.00440167, 0.004396313, 0.004397345, 0.004394255, 0.00439514, 
    0.004391179, 0.004393846, 0.004389137, 0.004391819, 0.004391397, 
    0.004393933, 0.004408984, 0.004406133, 0.004409152, 0.004408745, 
    0.004408929, 0.004411134, 0.004412243, 0.004414581, 0.004414157, 
    0.004412442, 0.004408563, 0.004409882, 0.004406567, 0.004406642, 
    0.004402952, 0.004404615, 0.004398422, 0.004400183, 0.004395103, 
    0.004396379, 0.004395162, 0.004395531, 0.004395157, 0.004397029, 
    0.004396227, 0.004397876, 0.004404303, 0.004402411, 0.004408053, 
    0.004411443, 0.004413709, 0.004415313, 0.004415086, 0.004414653, 
    0.004412432, 0.004410349, 0.004408761, 0.004407699, 0.004406653, 
    0.004403476, 0.004401807, 0.004398064, 0.004398744, 0.004397596, 
    0.004396506, 0.004394671, 0.004394974, 0.004394165, 0.004397629, 
    0.004395325, 0.00439913, 0.004398088, 0.004406351, 0.004409527, 
    0.004410863, 0.004412046, 0.004414911, 0.004412931, 0.004413711, 
    0.004411859, 0.00441068, 0.004411264, 0.00440767, 0.004409066, 
    0.004401708, 0.004404875, 0.004396633, 0.004398604, 0.004396162, 
    0.004397409, 0.004395271, 0.004397195, 0.004393865, 0.004393138, 
    0.004393635, 0.004391735, 0.004397301, 0.00439516, 0.00441128, 
    0.004411184, 0.004410742, 0.004412685, 0.004412805, 0.004414592, 
    0.004413004, 0.004412326, 0.004410614, 0.004409598, 0.004408634, 
    0.004406515, 0.004404147, 0.004400844, 0.004398476, 0.004396889, 
    0.004397864, 0.004397003, 0.004397964, 0.004398416, 0.00439341, 
    0.004396218, 0.004392009, 0.004392242, 0.004394145, 0.004392216, 
    0.004411118, 0.004411666, 0.004413563, 0.004412078, 0.004414787, 
    0.004413268, 0.004412394, 0.004409033, 0.004408299, 0.004407614, 
    0.004406264, 0.00440453, 0.00440149, 0.004398849, 0.004396444, 
    0.00439662, 0.004396558, 0.004396019, 0.004397352, 0.0043958, 
    0.004395538, 0.004396221, 0.004392273, 0.004393401, 0.004392247, 
    0.004392982, 0.004411488, 0.004410567, 0.004411065, 0.004410128, 
    0.004410786, 0.004407856, 0.004406977, 0.004402876, 0.004404563, 
    0.004401884, 0.004404292, 0.004403864, 0.004401789, 0.004404163, 
    0.004398991, 0.00440249, 0.004395998, 0.004399481, 0.004395779, 
    0.004396454, 0.004395339, 0.004394338, 0.004393084, 0.004390764, 
    0.004391302, 0.004389366, 0.004409196, 0.004408001, 0.004408109, 
    0.004406861, 0.004405937, 0.00440394, 0.004400736, 0.004401942, 
    0.004399732, 0.004399288, 0.004402646, 0.004400581, 0.004407203, 
    0.004406129, 0.004406771, 0.0044091, 0.004401659, 0.004405473, 
    0.004398437, 0.004400501, 0.00439448, 0.00439747, 0.004391597, 
    0.004389081, 0.00438673, 0.004383965, 0.004407352, 0.004408163, 
    0.004406713, 0.004404702, 0.004402846, 0.004400374, 0.004400124, 
    0.00439966, 0.004398463, 0.004397456, 0.00439951, 0.004397204, 
    0.004405873, 0.00440133, 0.004408468, 0.004406312, 0.004404822, 
    0.004405479, 0.00440208, 0.004401279, 0.004398022, 0.004399707, 
    0.004389699, 0.004394122, 0.004381874, 0.00438529, 0.004408447, 
    0.004407356, 0.00440356, 0.004405366, 0.004400211, 0.004398942, 
    0.004397914, 0.004396594, 0.004396454, 0.004395674, 0.004396953, 
    0.004395725, 0.004400369, 0.004398294, 0.004403998, 0.004402606, 
    0.004403247, 0.004403948, 0.004401785, 0.004399477, 0.004399433, 
    0.004398692, 0.004396596, 0.004400191, 0.004389118, 0.004395942, 
    0.004406168, 0.004404062, 0.004403768, 0.004404582, 0.00439907, 
    0.004401065, 0.004395693, 0.004397145, 0.004394768, 0.004395948, 
    0.004396122, 0.00439764, 0.004398585, 0.004400973, 0.004402918, 
    0.004404465, 0.004404105, 0.004402407, 0.004399337, 0.00439644, 
    0.004397073, 0.004394948, 0.004400585, 0.004398217, 0.00439913, 
    0.004396751, 0.004401973, 0.004397509, 0.004403112, 0.004402622, 
    0.004401105, 0.004398053, 0.004397386, 0.004396665, 0.004397111, 
    0.00439926, 0.004399615, 0.004401143, 0.004401562, 0.004402729, 
    0.004403693, 0.004402811, 0.004401884, 0.004399261, 0.004396897, 
    0.004394323, 0.004393696, 0.004390678, 0.004393127, 0.004389079, 
    0.004392509, 0.004386579, 0.004397259, 0.004392621, 0.004401037, 
    0.004400131, 0.004398486, 0.004394729, 0.004396762, 0.004394387, 
    0.004399629, 0.004402346, 0.004403056, 0.00440437, 0.004403026, 
    0.004403135, 0.00440185, 0.004402263, 0.004399174, 0.004400834, 
    0.004396125, 0.004394407, 0.004389567, 0.004386599, 0.00438359, 
    0.004382259, 0.004381855, 0.004381685,
  8.312036e-06, 8.311841e-06, 8.311886e-06, 8.311705e-06, 8.311816e-06, 
    8.311687e-06, 8.312009e-06, 8.311823e-06, 8.311949e-06, 8.312034e-06, 
    8.311284e-06, 8.311698e-06, 8.310906e-06, 8.31119e-06, 8.310472e-06, 
    8.310936e-06, 8.310377e-06, 8.310511e-06, 8.310158e-06, 8.310263e-06, 
    8.309733e-06, 8.310109e-06, 8.309481e-06, 8.309838e-06, 8.309774e-06, 
    8.310117e-06, 8.311642e-06, 8.31133e-06, 8.311655e-06, 8.311613e-06, 
    8.311637e-06, 8.311805e-06, 8.311869e-06, 8.312067e-06, 8.312036e-06, 
    8.311899e-06, 8.311595e-06, 8.311718e-06, 8.311445e-06, 8.311452e-06, 
    8.311097e-06, 8.311261e-06, 8.31063e-06, 8.310825e-06, 8.31026e-06, 
    8.310404e-06, 8.310262e-06, 8.310309e-06, 8.310261e-06, 8.310473e-06, 
    8.310382e-06, 8.310573e-06, 8.311226e-06, 8.311038e-06, 8.311559e-06, 
    8.311796e-06, 8.311997e-06, 8.312112e-06, 8.312097e-06, 8.31206e-06, 
    8.311898e-06, 8.311756e-06, 8.311631e-06, 8.311541e-06, 8.311452e-06, 
    8.311104e-06, 8.310962e-06, 8.310578e-06, 8.31067e-06, 8.310529e-06, 
    8.31042e-06, 8.310201e-06, 8.31024e-06, 8.310138e-06, 8.310547e-06, 
    8.310271e-06, 8.310718e-06, 8.310597e-06, 8.311345e-06, 8.311689e-06, 
    8.311757e-06, 8.311874e-06, 8.312082e-06, 8.311937e-06, 8.311993e-06, 
    8.311873e-06, 8.31178e-06, 8.31183e-06, 8.311538e-06, 8.311653e-06, 
    8.310953e-06, 8.311273e-06, 8.310432e-06, 8.310653e-06, 8.310381e-06, 
    8.310526e-06, 8.310269e-06, 8.310501e-06, 8.310106e-06, 8.310006e-06, 
    8.310072e-06, 8.309842e-06, 8.310511e-06, 8.310254e-06, 8.311828e-06, 
    8.311818e-06, 8.311788e-06, 8.311917e-06, 8.311929e-06, 8.312063e-06, 
    8.311952e-06, 8.311896e-06, 8.311781e-06, 8.311694e-06, 8.311615e-06, 
    8.311432e-06, 8.3112e-06, 8.310876e-06, 8.310638e-06, 8.310467e-06, 
    8.310578e-06, 8.31048e-06, 8.310586e-06, 8.31064e-06, 8.310038e-06, 
    8.310377e-06, 8.309876e-06, 8.309908e-06, 8.310132e-06, 8.309904e-06, 
    8.311814e-06, 8.31186e-06, 8.311989e-06, 8.311889e-06, 8.312079e-06, 
    8.311965e-06, 8.31189e-06, 8.311632e-06, 8.311591e-06, 8.311526e-06, 
    8.311414e-06, 8.311253e-06, 8.310944e-06, 8.310671e-06, 8.310417e-06, 
    8.310438e-06, 8.31043e-06, 8.310362e-06, 8.310516e-06, 8.310337e-06, 
    8.310299e-06, 8.310387e-06, 8.309911e-06, 8.310052e-06, 8.309908e-06, 
    8.310002e-06, 8.311848e-06, 8.311773e-06, 8.311812e-06, 8.311733e-06, 
    8.311782e-06, 8.311529e-06, 8.311448e-06, 8.311069e-06, 8.311251e-06, 
    8.310981e-06, 8.311231e-06, 8.311183e-06, 8.310937e-06, 8.311224e-06, 
    8.310671e-06, 8.311022e-06, 8.31036e-06, 8.310704e-06, 8.310335e-06, 
    8.310418e-06, 8.310289e-06, 8.31016e-06, 8.310011e-06, 8.309702e-06, 
    8.309778e-06, 8.309525e-06, 8.311664e-06, 8.311552e-06, 8.311577e-06, 
    8.311466e-06, 8.311379e-06, 8.311201e-06, 8.310874e-06, 8.311005e-06, 
    8.31078e-06, 8.310727e-06, 8.311078e-06, 8.310851e-06, 8.311486e-06, 
    8.311375e-06, 8.311453e-06, 8.311647e-06, 8.310953e-06, 8.311317e-06, 
    8.310632e-06, 8.310853e-06, 8.310177e-06, 8.310509e-06, 8.309816e-06, 
    8.309452e-06, 8.310021e-06, 8.310609e-06, 8.311506e-06, 8.311582e-06, 
    8.311457e-06, 8.311248e-06, 8.311088e-06, 8.310838e-06, 8.31082e-06, 
    8.310766e-06, 8.310643e-06, 8.31053e-06, 8.310733e-06, 8.310502e-06, 
    8.311317e-06, 8.310928e-06, 8.311596e-06, 8.311388e-06, 8.311267e-06, 
    8.311337e-06, 8.311024e-06, 8.31094e-06, 8.310577e-06, 8.310777e-06, 
    8.309529e-06, 8.310111e-06, 8.311093e-06, 8.310321e-06, 8.311605e-06, 
    8.311513e-06, 8.311148e-06, 8.311329e-06, 8.310829e-06, 8.310688e-06, 
    8.310584e-06, 8.310421e-06, 8.310415e-06, 8.310319e-06, 8.310474e-06, 
    8.31033e-06, 8.310837e-06, 8.31062e-06, 8.31121e-06, 8.311065e-06, 
    8.311138e-06, 8.311205e-06, 8.310992e-06, 8.310727e-06, 8.310746e-06, 
    8.310653e-06, 8.31034e-06, 8.310827e-06, 8.309404e-06, 8.310277e-06, 
    8.311408e-06, 8.311183e-06, 8.31118e-06, 8.311264e-06, 8.310702e-06, 
    8.310911e-06, 8.310324e-06, 8.310496e-06, 8.310219e-06, 8.310356e-06, 
    8.310375e-06, 8.310551e-06, 8.310651e-06, 8.310897e-06, 8.311094e-06, 
    8.311255e-06, 8.31122e-06, 8.311041e-06, 8.310715e-06, 8.310403e-06, 
    8.31047e-06, 8.31024e-06, 8.310866e-06, 8.310601e-06, 8.310697e-06, 
    8.310447e-06, 8.311003e-06, 8.310458e-06, 8.311125e-06, 8.311075e-06, 
    8.310915e-06, 8.310565e-06, 8.310522e-06, 8.31043e-06, 8.310492e-06, 
    8.310712e-06, 8.310758e-06, 8.310925e-06, 8.310958e-06, 8.311088e-06, 
    8.311181e-06, 8.31109e-06, 8.310986e-06, 8.310722e-06, 8.310454e-06, 
    8.310155e-06, 8.310089e-06, 8.309649e-06, 8.309974e-06, 8.309394e-06, 
    8.309838e-06, 8.30998e-06, 8.310461e-06, 8.309901e-06, 8.310916e-06, 
    8.310822e-06, 8.310619e-06, 8.31018e-06, 8.310448e-06, 8.310147e-06, 
    8.310762e-06, 8.311022e-06, 8.311118e-06, 8.311241e-06, 8.311114e-06, 
    8.311126e-06, 8.311e-06, 8.311043e-06, 8.310713e-06, 8.310894e-06, 
    8.310369e-06, 8.310155e-06, 8.309542e-06, 8.310021e-06, 8.310731e-06, 
    8.311021e-06, 8.31111e-06, 8.311145e-06,
  1.680188e-10, 1.68097e-10, 1.680819e-10, 1.681448e-10, 1.681102e-10, 
    1.681512e-10, 1.68035e-10, 1.680998e-10, 1.680586e-10, 1.680263e-10, 
    1.682666e-10, 1.681477e-10, 1.683944e-10, 1.683172e-10, 1.685127e-10, 
    1.683819e-10, 1.685393e-10, 1.685097e-10, 1.68601e-10, 1.685748e-10, 
    1.686905e-10, 1.68613e-10, 1.68752e-10, 1.686724e-10, 1.686845e-10, 
    1.686104e-10, 1.681723e-10, 1.682515e-10, 1.681674e-10, 1.681787e-10, 
    1.681738e-10, 1.681106e-10, 1.680784e-10, 1.680134e-10, 1.680253e-10, 
    1.680733e-10, 1.681838e-10, 1.681467e-10, 1.682419e-10, 1.682398e-10, 
    1.683459e-10, 1.682979e-10, 1.68478e-10, 1.684268e-10, 1.685759e-10, 
    1.685382e-10, 1.68574e-10, 1.685632e-10, 1.685741e-10, 1.685189e-10, 
    1.685425e-10, 1.684942e-10, 1.683068e-10, 1.683614e-10, 1.681987e-10, 
    1.681006e-10, 1.680377e-10, 1.679926e-10, 1.67999e-10, 1.68011e-10, 
    1.680736e-10, 1.681334e-10, 1.681789e-10, 1.682093e-10, 1.682394e-10, 
    1.68329e-10, 1.683783e-10, 1.68488e-10, 1.684688e-10, 1.685019e-10, 
    1.685344e-10, 1.685884e-10, 1.685796e-10, 1.686032e-10, 1.685015e-10, 
    1.685688e-10, 1.684577e-10, 1.68488e-10, 1.682451e-10, 1.681568e-10, 
    1.681173e-10, 1.680847e-10, 1.680038e-10, 1.680595e-10, 1.680375e-10, 
    1.680905e-10, 1.681239e-10, 1.681075e-10, 1.682101e-10, 1.6817e-10, 
    1.683813e-10, 1.682899e-10, 1.685306e-10, 1.684728e-10, 1.685446e-10, 
    1.685081e-10, 1.685705e-10, 1.685143e-10, 1.686122e-10, 1.686334e-10, 
    1.686189e-10, 1.686754e-10, 1.685111e-10, 1.685737e-10, 1.681069e-10, 
    1.681096e-10, 1.681223e-10, 1.680664e-10, 1.680631e-10, 1.680129e-10, 
    1.680578e-10, 1.680768e-10, 1.68126e-10, 1.681548e-10, 1.681823e-10, 
    1.682431e-10, 1.683108e-10, 1.684068e-10, 1.684765e-10, 1.685233e-10, 
    1.684948e-10, 1.685199e-10, 1.684917e-10, 1.684786e-10, 1.686253e-10, 
    1.685425e-10, 1.686673e-10, 1.686605e-10, 1.686037e-10, 1.686612e-10, 
    1.681115e-10, 1.680961e-10, 1.680419e-10, 1.680843e-10, 1.680075e-10, 
    1.680501e-10, 1.680745e-10, 1.681703e-10, 1.681921e-10, 1.682115e-10, 
    1.682505e-10, 1.683004e-10, 1.683881e-10, 1.684653e-10, 1.685364e-10, 
    1.685313e-10, 1.685331e-10, 1.685487e-10, 1.685096e-10, 1.685552e-10, 
    1.685626e-10, 1.685428e-10, 1.686595e-10, 1.686261e-10, 1.686603e-10, 
    1.686386e-10, 1.681011e-10, 1.681272e-10, 1.681131e-10, 1.681395e-10, 
    1.681207e-10, 1.682039e-10, 1.682289e-10, 1.683473e-10, 1.682992e-10, 
    1.683765e-10, 1.683073e-10, 1.683194e-10, 1.68378e-10, 1.683112e-10, 
    1.684606e-10, 1.683582e-10, 1.685493e-10, 1.684455e-10, 1.685558e-10, 
    1.685361e-10, 1.68569e-10, 1.685982e-10, 1.686355e-10, 1.687037e-10, 
    1.68688e-10, 1.687457e-10, 1.681664e-10, 1.682001e-10, 1.681976e-10, 
    1.682333e-10, 1.682597e-10, 1.683176e-10, 1.684103e-10, 1.683755e-10, 
    1.6844e-10, 1.684528e-10, 1.683552e-10, 1.684146e-10, 1.682231e-10, 
    1.682534e-10, 1.682357e-10, 1.681687e-10, 1.683829e-10, 1.682723e-10, 
    1.684776e-10, 1.684173e-10, 1.68594e-10, 1.685054e-10, 1.686793e-10, 
    1.687529e-10, 1.688476e-10, 1.689567e-10, 1.68219e-10, 1.68196e-10, 
    1.682377e-10, 1.682947e-10, 1.68349e-10, 1.684209e-10, 1.684285e-10, 
    1.684419e-10, 1.684772e-10, 1.685066e-10, 1.684457e-10, 1.685141e-10, 
    1.682594e-10, 1.683928e-10, 1.681869e-10, 1.68248e-10, 1.682915e-10, 
    1.682729e-10, 1.683717e-10, 1.683949e-10, 1.684894e-10, 1.684408e-10, 
    1.687342e-10, 1.686037e-10, 1.690416e-10, 1.689041e-10, 1.681879e-10, 
    1.682192e-10, 1.68328e-10, 1.682762e-10, 1.68426e-10, 1.684628e-10, 
    1.684933e-10, 1.685315e-10, 1.68536e-10, 1.685588e-10, 1.685214e-10, 
    1.685575e-10, 1.684211e-10, 1.68482e-10, 1.683161e-10, 1.68356e-10, 
    1.683378e-10, 1.683175e-10, 1.683802e-10, 1.684465e-10, 1.684487e-10, 
    1.684699e-10, 1.685284e-10, 1.684266e-10, 1.687497e-10, 1.685481e-10, 
    1.682534e-10, 1.683129e-10, 1.683224e-10, 1.682991e-10, 1.684591e-10, 
    1.684008e-10, 1.685583e-10, 1.685158e-10, 1.685858e-10, 1.685509e-10, 
    1.685457e-10, 1.685012e-10, 1.684734e-10, 1.684034e-10, 1.683469e-10, 
    1.683026e-10, 1.683129e-10, 1.683616e-10, 1.684508e-10, 1.685361e-10, 
    1.685172e-10, 1.685804e-10, 1.68415e-10, 1.684838e-10, 1.684569e-10, 
    1.685272e-10, 1.683745e-10, 1.685021e-10, 1.683417e-10, 1.683559e-10, 
    1.683997e-10, 1.684879e-10, 1.685087e-10, 1.685295e-10, 1.685168e-10, 
    1.684532e-10, 1.684431e-10, 1.683988e-10, 1.683862e-10, 1.683528e-10, 
    1.683249e-10, 1.683503e-10, 1.683767e-10, 1.684535e-10, 1.685226e-10, 
    1.685985e-10, 1.686174e-10, 1.687047e-10, 1.686326e-10, 1.687507e-10, 
    1.686486e-10, 1.688508e-10, 1.685107e-10, 1.686472e-10, 1.68402e-10, 
    1.684284e-10, 1.684755e-10, 1.685856e-10, 1.685269e-10, 1.68596e-10, 
    1.684428e-10, 1.683629e-10, 1.683433e-10, 1.683051e-10, 1.683442e-10, 
    1.68341e-10, 1.683784e-10, 1.683664e-10, 1.684561e-10, 1.684079e-10, 
    1.685454e-10, 1.685956e-10, 1.687393e-10, 1.688517e-10, 1.689733e-10, 
    1.690266e-10, 1.690429e-10, 1.690497e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  1.024205, 1.004775, 1.008553, 0.9928728, 1.001573, 0.9913033, 1.020268, 
    1.004002, 1.014387, 1.022458, 0.9624152, 0.9921733, 0.9314803, 0.9504818, 
    0.9027274, 0.9344367, 0.8963296, 0.9036449, 0.8816274, 0.8879369, 
    0.8597513, 0.8787149, 0.8451329, 0.8642825, 0.8612868, 0.8793399, 
    0.9861892, 0.9661211, 0.9873773, 0.9845167, 0.9858008, 1.001393, 
    1.009245, 1.025691, 1.022707, 1.010628, 0.9832303, 0.9925349, 0.9690835, 
    0.9696134, 0.9434814, 0.9552667, 0.91131, 0.9238108, 0.8876737, 
    0.8967658, 0.8881004, 0.8907286, 0.8880662, 0.9013998, 0.8956877, 
    0.9074184, 0.9530594, 0.9396528, 0.9796179, 1.003618, 1.019554, 1.030856, 
    1.029258, 1.026212, 1.010557, 0.9958328, 0.984606, 0.9770934, 0.9696895, 
    0.947261, 0.9353878, 0.9087805, 0.913586, 0.9054461, 0.8976703, 
    0.8846079, 0.8867586, 0.8810017, 0.9056623, 0.8892745, 0.9163225, 
    0.908927, 0.9676688, 0.9900254, 0.9995162, 1.007827, 1.02803, 1.014079, 
    1.019579, 1.006494, 0.9981754, 1.00229, 0.9768879, 0.986766, 0.9346839, 
    0.9571292, 0.8985773, 0.9125999, 0.8952156, 0.9040881, 0.8888831, 
    0.9025679, 0.8788594, 0.8736933, 0.8772236, 0.8636628, 0.9033261, 
    0.8880997, 1.002405, 1.001734, 0.9986082, 1.012346, 1.013187, 1.025773, 
    1.014575, 1.009804, 0.9976937, 0.9905266, 0.9837123, 0.9687244, 
    0.9519749, 0.928539, 0.9116911, 0.9003916, 0.9073213, 0.9012033, 
    0.9080421, 0.9112473, 0.8756287, 0.8956339, 0.8656136, 0.867276, 
    0.8808644, 0.8670886, 1.001263, 1.005124, 1.018525, 1.008039, 1.027143, 
    1.01645, 1.010299, 0.986558, 0.9813411, 0.9765005, 0.9669394, 0.9546636, 
    0.9331154, 0.9143545, 0.8972182, 0.8984743, 0.898032, 0.8942017, 
    0.9036875, 0.8926442, 0.8907896, 0.8956373, 0.8674985, 0.8755406, 
    0.8673112, 0.872548, 1.00387, 0.9973717, 1.000883, 0.9942795, 0.9989312, 
    0.9782391, 0.9720324, 0.9429735, 0.9549049, 0.9359157, 0.9529771, 
    0.9499543, 0.9352928, 0.9520559, 0.9153878, 0.94025, 0.8940528, 
    0.9188961, 0.8924951, 0.8972923, 0.8893501, 0.882234, 0.8732806, 
    0.8567502, 0.8605793, 0.8467507, 0.9876829, 0.9792492, 0.9799932, 
    0.971166, 0.9646356, 0.950478, 0.9277546, 0.9363022, 0.9206098, 
    0.9174579, 0.9412987, 0.9266618, 0.9736047, 0.9660242, 0.9705389, 
    0.9870169, 0.9343308, 0.9613808, 0.9114122, 0.9260815, 0.8832486, 
    0.9045569, 0.8626865, 0.844764, 0.8278925, 0.8081549, 0.9746469, 
    0.9803784, 0.9701164, 0.9559097, 0.9427258, 0.9251867, 0.9233924, 
    0.9201047, 0.9115888, 0.904426, 0.9190637, 0.9026303, 0.964263, 
    0.9319823, 0.9825437, 0.9673261, 0.956748, 0.9613903, 0.9372793, 
    0.9315932, 0.9084743, 0.9204286, 0.8491872, 0.8807287, 0.7931225, 
    0.8176312, 0.9823804, 0.9746673, 0.9478049, 0.9605895, 0.9240162, 
    0.9150059, 0.9076802, 0.8983106, 0.8972999, 0.8917469, 0.9008457, 
    0.892107, 0.9251493, 0.9103884, 0.9508784, 0.9410279, 0.9455605, 
    0.9505302, 0.9351889, 0.918833, 0.9184858, 0.9132386, 0.8984433, 
    0.923868, 0.8451091, 0.8937709, 0.9662542, 0.9513842, 0.9492624, 
    0.9550235, 0.9159092, 0.9300877, 0.8918827, 0.9022138, 0.885285, 
    0.8936983, 0.8949358, 0.9057378, 0.9124602, 0.9294373, 0.9432438, 
    0.9541883, 0.951644, 0.9396204, 0.9178327, 0.8972073, 0.9017264, 
    0.886572, 0.9266696, 0.9098616, 0.9163584, 0.8994157, 0.9365288, 
    0.9049209, 0.9446015, 0.9411252, 0.9303691, 0.9087197, 0.9039312, 
    0.8988132, 0.9019719, 0.9172798, 0.919788, 0.9306312, 0.9336231, 
    0.9418823, 0.9487171, 0.9424718, 0.9359112, 0.9172744, 0.9004673, 
    0.8821324, 0.8776445, 0.8561971, 0.8736542, 0.8448374, 0.8693339, 
    0.8269178, 0.9030917, 0.8700589, 0.9298804, 0.9234424, 0.9117916, 
    0.8850564, 0.8994955, 0.8826094, 0.9198865, 0.9392043, 0.9442032, 
    0.9535226, 0.9439901, 0.9447656, 0.9356411, 0.9385737, 0.9166554, 
    0.9284312, 0.8949662, 0.8827434, 0.8481994, 0.827, 0.8054078, 0.7958688, 
    0.7929651, 0.7917509,
  0.4113339, 0.3957348, 0.3987494, 0.3863026, 0.3931887, 0.3850658, 
    0.4081534, 0.3951194, 0.4034216, 0.4099215, 0.3625988, 0.3857512, 
    0.339186, 0.3534888, 0.3180384, 0.341394, 0.3134156, 0.3187046, 0.302908, 
    0.3073978, 0.2875732, 0.3008455, 0.2775321, 0.29072, 0.288638, 0.3012875, 
    0.3810479, 0.3654487, 0.3819798, 0.3797372, 0.3807434, 0.3930451, 
    0.3993014, 0.4125376, 0.4101226, 0.4004079, 0.3787306, 0.3860368, 
    0.3677364, 0.3681458, 0.34819, 0.3571308, 0.3242885, 0.3334874, 
    0.3072099, 0.3137304, 0.3075145, 0.3093939, 0.30749, 0.3170773, 
    0.3129538, 0.3214482, 0.3554487, 0.3453064, 0.3759103, 0.3948132, 
    0.4075778, 0.4167297, 0.4154311, 0.4129593, 0.4003513, 0.3886401, 
    0.3798077, 0.3739448, 0.3682046, 0.3510451, 0.3421061, 0.3224406, 
    0.3259549, 0.3200125, 0.3143825, 0.3050249, 0.3065569, 0.302464, 
    0.3201702, 0.308353, 0.3279636, 0.3225479, 0.3666416, 0.3840607, 
    0.391555, 0.3981688, 0.4144335, 0.4031737, 0.4075978, 0.3971057, 
    0.3904938, 0.3937588, 0.3737851, 0.3815004, 0.3415793, 0.3585522, 
    0.3150369, 0.3252324, 0.3126143, 0.3190266, 0.3080734, 0.3179237, 
    0.3009475, 0.2973042, 0.2997917, 0.2902892, 0.3184735, 0.3075137, 
    0.39385, 0.3933167, 0.3908368, 0.4017839, 0.402458, 0.4126034, 0.403572, 
    0.3997491, 0.3901126, 0.384455, 0.3791081, 0.3674588, 0.3546231, 
    0.3369955, 0.3245672, 0.316348, 0.3213777, 0.3169353, 0.3219028, 
    0.3242429, 0.2986665, 0.312915, 0.2916476, 0.2928074, 0.3023667, 
    0.2926766, 0.3929425, 0.3960142, 0.4067488, 0.3983384, 0.4137143, 
    0.4050784, 0.4001445, 0.3813366, 0.3772551, 0.3734835, 0.3660819, 
    0.3566708, 0.3404071, 0.3265181, 0.3140566, 0.3149627, 0.3146435, 
    0.3118852, 0.3187357, 0.3107668, 0.3094372, 0.3129177, 0.2929628, 
    0.2986049, 0.2928321, 0.2964997, 0.3950149, 0.3898575, 0.3926409, 
    0.3874129, 0.3910924, 0.3748356, 0.3700158, 0.3478062, 0.3568546, 
    0.3425018, 0.3553862, 0.3530883, 0.3420343, 0.3546854, 0.3272759, 
    0.3457546, 0.3117782, 0.3298559, 0.3106599, 0.31411, 0.3084075, 
    0.3033381, 0.2970144, 0.2854989, 0.2881478, 0.2786356, 0.3822199, 
    0.3756228, 0.3762034, 0.3693462, 0.3643075, 0.3534863, 0.3364127, 
    0.3427921, 0.3311211, 0.3287983, 0.3465452, 0.3356007, 0.3712349, 
    0.3653756, 0.3688608, 0.3816969, 0.3413154, 0.3618066, 0.3243632, 
    0.3351703, 0.3040585, 0.3193662, 0.2896102, 0.2772802, 0.2659042, 
    0.2528791, 0.3720437, 0.3765039, 0.3685346, 0.3576207, 0.3476202, 
    0.3345065, 0.3331777, 0.3307483, 0.3244927, 0.3192719, 0.3299802, 
    0.317969, 0.3640189, 0.339561, 0.3781942, 0.3663789, 0.358261, 0.3618146, 
    0.3435248, 0.3392712, 0.3222174, 0.3309875, 0.2802997, 0.3022699, 
    0.2431699, 0.2590936, 0.3780669, 0.3720598, 0.3514583, 0.3612006, 
    0.3336395, 0.3269962, 0.3216392, 0.3148441, 0.3141154, 0.3101233, 
    0.3166765, 0.3103816, 0.3344788, 0.323615, 0.3537905, 0.3463411, 
    0.3497605, 0.353526, 0.3419583, 0.32981, 0.329555, 0.3257, 0.3149374, 
    0.3335297, 0.2775138, 0.3115733, 0.3655539, 0.3541737, 0.3525635, 
    0.3569455, 0.3276596, 0.3381488, 0.3102207, 0.3176671, 0.3055071, 
    0.3115236, 0.312413, 0.3202252, 0.3251302, 0.3376643, 0.3480107, 
    0.3563089, 0.3543723, 0.3452822, 0.3290736, 0.3140483, 0.3173135, 
    0.306424, 0.3356069, 0.3232298, 0.3279893, 0.3156424, 0.3429617, 
    0.3196289, 0.3490359, 0.3464146, 0.3383584, 0.3223959, 0.3189126, 
    0.315207, 0.3174919, 0.3286669, 0.3305146, 0.3385539, 0.3407867, 
    0.3469848, 0.3521503, 0.3474289, 0.3424987, 0.3286632, 0.3164023, 
    0.3032658, 0.3000891, 0.2851161, 0.2972758, 0.2773286, 0.2942432, 
    0.2652518, 0.318302, 0.2947522, 0.3379946, 0.3332148, 0.3246401, 
    0.3053433, 0.3157, 0.3036039, 0.3305872, 0.344969, 0.3487351, 0.3558016, 
    0.3485742, 0.3491598, 0.3422969, 0.3444963, 0.328208, 0.336916, 
    0.3124347, 0.3036993, 0.2796249, 0.2653078, 0.2510919, 0.2449303, 
    0.2430694, 0.2422932,
  0.1873237, 0.1793951, 0.180924, 0.1746218, 0.1781051, 0.1739971, 0.1857037, 
    0.1790832, 0.1832968, 0.1866041, 0.1626971, 0.1743432, 0.151022, 
    0.1581418, 0.1405686, 0.1521185, 0.1382955, 0.1408965, 0.1331453, 
    0.1353432, 0.1256713, 0.1321372, 0.120805, 0.1272008, 0.1261886, 
    0.1323532, 0.1719694, 0.1641253, 0.1724395, 0.1713086, 0.1718159, 
    0.1780323, 0.1812042, 0.1879372, 0.1867065, 0.1817659, 0.1708013, 
    0.1744875, 0.1652729, 0.1654783, 0.1554995, 0.159961, 0.1436487, 
    0.1481963, 0.1352511, 0.1384502, 0.1354003, 0.1363216, 0.1353883, 
    0.1400956, 0.1380687, 0.142248, 0.1591205, 0.1540638, 0.169381, 
    0.1789281, 0.1854107, 0.190076, 0.1894131, 0.1881523, 0.1817372, 
    0.1758032, 0.1713442, 0.1683921, 0.1655078, 0.1569226, 0.1524724, 
    0.1427372, 0.1444713, 0.1415406, 0.1387706, 0.1341811, 0.1349312, 
    0.1329283, 0.1416183, 0.1358113, 0.1454635, 0.1427901, 0.1647236, 
    0.1734895, 0.1772779, 0.1806295, 0.1889041, 0.1831708, 0.1854209, 
    0.1800902, 0.1767408, 0.1783938, 0.1683117, 0.1721977, 0.1522106, 
    0.1606717, 0.1390922, 0.1441146, 0.1379019, 0.141055, 0.1356742, 
    0.1405121, 0.132187, 0.1304083, 0.1316224, 0.1269913, 0.1407827, 0.1354, 
    0.17844, 0.1781699, 0.1769144, 0.1824647, 0.1828071, 0.1879708, 
    0.1833732, 0.1814314, 0.176548, 0.1736886, 0.1709916, 0.1651335, 
    0.1587081, 0.1499351, 0.1437862, 0.1397369, 0.1422132, 0.1400258, 
    0.1424721, 0.1436262, 0.1310731, 0.1380496, 0.1276521, 0.1282167, 
    0.1328807, 0.128153, 0.1779804, 0.1795367, 0.1849888, 0.1807155, 
    0.1885373, 0.1841391, 0.1816321, 0.172115, 0.1700581, 0.1681601, 
    0.1644428, 0.1597311, 0.1516283, 0.1447494, 0.1386104, 0.1390557, 
    0.1388988, 0.137544, 0.1409118, 0.1369951, 0.1363429, 0.1380509, 
    0.1282924, 0.131043, 0.1282287, 0.1300159, 0.1790302, 0.1764189, 
    0.1778276, 0.1751828, 0.1770438, 0.1688402, 0.1664173, 0.1553083, 
    0.159823, 0.1526691, 0.1590892, 0.1579419, 0.1524367, 0.1587392, 
    0.1451237, 0.1542869, 0.1374915, 0.146399, 0.1369426, 0.1386367, 
    0.135838, 0.1333557, 0.1302669, 0.1246642, 0.1259504, 0.1213387, 
    0.1725606, 0.1692363, 0.1695286, 0.1660809, 0.1635532, 0.1581405, 
    0.149646, 0.1528133, 0.1470249, 0.1458761, 0.1546804, 0.1492435, 
    0.1670297, 0.1640887, 0.1658373, 0.1722967, 0.1520794, 0.1623003, 
    0.1436855, 0.1490301, 0.1337081, 0.1412223, 0.1266612, 0.1206833, 
    0.115198, 0.1089543, 0.1674362, 0.1696798, 0.1656735, 0.1602059, 
    0.1552157, 0.1487012, 0.1480429, 0.1468404, 0.1437494, 0.1411758, 
    0.1464605, 0.1405344, 0.1634086, 0.1512081, 0.1705311, 0.1645918, 
    0.1605261, 0.1623043, 0.1531776, 0.1510643, 0.1426271, 0.1469588, 
    0.1221441, 0.1328334, 0.1043264, 0.1119283, 0.1704669, 0.1674443, 
    0.1571286, 0.1619969, 0.1482717, 0.1449855, 0.1423421, 0.1389975, 
    0.1386393, 0.1366794, 0.1398984, 0.1368061, 0.1486875, 0.1433164, 
    0.1582924, 0.1545788, 0.1562821, 0.1581604, 0.1523989, 0.1463763, 
    0.1462502, 0.1443454, 0.1390433, 0.1482173, 0.1207962, 0.1373909, 
    0.164178, 0.1584837, 0.15768, 0.1598684, 0.1453133, 0.1505072, 0.1367271, 
    0.1403858, 0.1344171, 0.1373665, 0.1378031, 0.1416453, 0.1440641, 
    0.1502668, 0.1554102, 0.1595502, 0.1585829, 0.1540518, 0.1460122, 
    0.1386064, 0.1402118, 0.1348661, 0.1492465, 0.1431264, 0.1454762, 
    0.1393899, 0.1528976, 0.1413517, 0.1559209, 0.1546153, 0.1506112, 
    0.1427152, 0.1409989, 0.1391758, 0.1402996, 0.1458111, 0.1467248, 
    0.1507082, 0.1518168, 0.1548992, 0.1574738, 0.1551204, 0.1526675, 
    0.1458093, 0.1397636, 0.1333204, 0.1317677, 0.1244784, 0.1303944, 
    0.1207067, 0.128916, 0.1148844, 0.1406983, 0.129164, 0.1504307, 
    0.1480613, 0.1438222, 0.1343369, 0.1394182, 0.1334858, 0.1467608, 
    0.1538959, 0.155771, 0.1592968, 0.1556909, 0.1559827, 0.1525672, 
    0.1536607, 0.1455843, 0.1498956, 0.1378138, 0.1335324, 0.1218174, 
    0.1149112, 0.1081007, 0.1051638, 0.1042786, 0.1039096,
  0.04576219, 0.04345123, 0.04389507, 0.04207106, 0.04307738, 0.04189106, 
    0.04528815, 0.04336079, 0.04458559, 0.04555149, 0.03866079, 0.04199079, 
    0.03537561, 0.03737251, 0.03248139, 0.03568183, 0.03185815, 0.03257148, 
    0.03045431, 0.03105198, 0.02843791, 0.03018086, 0.02713869, 0.02884851, 
    0.02857666, 0.03023941, 0.04130784, 0.03906637, 0.04144289, 0.04111811, 
    0.04126373, 0.04305632, 0.04397652, 0.04594196, 0.04558146, 0.04413984, 
    0.04097256, 0.04203235, 0.03939275, 0.03945125, 0.03662903, 0.03788599, 
    0.03332941, 0.03458877, 0.03102689, 0.03190048, 0.03106755, 0.03131873, 
    0.03106428, 0.03235152, 0.03179608, 0.03294326, 0.03764858, 0.03622625, 
    0.04056557, 0.04331584, 0.04520252, 0.04656971, 0.04637498, 0.04600501, 
    0.04413148, 0.04241187, 0.04112829, 0.04028265, 0.03945966, 0.03702914, 
    0.03578074, 0.03307805, 0.03355657, 0.03274858, 0.03198821, 0.03073571, 
    0.0309398, 0.0303954, 0.03276993, 0.03117956, 0.03383094, 0.03309263, 
    0.0392365, 0.04174492, 0.04283804, 0.0438095, 0.04622556, 0.04454889, 
    0.04520549, 0.0436529, 0.04268271, 0.04316099, 0.04025967, 0.04137339, 
    0.03570756, 0.03808696, 0.03207634, 0.03345803, 0.03175046, 0.03261504, 
    0.03114219, 0.03246588, 0.03019438, 0.02971298, 0.03004142, 0.02879219, 
    0.03254021, 0.03106745, 0.04317439, 0.04309614, 0.04273288, 0.04434321, 
    0.04444293, 0.0459518, 0.04460787, 0.04404256, 0.04262697, 0.04180222, 
    0.04102712, 0.03935309, 0.03753223, 0.03507256, 0.03336738, 0.03225308, 
    0.03293369, 0.03233235, 0.03300498, 0.0333232, 0.02989274, 0.03179087, 
    0.02896986, 0.02912179, 0.03038248, 0.02910465, 0.04304127, 0.04349228, 
    0.04507926, 0.04383447, 0.04611792, 0.04483123, 0.04410094, 0.04134968, 
    0.04075947, 0.04021632, 0.03915657, 0.03782103, 0.03554485, 0.03363344, 
    0.03194435, 0.03206633, 0.03202335, 0.03165257, 0.03257567, 0.03150259, 
    0.03132454, 0.03179122, 0.02914217, 0.02988459, 0.02912503, 0.02960696, 
    0.04334541, 0.04258968, 0.04299705, 0.04223284, 0.0427703, 0.04041082, 
    0.03971883, 0.03657536, 0.03784699, 0.03583574, 0.03763976, 0.03731615, 
    0.03577078, 0.03754099, 0.03373696, 0.0362888, 0.03163822, 0.03409006, 
    0.03148825, 0.03195154, 0.03118683, 0.03051143, 0.02967477, 0.02816812, 
    0.02851274, 0.02728063, 0.0414777, 0.04052416, 0.04060781, 0.03962293, 
    0.03890375, 0.03737214, 0.03499205, 0.03587608, 0.03426356, 0.03394516, 
    0.03639911, 0.03487998, 0.03989351, 0.03905591, 0.0395535, 0.04140187, 
    0.0356709, 0.03854822, 0.03333959, 0.03482061, 0.03060715, 0.03266104, 
    0.02870351, 0.02710633, 0.02565541, 0.0240216, 0.04000954, 0.04065112, 
    0.03950683, 0.03795524, 0.03654933, 0.03472912, 0.03454616, 0.03421239, 
    0.03335722, 0.03264825, 0.03410707, 0.032472, 0.03886273, 0.03542755, 
    0.04089506, 0.03919898, 0.03804576, 0.03854933, 0.03597801, 0.03538739, 
    0.03304772, 0.03424521, 0.02749512, 0.03036966, 0.02282303, 0.02479745, 
    0.04087666, 0.04001184, 0.0370871, 0.03846219, 0.03460971, 0.03369873, 
    0.03296918, 0.03205038, 0.03195227, 0.03141637, 0.03229741, 0.03145096, 
    0.0347253, 0.03323773, 0.03741496, 0.03637062, 0.03684893, 0.03737773, 
    0.03576018, 0.03408376, 0.03404879, 0.0335218, 0.032063, 0.0345946, 
    0.02713639, 0.03161079, 0.03908129, 0.03746894, 0.03724236, 0.03785981, 
    0.03378939, 0.035232, 0.03142941, 0.03243119, 0.03079989, 0.03160406, 
    0.03172342, 0.03277738, 0.03344409, 0.03516499, 0.03660395, 0.03776992, 
    0.03749688, 0.03622287, 0.03398287, 0.03194325, 0.03238343, 0.03092206, 
    0.03488083, 0.03318534, 0.03383448, 0.03215793, 0.03589967, 0.03269666, 
    0.03674742, 0.03638088, 0.03526101, 0.03307198, 0.03259962, 0.03209925, 
    0.03240752, 0.03392718, 0.03418034, 0.03528806, 0.0355975, 0.03646052, 
    0.03718428, 0.03652258, 0.03583529, 0.03392667, 0.03226042, 0.03050184, 
    0.03008075, 0.02811844, 0.02970926, 0.02711258, 0.02931027, 0.02557294, 
    0.03251706, 0.02937711, 0.03521067, 0.03455126, 0.03337733, 0.0307781, 
    0.0321657, 0.03054676, 0.0341903, 0.03617921, 0.0367053, 0.03769835, 
    0.03668278, 0.03676477, 0.03580723, 0.0361133, 0.03386438, 0.03506156, 
    0.03172634, 0.03055942, 0.02740807, 0.02557998, 0.0237997, 0.0230391, 
    0.0228107, 0.02271563,
  0.003994536, 0.003745579, 0.003793125, 0.003598556, 0.003705629, 
    0.003579474, 0.003943187, 0.003735907, 0.003867351, 0.003971694, 
    0.003240785, 0.003590044, 0.002903856, 0.003107728, 0.002613652, 
    0.002934932, 0.002552004, 0.002622586, 0.002414273, 0.002472716, 
    0.002219269, 0.002387631, 0.002095438, 0.002258702, 0.002232577, 
    0.00239333, 0.003517796, 0.003282915, 0.003532058, 0.003497782, 
    0.003513141, 0.003703383, 0.003801867, 0.004014044, 0.003974942, 
    0.003819402, 0.003482445, 0.003594449, 0.003316895, 0.003322994, 
    0.003031483, 0.003160617, 0.002698018, 0.002824329, 0.002470258, 
    0.002556179, 0.002474243, 0.002498893, 0.002473923, 0.002600779, 
    0.00254588, 0.002659531, 0.003136141, 0.002990345, 0.003439632, 
    0.003731105, 0.003933928, 0.004082331, 0.004061122, 0.004020892, 
    0.003818504, 0.003634742, 0.003498854, 0.003409936, 0.003323871, 
    0.003072469, 0.002944982, 0.002672953, 0.002720712, 0.002640172, 
    0.002564841, 0.002441754, 0.002461725, 0.002408529, 0.002642293, 
    0.00248523, 0.002748175, 0.002674405, 0.003300623, 0.003563996, 
    0.003680106, 0.003783949, 0.004044864, 0.0038634, 0.00393425, 
    0.003767165, 0.003663556, 0.003714556, 0.003407527, 0.003524717, 
    0.002937544, 0.00318137, 0.002573549, 0.002710863, 0.002541381, 
    0.002626908, 0.002481564, 0.002612111, 0.002388947, 0.002342188, 
    0.002374069, 0.002253283, 0.002619483, 0.002474234, 0.003715986, 
    0.003707632, 0.003668898, 0.003841263, 0.003851992, 0.004015113, 
    0.003869752, 0.003808954, 0.00365762, 0.003570063, 0.003488191, 
    0.003312762, 0.00312416, 0.002873172, 0.002701808, 0.00259103, 
    0.002658579, 0.002598879, 0.002665675, 0.002697397, 0.002359626, 
    0.002545366, 0.002270382, 0.002285026, 0.00240727, 0.002283373, 
    0.003701776, 0.00374997, 0.003920607, 0.003786625, 0.00403316, 
    0.003893831, 0.003815224, 0.003522214, 0.003460014, 0.003402984, 
    0.003292294, 0.003153916, 0.002921021, 0.002728401, 0.00256051, 
    0.00257256, 0.002568312, 0.002531735, 0.002623002, 0.002516969, 
    0.002499465, 0.0025454, 0.002286992, 0.002358834, 0.002285338, 
    0.002331915, 0.00373426, 0.003653653, 0.003697057, 0.003615723, 
    0.003672884, 0.003423385, 0.003350927, 0.003025996, 0.003156594, 
    0.002950574, 0.003135232, 0.003101935, 0.002943972, 0.00312506, 
    0.002738764, 0.002996728, 0.002530321, 0.002774168, 0.002515559, 
    0.00256122, 0.002485942, 0.002419847, 0.002338484, 0.002193434, 
    0.002226443, 0.002108895, 0.003535735, 0.003435283, 0.003444068, 
    0.003340909, 0.003266003, 0.003107689, 0.00286503, 0.002954675, 
    0.002791595, 0.002759626, 0.003007985, 0.002853708, 0.003369184, 
    0.003281823, 0.003333662, 0.003527725, 0.002933819, 0.003229109, 
    0.002699035, 0.002847712, 0.002429192, 0.002631477, 0.002244759, 
    0.002092374, 0.001955873, 0.001804454, 0.003381324, 0.00344862, 
    0.003328791, 0.003167766, 0.003023334, 0.00283848, 0.002820035, 
    0.002786453, 0.002700793, 0.002630205, 0.002775875, 0.002612717, 
    0.003261747, 0.002909121, 0.003474282, 0.003296711, 0.003177114, 
    0.003229221, 0.002965049, 0.002905047, 0.002669933, 0.00278975, 
    0.002129267, 0.002406022, 0.001694966, 0.001876052, 0.003472344, 
    0.003381565, 0.003078413, 0.003220191, 0.002826439, 0.002734935, 
    0.00266211, 0.002570984, 0.002561292, 0.00250849, 0.002595419, 
    0.002511891, 0.002838095, 0.00268887, 0.003112092, 0.003005077, 
    0.003053991, 0.003108264, 0.002942889, 0.002773534, 0.002770022, 
    0.002717237, 0.002572238, 0.002824916, 0.002095225, 0.002527626, 
    0.00328446, 0.003117648, 0.003094352, 0.003157916, 0.002744013, 
    0.002889305, 0.002509772, 0.002608672, 0.002448031, 0.002526956, 
    0.002538716, 0.002643033, 0.00270947, 0.002882523, 0.003028918, 
    0.003148645, 0.00312052, 0.00299, 0.002763408, 0.002560402, 0.002603941, 
    0.002459988, 0.002853793, 0.002683647, 0.002748531, 0.002581617, 
    0.002957076, 0.002635019, 0.003043596, 0.003006123, 0.002892243, 
    0.00267235, 0.002625378, 0.002575815, 0.002606326, 0.002757824, 
    0.002783232, 0.002894982, 0.002926364, 0.003014256, 0.003088386, 
    0.003020599, 0.002950527, 0.002757771, 0.002591758, 0.002418911, 
    0.002377893, 0.002188687, 0.002341829, 0.002092971, 0.002303225, 
    0.001948174, 0.00261719, 0.00230968, 0.002887144, 0.002820548, 
    0.002702804, 0.002445902, 0.002582385, 0.002423297, 0.002784233, 
    0.00298555, 0.003039285, 0.003141268, 0.003036981, 0.003045373, 
    0.002947673, 0.002978829, 0.002751527, 0.002872057, 0.002539004, 
    0.002424533, 0.002120994, 0.00194883, 0.001784079, 0.001714601, 
    0.001693847, 0.001685222,
  0.0001100816, 0.0001015489, 0.0001031674, 9.657819e-05, 0.0001001931, 
    9.593687e-05, 0.00010831, 0.0001012204, 0.0001057046, 0.0001092927, 
    8.470473e-05, 9.629199e-05, 7.382834e-05, 8.037269e-05, 6.471662e-05, 
    7.481847e-05, 6.281333e-05, 6.499336e-05, 5.86039e-05, 6.038274e-05, 
    5.274922e-05, 5.779663e-05, 4.909829e-05, 5.392287e-05, 5.314471e-05, 
    5.796912e-05, 9.386994e-05, 8.608603e-05, 9.434706e-05, 9.32013e-05, 
    9.371434e-05, 0.000100117, 0.0001034656, 0.0001107561, 0.0001094048, 
    0.0001040642, 9.268957e-05, 9.644002e-05, 8.720325e-05, 8.740414e-05, 
    7.791179e-05, 8.208893e-05, 6.73399e-05, 7.130691e-05, 6.030769e-05, 
    6.294182e-05, 6.042936e-05, 6.118302e-05, 6.041959e-05, 6.431818e-05, 
    6.262486e-05, 6.614051e-05, 8.129374e-05, 7.659065e-05, 9.126414e-05, 
    0.0001010574, 0.0001079912, 0.0001131243, 0.0001123876, 0.0001109932, 
    0.0001040335, 9.779676e-05, 9.323705e-05, 9.02781e-05, 8.743304e-05, 
    7.923283e-05, 7.513925e-05, 6.655831e-05, 6.804917e-05, 6.553891e-05, 
    6.320866e-05, 5.9439e-05, 6.004737e-05, 5.842968e-05, 6.560474e-05, 
    6.076508e-05, 6.890956e-05, 6.660348e-05, 8.666801e-05, 9.541727e-05, 
    9.932904e-05, 0.0001028546, 0.0001118236, 0.0001055692, 0.0001080023, 
    0.000102283, 9.876936e-05, 0.0001004957, 9.019821e-05, 9.410139e-05, 
    7.490179e-05, 8.276444e-05, 6.347713e-05, 6.774117e-05, 6.248649e-05, 
    6.512734e-05, 6.065301e-05, 6.466882e-05, 5.783646e-05, 5.642502e-05, 
    5.738659e-05, 5.376125e-05, 6.489718e-05, 6.042912e-05, 0.0001005442, 
    0.000100261, 9.894988e-05, 0.0001048114, 0.0001051786, 0.0001107931, 
    0.0001057869, 0.0001037074, 9.856883e-05, 9.562086e-05, 9.288118e-05, 
    8.706722e-05, 8.090514e-05, 7.285335e-05, 6.745826e-05, 6.40168e-05, 
    6.611085e-05, 6.42594e-05, 6.633166e-05, 6.73205e-05, 5.695057e-05, 
    6.260907e-05, 5.427152e-05, 5.470928e-05, 5.839152e-05, 5.465982e-05, 
    0.0001000625, 0.0001016981, 0.0001075329, 0.0001029458, 0.000111418, 
    0.0001066128, 0.0001039215, 9.401773e-05, 9.194211e-05, 9.00476e-05, 
    8.639396e-05, 8.187106e-05, 7.437485e-05, 6.828988e-05, 6.307519e-05, 
    6.344661e-05, 6.331563e-05, 6.219009e-05, 6.500624e-05, 6.173688e-05, 
    6.120053e-05, 6.261009e-05, 5.47681e-05, 5.692664e-05, 5.471861e-05, 
    5.611584e-05, 0.0001011644, 9.843487e-05, 9.99027e-05, 9.715588e-05, 
    9.908468e-05, 9.072444e-05, 8.83255e-05, 7.773538e-05, 8.195813e-05, 
    7.531782e-05, 8.126424e-05, 8.018516e-05, 7.510704e-05, 8.093425e-05, 
    6.861454e-05, 7.679538e-05, 6.214666e-05, 6.972605e-05, 6.169364e-05, 
    6.309706e-05, 6.078681e-05, 5.877309e-05, 5.631349e-05, 5.198309e-05, 
    5.29623e-05, 4.949241e-05, 9.447013e-05, 9.111959e-05, 9.141158e-05, 
    8.799478e-05, 8.55308e-05, 8.037141e-05, 7.25951e-05, 7.544882e-05, 
    7.027436e-05, 6.926896e-05, 7.715655e-05, 7.22363e-05, 8.892867e-05, 
    8.605004e-05, 8.775578e-05, 9.420207e-05, 7.478293e-05, 8.432258e-05, 
    6.737164e-05, 7.204641e-05, 5.905697e-05, 6.526907e-05, 5.350726e-05, 
    4.900867e-05, 4.504903e-05, 4.073846e-05, 8.93302e-05, 9.156296e-05, 
    8.759519e-05, 8.232155e-05, 7.76497e-05, 7.175426e-05, 7.117127e-05, 
    7.011246e-05, 6.742654e-05, 6.522958e-05, 6.977966e-05, 6.468761e-05, 
    8.539138e-05, 7.399586e-05, 9.241742e-05, 8.653924e-05, 8.262581e-05, 
    8.432622e-05, 7.57805e-05, 7.386618e-05, 6.646424e-05, 7.021627e-05, 
    5.009037e-05, 5.83537e-05, 3.767778e-05, 4.276571e-05, 9.235281e-05, 
    8.933814e-05, 7.942466e-05, 8.403102e-05, 7.137356e-05, 6.84945e-05, 
    6.622072e-05, 6.339804e-05, 6.309929e-05, 6.147695e-05, 6.415243e-05, 
    6.158118e-05, 7.174208e-05, 6.705439e-05, 8.051397e-05, 7.70632e-05, 
    7.863659e-05, 8.039001e-05, 7.507232e-05, 6.970605e-05, 6.95956e-05, 
    6.794049e-05, 6.343688e-05, 7.132546e-05, 4.909219e-05, 6.206404e-05, 
    8.613657e-05, 8.069407e-05, 7.993982e-05, 8.200108e-05, 6.877903e-05, 
    7.336561e-05, 6.151622e-05, 6.456238e-05, 5.963006e-05, 6.204334e-05, 
    6.240459e-05, 6.562772e-05, 6.769763e-05, 7.315016e-05, 7.782929e-05, 
    8.169977e-05, 8.078707e-05, 7.657956e-05, 6.938781e-05, 6.307191e-05, 
    6.441599e-05, 5.999441e-05, 7.223893e-05, 6.689153e-05, 6.892077e-05, 
    6.372607e-05, 7.552559e-05, 6.537908e-05, 7.830167e-05, 7.709675e-05, 
    7.345897e-05, 6.653956e-05, 6.507989e-05, 6.354705e-05, 6.448977e-05, 
    6.92124e-05, 7.001109e-05, 7.354603e-05, 7.454516e-05, 7.735795e-05, 
    7.974687e-05, 7.756178e-05, 7.531633e-05, 6.921073e-05, 6.403931e-05, 
    5.874468e-05, 5.750212e-05, 5.184264e-05, 5.641427e-05, 4.902622e-05, 
    5.525453e-05, 4.482786e-05, 6.482624e-05, 5.544804e-05, 7.329693e-05, 
    7.11875e-05, 6.748938e-05, 5.956531e-05, 6.374978e-05, 5.88779e-05, 
    7.00426e-05, 7.643696e-05, 7.816288e-05, 8.146017e-05, 7.808871e-05, 
    7.835891e-05, 7.522509e-05, 7.622157e-05, 6.901474e-05, 7.281793e-05, 
    6.241346e-05, 5.891542e-05, 4.984734e-05, 4.484662e-05, 4.016519e-05, 
    3.822307e-05, 3.764673e-05, 3.740777e-05,
  8.462572e-07, 7.610096e-07, 7.770259e-07, 7.122837e-07, 7.476488e-07, 
    7.06049e-07, 8.283956e-07, 7.577677e-07, 8.022802e-07, 8.382931e-07, 
    5.988798e-07, 7.094998e-07, 4.990146e-07, 5.586182e-07, 4.186445e-07, 
    5.079355e-07, 4.022677e-07, 4.210375e-07, 3.665845e-07, 3.815715e-07, 
    3.182546e-07, 3.598286e-07, 2.889328e-07, 3.278165e-07, 3.214694e-07, 
    3.612698e-07, 6.860377e-07, 6.118466e-07, 6.906457e-07, 6.795918e-07, 
    6.845364e-07, 7.469009e-07, 7.799859e-07, 8.530792e-07, 8.394236e-07, 
    7.859322e-07, 6.746675e-07, 7.10939e-07, 6.223773e-07, 6.242753e-07, 
    5.360293e-07, 5.744934e-07, 4.414551e-07, 4.764585e-07, 3.809365e-07, 
    4.033682e-07, 3.819662e-07, 3.883582e-07, 3.818835e-07, 4.152035e-07, 
    4.006538e-07, 4.309916e-07, 5.671257e-07, 5.239891e-07, 6.609923e-07, 
    7.561608e-07, 8.251904e-07, 8.771259e-07, 8.696305e-07, 8.554802e-07, 
    7.856272e-07, 7.241626e-07, 6.799356e-07, 6.515687e-07, 6.245485e-07, 
    5.481304e-07, 5.108328e-07, 4.346304e-07, 4.476689e-07, 4.257651e-07, 
    4.056566e-07, 3.736034e-07, 3.787356e-07, 3.651242e-07, 4.263361e-07, 
    3.848107e-07, 4.55233e-07, 4.350239e-07, 6.173283e-07, 7.010062e-07, 
    7.391623e-07, 7.739253e-07, 8.639013e-07, 8.009288e-07, 8.253019e-07, 
    7.68265e-07, 7.336751e-07, 7.50626e-07, 6.508064e-07, 6.882721e-07, 
    5.086874e-07, 5.807693e-07, 4.079621e-07, 4.449681e-07, 3.994699e-07, 
    4.221972e-07, 3.838606e-07, 4.182309e-07, 3.601613e-07, 3.484163e-07, 
    3.564082e-07, 3.264956e-07, 4.202053e-07, 3.819642e-07, 7.511038e-07, 
    7.483166e-07, 7.354435e-07, 7.933703e-07, 7.970301e-07, 8.534541e-07, 
    8.031022e-07, 7.823863e-07, 7.317114e-07, 7.02981e-07, 6.765101e-07, 
    6.210929e-07, 5.63533e-07, 4.902648e-07, 4.424905e-07, 4.126052e-07, 
    4.307335e-07, 4.146964e-07, 4.326554e-07, 4.412851e-07, 3.527792e-07, 
    4.005187e-07, 3.306694e-07, 3.342596e-07, 3.648046e-07, 3.338536e-07, 
    7.463649e-07, 7.624827e-07, 8.205869e-07, 7.748284e-07, 8.597855e-07, 
    8.113634e-07, 7.845139e-07, 6.874646e-07, 6.674885e-07, 6.493703e-07, 
    6.147438e-07, 5.724726e-07, 5.039337e-07, 4.497824e-07, 4.045115e-07, 
    4.076997e-07, 4.065748e-07, 3.96937e-07, 4.211489e-07, 3.930711e-07, 
    3.885072e-07, 4.005273e-07, 3.347427e-07, 3.525801e-07, 3.343363e-07, 
    3.458551e-07, 7.572144e-07, 7.304005e-07, 7.447938e-07, 7.179097e-07, 
    7.367651e-07, 6.558311e-07, 6.329979e-07, 5.344185e-07, 5.732801e-07, 
    5.124472e-07, 5.668526e-07, 5.568896e-07, 5.105422e-07, 5.638016e-07, 
    4.526368e-07, 5.258515e-07, 3.965662e-07, 4.624385e-07, 3.927027e-07, 
    4.046991e-07, 3.849948e-07, 3.680042e-07, 3.474917e-07, 3.120475e-07, 
    3.199853e-07, 2.920663e-07, 6.918352e-07, 6.59609e-07, 6.624035e-07, 
    6.298633e-07, 6.066253e-07, 5.586062e-07, 4.879528e-07, 5.136321e-07, 
    4.6729e-07, 4.584013e-07, 5.291386e-07, 4.847454e-07, 6.387215e-07, 
    6.115069e-07, 6.27601e-07, 6.892448e-07, 5.076142e-07, 5.953023e-07, 
    4.417327e-07, 4.830495e-07, 3.703888e-07, 4.234255e-07, 3.244228e-07, 
    2.882217e-07, 2.572e-07, 2.243959e-07, 6.425383e-07, 6.638537e-07, 
    6.260815e-07, 5.766532e-07, 5.336358e-07, 4.804432e-07, 4.752518e-07, 
    4.658561e-07, 4.422128e-07, 4.230829e-07, 4.629119e-07, 4.183932e-07, 
    6.053177e-07, 5.00521e-07, 6.720515e-07, 6.161134e-07, 5.794802e-07, 
    5.953358e-07, 5.166357e-07, 4.993541e-07, 4.338104e-07, 4.667753e-07, 
    2.96836e-07, 3.644881e-07, 2.017592e-07, 2.396935e-07, 6.714307e-07, 
    6.426136e-07, 5.498916e-07, 5.925763e-07, 4.770517e-07, 4.515806e-07, 
    4.316895e-07, 4.072827e-07, 4.047183e-07, 3.908578e-07, 4.137741e-07, 
    3.917448e-07, 4.803347e-07, 4.38959e-07, 5.59921e-07, 5.282885e-07, 
    5.426604e-07, 5.587776e-07, 5.102273e-07, 4.622613e-07, 4.612848e-07, 
    4.467157e-07, 4.076179e-07, 4.766236e-07, 2.888854e-07, 3.958623e-07, 
    6.123203e-07, 5.615838e-07, 5.546297e-07, 5.736783e-07, 4.540838e-07, 
    4.948573e-07, 3.911919e-07, 4.173114e-07, 3.752133e-07, 3.956842e-07, 
    3.987697e-07, 4.265355e-07, 4.445866e-07, 4.929245e-07, 5.352756e-07, 
    5.708848e-07, 5.624418e-07, 5.238882e-07, 4.594503e-07, 4.044836e-07, 
    4.160478e-07, 3.782881e-07, 4.847686e-07, 4.37537e-07, 4.553322e-07, 
    4.101025e-07, 5.143271e-07, 4.243801e-07, 5.395939e-07, 5.285939e-07, 
    4.956952e-07, 4.344671e-07, 4.217865e-07, 4.085631e-07, 4.166843e-07, 
    4.579026e-07, 4.649588e-07, 4.964769e-07, 5.054688e-07, 5.309741e-07, 
    5.528537e-07, 5.328334e-07, 5.124336e-07, 4.578877e-07, 4.127994e-07, 
    3.677658e-07, 3.573711e-07, 3.109133e-07, 3.483277e-07, 2.883617e-07, 
    3.387455e-07, 2.554926e-07, 4.195925e-07, 3.403394e-07, 4.942407e-07, 
    4.753961e-07, 4.427633e-07, 3.746682e-07, 4.103065e-07, 3.688845e-07, 
    4.652376e-07, 5.225926e-07, 5.383242e-07, 5.686658e-07, 5.37646e-07, 
    5.401177e-07, 5.116081e-07, 5.20636e-07, 4.561598e-07, 4.899472e-07, 
    3.988456e-07, 3.691996e-07, 2.94895e-07, 2.556369e-07, 2.201129e-07, 
    2.057503e-07, 2.015324e-07, 1.997897e-07,
  1.022341e-09, 8.438348e-10, 8.765592e-10, 7.467173e-10, 8.168341e-10, 
    7.345637e-10, 9.840733e-10, 8.372589e-10, 9.289362e-10, 1.005222e-09, 
    5.360756e-10, 7.412825e-10, 3.708298e-10, 4.669836e-10, 2.540601e-10, 
    3.847323e-10, 2.322727e-10, 2.573026e-10, 1.873837e-10, 2.057934e-10, 
    1.326946e-10, 1.793018e-10, 1.032762e-10, 1.429222e-10, 1.360992e-10, 
    1.810144e-10, 6.959859e-10, 5.58994e-10, 7.048101e-10, 6.83703e-10, 
    6.931188e-10, 8.153314e-10, 8.826515e-10, 1.037072e-09, 1.007647e-09, 
    8.949239e-10, 6.743667e-10, 7.440893e-10, 5.778331e-10, 5.812513e-10, 
    4.296515e-10, 4.938429e-10, 2.855819e-10, 3.364856e-10, 2.05e-10, 
    2.337133e-10, 2.062871e-10, 2.143434e-10, 2.061836e-10, 2.494217e-10, 
    2.301644e-10, 2.709553e-10, 4.813147e-10, 4.101911e-10, 6.486557e-10, 
    8.340071e-10, 9.772543e-10, 1.089507e-09, 1.073079e-09, 1.042273e-09, 
    8.942931e-10, 7.700463e-10, 6.843552e-10, 6.311267e-10, 5.817438e-10, 
    4.495218e-10, 3.89285e-10, 2.760109e-10, 2.943989e-10, 2.637552e-10, 
    2.36721e-10, 1.95924e-10, 2.022597e-10, 1.856254e-10, 2.645377e-10, 
    2.098584e-10, 3.052613e-10, 2.765587e-10, 5.687779e-10, 7.247787e-10, 
    7.998308e-10, 8.701941e-10, 1.060574e-09, 9.261105e-10, 9.774916e-10, 
    8.586098e-10, 7.888917e-10, 8.228263e-10, 6.297158e-10, 7.0026e-10, 
    3.859117e-10, 5.046004e-10, 2.397656e-10, 2.905547e-10, 2.286227e-10, 
    2.588796e-10, 2.086629e-10, 2.534997e-10, 1.796967e-10, 1.659646e-10, 
    1.752629e-10, 1.414908e-10, 2.561727e-10, 2.062849e-10, 8.237894e-10, 
    8.181769e-10, 7.924107e-10, 9.103509e-10, 9.179708e-10, 1.037883e-09, 
    9.306566e-10, 8.875981e-10, 7.849892e-10, 7.286052e-10, 6.778544e-10, 
    5.755243e-10, 4.752456e-10, 3.573684e-10, 2.870444e-10, 2.459405e-10, 
    2.705978e-10, 2.487405e-10, 2.732621e-10, 2.853416e-10, 1.710165e-10, 
    2.299885e-10, 1.460317e-10, 1.49983e-10, 1.852415e-10, 1.49534e-10, 
    8.142539e-10, 8.468271e-10, 9.674851e-10, 8.720457e-10, 1.051616e-09, 
    9.480031e-10, 8.919922e-10, 6.987157e-10, 6.608281e-10, 6.270607e-10, 
    5.641531e-10, 4.903959e-10, 3.784728e-10, 2.974203e-10, 2.35214e-10, 
    2.394181e-10, 2.379317e-10, 2.253375e-10, 2.574538e-10, 2.203577e-10, 
    2.145331e-10, 2.299993e-10, 1.505178e-10, 1.707842e-10, 1.500678e-10, 
    1.630261e-10, 8.36136e-10, 7.82388e-10, 8.111e-10, 7.577376e-10, 
    7.950448e-10, 6.390375e-10, 5.970469e-10, 4.270312e-10, 4.917726e-10, 
    3.918295e-10, 4.80852e-10, 4.640896e-10, 3.888286e-10, 4.75697e-10, 
    3.015184e-10, 4.131823e-10, 2.24858e-10, 3.157418e-10, 2.198854e-10, 
    2.354606e-10, 2.100896e-10, 1.890995e-10, 1.649013e-10, 1.26218e-10, 
    1.345226e-10, 1.06275e-10, 7.070934e-10, 6.460734e-10, 6.512931e-10, 
    5.913536e-10, 5.497232e-10, 4.669629e-10, 3.538403e-10, 3.937001e-10, 
    3.228654e-10, 3.098534e-10, 4.184755e-10, 3.489672e-10, 6.074842e-10, 
    5.583866e-10, 5.872573e-10, 7.021241e-10, 3.842278e-10, 5.298056e-10, 
    2.859738e-10, 3.463994e-10, 1.919947e-10, 2.60555e-10, 1.392572e-10, 
    1.026011e-10, 7.496886e-11, 4.992519e-11, 6.144772e-10, 6.540076e-10, 
    5.845104e-10, 4.975372e-10, 4.257583e-10, 3.424674e-10, 3.346816e-10, 
    3.207537e-10, 2.866516e-10, 2.600866e-10, 3.164334e-10, 2.53719e-10, 
    5.474141e-10, 3.731641e-10, 6.694229e-10, 5.666017e-10, 5.023845e-10, 
    5.29863e-10, 3.98458e-10, 3.713541e-10, 2.748686e-10, 3.221068e-10, 
    1.109088e-10, 1.848622e-10, 3.536804e-11, 6.104427e-11, 6.682508e-10, 
    6.14615e-10, 4.524367e-10, 5.250456e-10, 3.373738e-10, 2.999989e-10, 
    2.719219e-10, 2.388672e-10, 2.354859e-10, 2.175257e-10, 2.475041e-10, 
    2.186589e-10, 3.42304e-10, 2.820673e-10, 4.691679e-10, 4.171044e-10, 
    4.404999e-10, 4.6725e-10, 3.883301e-10, 3.154816e-10, 3.140535e-10, 
    2.930406e-10, 2.393136e-10, 3.367327e-10, 1.032329e-10, 2.239519e-10, 
    5.598323e-10, 4.719639e-10, 4.60315e-10, 4.92451e-10, 3.036023e-10, 
    3.644112e-10, 2.179523e-10, 2.522584e-10, 1.979031e-10, 2.237192e-10, 
    2.277127e-10, 2.648113e-10, 2.900132e-10, 3.614413e-10, 4.284243e-10, 
    4.876926e-10, 4.734057e-10, 4.100292e-10, 3.113799e-10, 2.351778e-10, 
    2.505569e-10, 2.017042e-10, 3.490016e-10, 2.800726e-10, 3.054056e-10, 
    2.426049e-10, 3.947996e-10, 2.618614e-10, 4.354714e-10, 4.175965e-10, 
    3.657016e-10, 2.757837e-10, 2.583206e-10, 2.405619e-10, 2.514131e-10, 
    3.091296e-10, 3.194348e-10, 3.669064e-10, 3.808689e-10, 4.214424e-10, 
    4.573558e-10, 4.244554e-10, 3.918077e-10, 3.091074e-10, 2.462006e-10, 
    1.888112e-10, 1.763961e-10, 1.2505e-10, 1.658636e-10, 1.027354e-10, 
    1.549814e-10, 7.355739e-11, 2.553439e-10, 1.567702e-10, 3.634625e-10, 
    3.348971e-10, 2.874311e-10, 1.972331e-10, 2.428762e-10, 1.901671e-10, 
    3.198443e-10, 4.079545e-10, 4.333952e-10, 4.839241e-10, 4.322875e-10, 
    4.36329e-10, 3.905047e-10, 4.048257e-10, 3.066024e-10, 3.568821e-10, 
    2.278116e-10, 1.905492e-10, 1.09013e-10, 7.367554e-11, 4.699335e-11, 
    3.77644e-11, 3.523394e-11, 3.421278e-11,
  4.04842e-13, 4.041397e-13, 4.042685e-13, 4.037571e-13, 4.040333e-13, 
    4.037092e-13, 4.046915e-13, 4.041138e-13, 4.044746e-13, 4.047747e-13, 
    4.029258e-13, 4.037356e-13, 4.02272e-13, 4.026527e-13, 4.01809e-13, 
    4.023271e-13, 4.017224e-13, 4.018219e-13, 4.01544e-13, 4.016172e-13, 
    4.013263e-13, 4.015119e-13, 4.01209e-13, 4.013671e-13, 4.013399e-13, 
    4.015187e-13, 4.03557e-13, 4.030164e-13, 4.035918e-13, 4.035086e-13, 
    4.035457e-13, 4.040274e-13, 4.042925e-13, 4.048999e-13, 4.047842e-13, 
    4.043408e-13, 4.034718e-13, 4.037467e-13, 4.030908e-13, 4.031043e-13, 
    4.025049e-13, 4.027589e-13, 4.019341e-13, 4.021359e-13, 4.016141e-13, 
    4.017282e-13, 4.016192e-13, 4.016512e-13, 4.016188e-13, 4.017906e-13, 
    4.017141e-13, 4.01876e-13, 4.027093e-13, 4.024279e-13, 4.033703e-13, 
    4.04101e-13, 4.046647e-13, 4.05106e-13, 4.050414e-13, 4.049203e-13, 
    4.043383e-13, 4.03849e-13, 4.035112e-13, 4.033012e-13, 4.031062e-13, 
    4.025836e-13, 4.023451e-13, 4.018961e-13, 4.019691e-13, 4.018475e-13, 
    4.017401e-13, 4.01578e-13, 4.016032e-13, 4.01537e-13, 4.018506e-13, 
    4.016334e-13, 4.020121e-13, 4.018983e-13, 4.03055e-13, 4.036706e-13, 
    4.039664e-13, 4.042435e-13, 4.049923e-13, 4.044635e-13, 4.046656e-13, 
    4.041978e-13, 4.039233e-13, 4.040569e-13, 4.032956e-13, 4.035739e-13, 
    4.023318e-13, 4.028014e-13, 4.017522e-13, 4.019538e-13, 4.017079e-13, 
    4.018281e-13, 4.016286e-13, 4.018068e-13, 4.015134e-13, 4.014588e-13, 
    4.014958e-13, 4.013614e-13, 4.018174e-13, 4.016192e-13, 4.040607e-13, 
    4.040386e-13, 4.039371e-13, 4.044015e-13, 4.044315e-13, 4.049031e-13, 
    4.044814e-13, 4.043119e-13, 4.039079e-13, 4.036857e-13, 4.034855e-13, 
    4.030816e-13, 4.026853e-13, 4.022187e-13, 4.019399e-13, 4.017767e-13, 
    4.018746e-13, 4.017878e-13, 4.018852e-13, 4.019331e-13, 4.014789e-13, 
    4.017134e-13, 4.013795e-13, 4.013952e-13, 4.015355e-13, 4.013934e-13, 
    4.040232e-13, 4.041515e-13, 4.046263e-13, 4.042507e-13, 4.04957e-13, 
    4.045496e-13, 4.043292e-13, 4.035678e-13, 4.034184e-13, 4.032851e-13, 
    4.030367e-13, 4.027452e-13, 4.023023e-13, 4.01981e-13, 4.017341e-13, 
    4.017508e-13, 4.017449e-13, 4.016949e-13, 4.018225e-13, 4.016751e-13, 
    4.01652e-13, 4.017134e-13, 4.013973e-13, 4.01478e-13, 4.013955e-13, 
    4.014471e-13, 4.041093e-13, 4.038976e-13, 4.040108e-13, 4.038005e-13, 
    4.039475e-13, 4.033324e-13, 4.031666e-13, 4.024946e-13, 4.027507e-13, 
    4.023552e-13, 4.027075e-13, 4.026412e-13, 4.023433e-13, 4.026871e-13, 
    4.019973e-13, 4.024397e-13, 4.01693e-13, 4.020537e-13, 4.016732e-13, 
    4.017351e-13, 4.016343e-13, 4.015508e-13, 4.014546e-13, 4.013005e-13, 
    4.013336e-13, 4.01221e-13, 4.036008e-13, 4.033602e-13, 4.033808e-13, 
    4.031442e-13, 4.029797e-13, 4.026526e-13, 4.022047e-13, 4.023626e-13, 
    4.02082e-13, 4.020304e-13, 4.024607e-13, 4.021854e-13, 4.032078e-13, 
    4.030139e-13, 4.03128e-13, 4.035812e-13, 4.023251e-13, 4.02901e-13, 
    4.019356e-13, 4.021752e-13, 4.015624e-13, 4.018348e-13, 4.013525e-13, 
    4.012064e-13, 4.010961e-13, 4.00996e-13, 4.032354e-13, 4.033915e-13, 
    4.031171e-13, 4.027735e-13, 4.024895e-13, 4.021596e-13, 4.021288e-13, 
    4.020736e-13, 4.019383e-13, 4.018329e-13, 4.020565e-13, 4.018076e-13, 
    4.029706e-13, 4.022813e-13, 4.034523e-13, 4.030464e-13, 4.027926e-13, 
    4.029012e-13, 4.023814e-13, 4.022741e-13, 4.018916e-13, 4.02079e-13, 
    4.012395e-13, 4.01534e-13, 4.009378e-13, 4.010405e-13, 4.034476e-13, 
    4.03236e-13, 4.025951e-13, 4.028822e-13, 4.021394e-13, 4.019913e-13, 
    4.018799e-13, 4.017486e-13, 4.017352e-13, 4.016639e-13, 4.017829e-13, 
    4.016684e-13, 4.02159e-13, 4.019201e-13, 4.026613e-13, 4.024553e-13, 
    4.025479e-13, 4.026537e-13, 4.023414e-13, 4.020527e-13, 4.02047e-13, 
    4.019637e-13, 4.017504e-13, 4.021369e-13, 4.012089e-13, 4.016894e-13, 
    4.030197e-13, 4.026723e-13, 4.026263e-13, 4.027534e-13, 4.020056e-13, 
    4.022466e-13, 4.016655e-13, 4.018018e-13, 4.015859e-13, 4.016885e-13, 
    4.017043e-13, 4.018516e-13, 4.019517e-13, 4.022348e-13, 4.025001e-13, 
    4.027345e-13, 4.026781e-13, 4.024273e-13, 4.020364e-13, 4.01734e-13, 
    4.017951e-13, 4.01601e-13, 4.021855e-13, 4.019122e-13, 4.020127e-13, 
    4.017635e-13, 4.02367e-13, 4.018399e-13, 4.02528e-13, 4.024572e-13, 
    4.022517e-13, 4.018952e-13, 4.018259e-13, 4.017554e-13, 4.017985e-13, 
    4.020275e-13, 4.020684e-13, 4.022565e-13, 4.023118e-13, 4.024725e-13, 
    4.026146e-13, 4.024844e-13, 4.023551e-13, 4.020274e-13, 4.017778e-13, 
    4.015497e-13, 4.015003e-13, 4.012959e-13, 4.014584e-13, 4.012069e-13, 
    4.014151e-13, 4.010905e-13, 4.018141e-13, 4.014222e-13, 4.022428e-13, 
    4.021296e-13, 4.019414e-13, 4.015832e-13, 4.017646e-13, 4.015551e-13, 
    4.0207e-13, 4.024191e-13, 4.025198e-13, 4.027197e-13, 4.025154e-13, 
    4.025314e-13, 4.023499e-13, 4.024067e-13, 4.020175e-13, 4.022168e-13, 
    4.017047e-13, 4.015566e-13, 4.012319e-13, 4.010909e-13, 4.009843e-13, 
    4.009474e-13, 4.009373e-13, 4.009332e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949657e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 
    8.949655e-07, 8.949656e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949656e-07, 
    8.949656e-07, 8.949657e-07, 8.949657e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949653e-07, 8.949652e-07, 8.949654e-07, 8.949653e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949657e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949656e-07, 8.949656e-07, 8.949657e-07, 8.949656e-07, 8.949657e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.94965e-07, 8.949651e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.94965e-07, 8.94965e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.760409e-16, 6.778689e-16, 6.775138e-16, 6.789867e-16, 6.7817e-16, 
    6.791341e-16, 6.764119e-16, 6.779412e-16, 6.769652e-16, 6.762059e-16, 
    6.818409e-16, 6.790525e-16, 6.847346e-16, 6.829595e-16, 6.874156e-16, 
    6.844582e-16, 6.880114e-16, 6.873309e-16, 6.893794e-16, 6.887928e-16, 
    6.914089e-16, 6.8965e-16, 6.927641e-16, 6.909893e-16, 6.912668e-16, 
    6.895919e-16, 6.796146e-16, 6.814938e-16, 6.79503e-16, 6.797712e-16, 
    6.79651e-16, 6.781867e-16, 6.77448e-16, 6.759015e-16, 6.761824e-16, 
    6.773185e-16, 6.798917e-16, 6.79019e-16, 6.812187e-16, 6.81169e-16, 
    6.836142e-16, 6.825121e-16, 6.866168e-16, 6.854514e-16, 6.888173e-16, 
    6.879714e-16, 6.887775e-16, 6.885332e-16, 6.887807e-16, 6.875399e-16, 
    6.880716e-16, 6.869796e-16, 6.827185e-16, 6.839718e-16, 6.802308e-16, 
    6.779766e-16, 6.764789e-16, 6.75415e-16, 6.755654e-16, 6.758521e-16, 
    6.773251e-16, 6.787093e-16, 6.797633e-16, 6.804679e-16, 6.811619e-16, 
    6.832594e-16, 6.843697e-16, 6.868521e-16, 6.864049e-16, 6.871628e-16, 
    6.878873e-16, 6.891021e-16, 6.889023e-16, 6.894372e-16, 6.871432e-16, 
    6.88668e-16, 6.861499e-16, 6.86839e-16, 6.813487e-16, 6.792546e-16, 
    6.783622e-16, 6.77582e-16, 6.75681e-16, 6.769939e-16, 6.764765e-16, 
    6.777077e-16, 6.784893e-16, 6.781028e-16, 6.804872e-16, 6.795605e-16, 
    6.844355e-16, 6.823374e-16, 6.878028e-16, 6.864968e-16, 6.881157e-16, 
    6.872899e-16, 6.887045e-16, 6.874315e-16, 6.896364e-16, 6.901159e-16, 
    6.897882e-16, 6.910472e-16, 6.873608e-16, 6.887773e-16, 6.780919e-16, 
    6.781549e-16, 6.784487e-16, 6.771569e-16, 6.770779e-16, 6.758937e-16, 
    6.769476e-16, 6.773961e-16, 6.785347e-16, 6.792075e-16, 6.79847e-16, 
    6.812521e-16, 6.828196e-16, 6.850096e-16, 6.865814e-16, 6.876341e-16, 
    6.869888e-16, 6.875585e-16, 6.869215e-16, 6.86623e-16, 6.899361e-16, 
    6.880765e-16, 6.908662e-16, 6.907121e-16, 6.894499e-16, 6.907294e-16, 
    6.781992e-16, 6.778365e-16, 6.765758e-16, 6.775625e-16, 6.757647e-16, 
    6.76771e-16, 6.773492e-16, 6.795795e-16, 6.800695e-16, 6.805233e-16, 
    6.814194e-16, 6.825686e-16, 6.845824e-16, 6.863329e-16, 6.879295e-16, 
    6.878126e-16, 6.878537e-16, 6.8821e-16, 6.873271e-16, 6.883549e-16, 
    6.885272e-16, 6.880765e-16, 6.906914e-16, 6.899448e-16, 6.907088e-16, 
    6.902227e-16, 6.779544e-16, 6.785648e-16, 6.78235e-16, 6.78855e-16, 
    6.784181e-16, 6.803597e-16, 6.809414e-16, 6.83661e-16, 6.825459e-16, 
    6.843208e-16, 6.827264e-16, 6.830089e-16, 6.843779e-16, 6.828127e-16, 
    6.862361e-16, 6.839153e-16, 6.882239e-16, 6.859084e-16, 6.883688e-16, 
    6.879226e-16, 6.886615e-16, 6.893228e-16, 6.901546e-16, 6.916878e-16, 
    6.91333e-16, 6.926146e-16, 6.794745e-16, 6.802653e-16, 6.80196e-16, 
    6.810234e-16, 6.81635e-16, 6.829602e-16, 6.850831e-16, 6.842853e-16, 
    6.8575e-16, 6.860439e-16, 6.838185e-16, 6.851849e-16, 6.807945e-16, 
    6.815043e-16, 6.81082e-16, 6.795367e-16, 6.844687e-16, 6.819392e-16, 
    6.866073e-16, 6.852394e-16, 6.892284e-16, 6.872455e-16, 6.911375e-16, 
    6.927975e-16, 6.943598e-16, 6.961815e-16, 6.806971e-16, 6.801599e-16, 
    6.811219e-16, 6.824513e-16, 6.836849e-16, 6.853228e-16, 6.854905e-16, 
    6.85797e-16, 6.865911e-16, 6.872584e-16, 6.858936e-16, 6.874256e-16, 
    6.816682e-16, 6.846882e-16, 6.799564e-16, 6.813823e-16, 6.823731e-16, 
    6.819389e-16, 6.841941e-16, 6.847251e-16, 6.868808e-16, 6.85767e-16, 
    6.923877e-16, 6.894619e-16, 6.975682e-16, 6.95307e-16, 6.799721e-16, 
    6.806954e-16, 6.832097e-16, 6.820139e-16, 6.854322e-16, 6.862724e-16, 
    6.869554e-16, 6.878274e-16, 6.879218e-16, 6.884383e-16, 6.875918e-16, 
    6.88405e-16, 6.853263e-16, 6.867028e-16, 6.829229e-16, 6.838435e-16, 
    6.834202e-16, 6.829555e-16, 6.843893e-16, 6.85915e-16, 6.859481e-16, 
    6.864369e-16, 6.878125e-16, 6.854461e-16, 6.927638e-16, 6.882477e-16, 
    6.814837e-16, 6.828746e-16, 6.830738e-16, 6.825351e-16, 6.861882e-16, 
    6.848654e-16, 6.884258e-16, 6.874644e-16, 6.890394e-16, 6.882569e-16, 
    6.881417e-16, 6.871362e-16, 6.865097e-16, 6.84926e-16, 6.836364e-16, 
    6.826133e-16, 6.828513e-16, 6.839749e-16, 6.860084e-16, 6.879301e-16, 
    6.875092e-16, 6.889197e-16, 6.851846e-16, 6.867516e-16, 6.86146e-16, 
    6.877248e-16, 6.842639e-16, 6.872098e-16, 6.835098e-16, 6.838347e-16, 
    6.848392e-16, 6.868575e-16, 6.873045e-16, 6.877806e-16, 6.874869e-16, 
    6.860601e-16, 6.858264e-16, 6.848149e-16, 6.845352e-16, 6.83764e-16, 
    6.83125e-16, 6.837087e-16, 6.843214e-16, 6.860609e-16, 6.876266e-16, 
    6.893321e-16, 6.897494e-16, 6.917378e-16, 6.901186e-16, 6.927889e-16, 
    6.905178e-16, 6.944476e-16, 6.873812e-16, 6.90452e-16, 6.84885e-16, 
    6.854858e-16, 6.865714e-16, 6.890596e-16, 6.877174e-16, 6.892872e-16, 
    6.858173e-16, 6.840134e-16, 6.83547e-16, 6.826754e-16, 6.83567e-16, 
    6.834945e-16, 6.843471e-16, 6.840732e-16, 6.861187e-16, 6.850203e-16, 
    6.881387e-16, 6.89275e-16, 6.924801e-16, 6.944413e-16, 6.96436e-16, 
    6.973155e-16, 6.975831e-16, 6.97695e-16 ;

 CWDC_TO_LITR2C =
  5.137911e-16, 5.151804e-16, 5.149105e-16, 5.160299e-16, 5.154092e-16, 
    5.16142e-16, 5.14073e-16, 5.152353e-16, 5.144936e-16, 5.139165e-16, 
    5.181991e-16, 5.160799e-16, 5.203983e-16, 5.190492e-16, 5.224358e-16, 
    5.201882e-16, 5.228886e-16, 5.223715e-16, 5.239283e-16, 5.234826e-16, 
    5.254707e-16, 5.24134e-16, 5.265007e-16, 5.251519e-16, 5.253628e-16, 
    5.240898e-16, 5.16507e-16, 5.179353e-16, 5.164223e-16, 5.166261e-16, 
    5.165347e-16, 5.154219e-16, 5.148605e-16, 5.136851e-16, 5.138986e-16, 
    5.14762e-16, 5.167177e-16, 5.160545e-16, 5.177262e-16, 5.176885e-16, 
    5.195468e-16, 5.187092e-16, 5.218288e-16, 5.209431e-16, 5.235011e-16, 
    5.228583e-16, 5.234709e-16, 5.232852e-16, 5.234733e-16, 5.225303e-16, 
    5.229344e-16, 5.221044e-16, 5.188661e-16, 5.198186e-16, 5.169754e-16, 
    5.152622e-16, 5.14124e-16, 5.133154e-16, 5.134297e-16, 5.136476e-16, 
    5.147671e-16, 5.158191e-16, 5.166201e-16, 5.171556e-16, 5.17683e-16, 
    5.192772e-16, 5.20121e-16, 5.220076e-16, 5.216677e-16, 5.222438e-16, 
    5.227943e-16, 5.237176e-16, 5.235657e-16, 5.239723e-16, 5.222288e-16, 
    5.233877e-16, 5.21474e-16, 5.219977e-16, 5.17825e-16, 5.162335e-16, 
    5.155552e-16, 5.149623e-16, 5.135176e-16, 5.145154e-16, 5.141221e-16, 
    5.150578e-16, 5.156518e-16, 5.153581e-16, 5.171702e-16, 5.16466e-16, 
    5.20171e-16, 5.185765e-16, 5.227301e-16, 5.217375e-16, 5.229679e-16, 
    5.223403e-16, 5.234154e-16, 5.224479e-16, 5.241237e-16, 5.244881e-16, 
    5.24239e-16, 5.251959e-16, 5.223942e-16, 5.234708e-16, 5.153498e-16, 
    5.153977e-16, 5.15621e-16, 5.146392e-16, 5.145792e-16, 5.136792e-16, 
    5.144802e-16, 5.14821e-16, 5.156864e-16, 5.161977e-16, 5.166837e-16, 
    5.177516e-16, 5.189429e-16, 5.206073e-16, 5.218019e-16, 5.226019e-16, 
    5.221115e-16, 5.225445e-16, 5.220604e-16, 5.218335e-16, 5.243515e-16, 
    5.229381e-16, 5.250583e-16, 5.249412e-16, 5.239819e-16, 5.249543e-16, 
    5.154314e-16, 5.151557e-16, 5.141977e-16, 5.149475e-16, 5.135812e-16, 
    5.14346e-16, 5.147854e-16, 5.164804e-16, 5.168528e-16, 5.171977e-16, 
    5.178787e-16, 5.187521e-16, 5.202826e-16, 5.21613e-16, 5.228264e-16, 
    5.227375e-16, 5.227688e-16, 5.230396e-16, 5.223686e-16, 5.231497e-16, 
    5.232806e-16, 5.229381e-16, 5.249254e-16, 5.24358e-16, 5.249387e-16, 
    5.245693e-16, 5.152454e-16, 5.157092e-16, 5.154586e-16, 5.159298e-16, 
    5.155977e-16, 5.170734e-16, 5.175154e-16, 5.195823e-16, 5.187348e-16, 
    5.200838e-16, 5.188721e-16, 5.190868e-16, 5.201272e-16, 5.189376e-16, 
    5.215394e-16, 5.197756e-16, 5.230501e-16, 5.212904e-16, 5.231603e-16, 
    5.228211e-16, 5.233827e-16, 5.238853e-16, 5.245175e-16, 5.256827e-16, 
    5.254131e-16, 5.263871e-16, 5.164006e-16, 5.170016e-16, 5.16949e-16, 
    5.175778e-16, 5.180426e-16, 5.190498e-16, 5.206632e-16, 5.200568e-16, 
    5.211701e-16, 5.213933e-16, 5.197021e-16, 5.207405e-16, 5.174039e-16, 
    5.179433e-16, 5.176223e-16, 5.164479e-16, 5.201962e-16, 5.182738e-16, 
    5.218215e-16, 5.207819e-16, 5.238136e-16, 5.223066e-16, 5.252646e-16, 
    5.265261e-16, 5.277134e-16, 5.290979e-16, 5.173298e-16, 5.169215e-16, 
    5.176526e-16, 5.18663e-16, 5.196005e-16, 5.208453e-16, 5.209727e-16, 
    5.212057e-16, 5.218092e-16, 5.223164e-16, 5.212791e-16, 5.224435e-16, 
    5.180678e-16, 5.20363e-16, 5.167669e-16, 5.178505e-16, 5.186036e-16, 
    5.182736e-16, 5.199875e-16, 5.20391e-16, 5.220294e-16, 5.211829e-16, 
    5.262146e-16, 5.23991e-16, 5.301518e-16, 5.284333e-16, 5.167788e-16, 
    5.173285e-16, 5.192394e-16, 5.183306e-16, 5.209285e-16, 5.21567e-16, 
    5.220861e-16, 5.227488e-16, 5.228206e-16, 5.23213e-16, 5.225698e-16, 
    5.231878e-16, 5.20848e-16, 5.218942e-16, 5.190214e-16, 5.197211e-16, 
    5.193993e-16, 5.190462e-16, 5.201359e-16, 5.212954e-16, 5.213206e-16, 
    5.21692e-16, 5.227375e-16, 5.20939e-16, 5.265005e-16, 5.230682e-16, 
    5.179276e-16, 5.189847e-16, 5.191361e-16, 5.187267e-16, 5.21503e-16, 
    5.204977e-16, 5.232036e-16, 5.22473e-16, 5.236699e-16, 5.230752e-16, 
    5.229877e-16, 5.222236e-16, 5.217474e-16, 5.205437e-16, 5.195637e-16, 
    5.187861e-16, 5.18967e-16, 5.198209e-16, 5.213664e-16, 5.228269e-16, 
    5.22507e-16, 5.23579e-16, 5.207403e-16, 5.219312e-16, 5.214709e-16, 
    5.226708e-16, 5.200406e-16, 5.222795e-16, 5.194675e-16, 5.197144e-16, 
    5.204778e-16, 5.220117e-16, 5.223514e-16, 5.227133e-16, 5.224901e-16, 
    5.214056e-16, 5.212281e-16, 5.204593e-16, 5.202467e-16, 5.196606e-16, 
    5.19175e-16, 5.196187e-16, 5.200843e-16, 5.214063e-16, 5.225962e-16, 
    5.238924e-16, 5.242095e-16, 5.257207e-16, 5.244901e-16, 5.265195e-16, 
    5.247935e-16, 5.277802e-16, 5.224097e-16, 5.247435e-16, 5.205126e-16, 
    5.209693e-16, 5.217943e-16, 5.236853e-16, 5.226652e-16, 5.238583e-16, 
    5.212211e-16, 5.198502e-16, 5.194957e-16, 5.188333e-16, 5.195109e-16, 
    5.194558e-16, 5.201038e-16, 5.198956e-16, 5.214502e-16, 5.206154e-16, 
    5.229854e-16, 5.23849e-16, 5.262849e-16, 5.277754e-16, 5.292914e-16, 
    5.299598e-16, 5.301632e-16, 5.302482e-16 ;

 CWDC_TO_LITR3C =
  1.622498e-16, 1.626885e-16, 1.626033e-16, 1.629568e-16, 1.627608e-16, 
    1.629922e-16, 1.623389e-16, 1.627059e-16, 1.624717e-16, 1.622894e-16, 
    1.636418e-16, 1.629726e-16, 1.643363e-16, 1.639103e-16, 1.649797e-16, 
    1.6427e-16, 1.651227e-16, 1.649594e-16, 1.654511e-16, 1.653103e-16, 
    1.659381e-16, 1.65516e-16, 1.662634e-16, 1.658374e-16, 1.65904e-16, 
    1.65502e-16, 1.631075e-16, 1.635585e-16, 1.630807e-16, 1.631451e-16, 
    1.631162e-16, 1.627648e-16, 1.625875e-16, 1.622164e-16, 1.622838e-16, 
    1.625564e-16, 1.63174e-16, 1.629646e-16, 1.634925e-16, 1.634806e-16, 
    1.640674e-16, 1.638029e-16, 1.64788e-16, 1.645083e-16, 1.653162e-16, 
    1.651131e-16, 1.653066e-16, 1.65248e-16, 1.653074e-16, 1.650096e-16, 
    1.651372e-16, 1.648751e-16, 1.638524e-16, 1.641532e-16, 1.632554e-16, 
    1.627144e-16, 1.623549e-16, 1.620996e-16, 1.621357e-16, 1.622045e-16, 
    1.62558e-16, 1.628902e-16, 1.631432e-16, 1.633123e-16, 1.634789e-16, 
    1.639823e-16, 1.642487e-16, 1.648445e-16, 1.647372e-16, 1.649191e-16, 
    1.650929e-16, 1.653845e-16, 1.653366e-16, 1.654649e-16, 1.649144e-16, 
    1.652803e-16, 1.64676e-16, 1.648414e-16, 1.635237e-16, 1.630211e-16, 
    1.628069e-16, 1.626197e-16, 1.621635e-16, 1.624785e-16, 1.623544e-16, 
    1.626498e-16, 1.628374e-16, 1.627447e-16, 1.633169e-16, 1.630945e-16, 
    1.642645e-16, 1.63761e-16, 1.650727e-16, 1.647592e-16, 1.651478e-16, 
    1.649496e-16, 1.652891e-16, 1.649835e-16, 1.655127e-16, 1.656278e-16, 
    1.655492e-16, 1.658513e-16, 1.649666e-16, 1.653066e-16, 1.627421e-16, 
    1.627572e-16, 1.628277e-16, 1.625176e-16, 1.624987e-16, 1.622145e-16, 
    1.624674e-16, 1.625751e-16, 1.628483e-16, 1.630098e-16, 1.631633e-16, 
    1.635005e-16, 1.638767e-16, 1.644023e-16, 1.647795e-16, 1.650322e-16, 
    1.648773e-16, 1.65014e-16, 1.648612e-16, 1.647895e-16, 1.655847e-16, 
    1.651384e-16, 1.658079e-16, 1.657709e-16, 1.65468e-16, 1.657751e-16, 
    1.627678e-16, 1.626808e-16, 1.623782e-16, 1.62615e-16, 1.621835e-16, 
    1.62425e-16, 1.625638e-16, 1.630991e-16, 1.632167e-16, 1.633256e-16, 
    1.635407e-16, 1.638164e-16, 1.642998e-16, 1.647199e-16, 1.651031e-16, 
    1.65075e-16, 1.650849e-16, 1.651704e-16, 1.649585e-16, 1.652052e-16, 
    1.652465e-16, 1.651384e-16, 1.657659e-16, 1.655867e-16, 1.657701e-16, 
    1.656535e-16, 1.627091e-16, 1.628556e-16, 1.627764e-16, 1.629252e-16, 
    1.628203e-16, 1.632863e-16, 1.634259e-16, 1.640786e-16, 1.63811e-16, 
    1.64237e-16, 1.638543e-16, 1.639221e-16, 1.642507e-16, 1.638751e-16, 
    1.646967e-16, 1.641397e-16, 1.651737e-16, 1.64618e-16, 1.652085e-16, 
    1.651014e-16, 1.652787e-16, 1.654375e-16, 1.656371e-16, 1.660051e-16, 
    1.659199e-16, 1.662275e-16, 1.630739e-16, 1.632637e-16, 1.63247e-16, 
    1.634456e-16, 1.635924e-16, 1.639105e-16, 1.644199e-16, 1.642285e-16, 
    1.6458e-16, 1.646505e-16, 1.641164e-16, 1.644444e-16, 1.633907e-16, 
    1.63561e-16, 1.634597e-16, 1.630888e-16, 1.642725e-16, 1.636654e-16, 
    1.647857e-16, 1.644575e-16, 1.654148e-16, 1.649389e-16, 1.65873e-16, 
    1.662714e-16, 1.666463e-16, 1.670835e-16, 1.633673e-16, 1.632384e-16, 
    1.634693e-16, 1.637883e-16, 1.640844e-16, 1.644775e-16, 1.645177e-16, 
    1.645913e-16, 1.647819e-16, 1.64942e-16, 1.646145e-16, 1.649822e-16, 
    1.636004e-16, 1.643252e-16, 1.631896e-16, 1.635317e-16, 1.637696e-16, 
    1.636653e-16, 1.642066e-16, 1.64334e-16, 1.648514e-16, 1.645841e-16, 
    1.66173e-16, 1.654709e-16, 1.674164e-16, 1.668737e-16, 1.631933e-16, 
    1.633669e-16, 1.639703e-16, 1.636833e-16, 1.645037e-16, 1.647054e-16, 
    1.648693e-16, 1.650786e-16, 1.651012e-16, 1.652252e-16, 1.65022e-16, 
    1.652172e-16, 1.644783e-16, 1.648087e-16, 1.639015e-16, 1.641225e-16, 
    1.640208e-16, 1.639093e-16, 1.642534e-16, 1.646196e-16, 1.646276e-16, 
    1.647449e-16, 1.65075e-16, 1.645071e-16, 1.662633e-16, 1.651794e-16, 
    1.635561e-16, 1.638899e-16, 1.639377e-16, 1.638084e-16, 1.646852e-16, 
    1.643677e-16, 1.652222e-16, 1.649915e-16, 1.653694e-16, 1.651817e-16, 
    1.65154e-16, 1.649127e-16, 1.647623e-16, 1.643822e-16, 1.640727e-16, 
    1.638272e-16, 1.638843e-16, 1.64154e-16, 1.64642e-16, 1.651032e-16, 
    1.650022e-16, 1.653407e-16, 1.644443e-16, 1.648204e-16, 1.64675e-16, 
    1.650539e-16, 1.642233e-16, 1.649304e-16, 1.640424e-16, 1.641203e-16, 
    1.643614e-16, 1.648458e-16, 1.649531e-16, 1.650673e-16, 1.649969e-16, 
    1.646544e-16, 1.645983e-16, 1.643556e-16, 1.642884e-16, 1.641034e-16, 
    1.6395e-16, 1.640901e-16, 1.642371e-16, 1.646546e-16, 1.650304e-16, 
    1.654397e-16, 1.655398e-16, 1.660171e-16, 1.656285e-16, 1.662693e-16, 
    1.657243e-16, 1.666674e-16, 1.649715e-16, 1.657085e-16, 1.643724e-16, 
    1.645166e-16, 1.647771e-16, 1.653743e-16, 1.650522e-16, 1.654289e-16, 
    1.645962e-16, 1.641632e-16, 1.640513e-16, 1.638421e-16, 1.640561e-16, 
    1.640387e-16, 1.642433e-16, 1.641776e-16, 1.646685e-16, 1.644049e-16, 
    1.651533e-16, 1.65426e-16, 1.661952e-16, 1.666659e-16, 1.671446e-16, 
    1.673557e-16, 1.6742e-16, 1.674468e-16 ;

 CWDC_vr =
  5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  1.027582e-18, 1.030361e-18, 1.029821e-18, 1.03206e-18, 1.030818e-18, 
    1.032284e-18, 1.028146e-18, 1.030471e-18, 1.028987e-18, 1.027833e-18, 
    1.036398e-18, 1.03216e-18, 1.040797e-18, 1.038099e-18, 1.044872e-18, 
    1.040376e-18, 1.045777e-18, 1.044743e-18, 1.047857e-18, 1.046965e-18, 
    1.050941e-18, 1.048268e-18, 1.053001e-18, 1.050304e-18, 1.050726e-18, 
    1.04818e-18, 1.033014e-18, 1.035871e-18, 1.032845e-18, 1.033252e-18, 
    1.033069e-18, 1.030844e-18, 1.029721e-18, 1.02737e-18, 1.027797e-18, 
    1.029524e-18, 1.033435e-18, 1.032109e-18, 1.035452e-18, 1.035377e-18, 
    1.039094e-18, 1.037418e-18, 1.043658e-18, 1.041886e-18, 1.047002e-18, 
    1.045717e-18, 1.046942e-18, 1.04657e-18, 1.046947e-18, 1.045061e-18, 
    1.045869e-18, 1.044209e-18, 1.037732e-18, 1.039637e-18, 1.033951e-18, 
    1.030524e-18, 1.028248e-18, 1.026631e-18, 1.026859e-18, 1.027295e-18, 
    1.029534e-18, 1.031638e-18, 1.03324e-18, 1.034311e-18, 1.035366e-18, 
    1.038554e-18, 1.040242e-18, 1.044015e-18, 1.043335e-18, 1.044487e-18, 
    1.045589e-18, 1.047435e-18, 1.047132e-18, 1.047945e-18, 1.044458e-18, 
    1.046775e-18, 1.042948e-18, 1.043995e-18, 1.03565e-18, 1.032467e-18, 
    1.031111e-18, 1.029925e-18, 1.027035e-18, 1.029031e-18, 1.028244e-18, 
    1.030116e-18, 1.031304e-18, 1.030716e-18, 1.03434e-18, 1.032932e-18, 
    1.040342e-18, 1.037153e-18, 1.04546e-18, 1.043475e-18, 1.045936e-18, 
    1.044681e-18, 1.046831e-18, 1.044896e-18, 1.048247e-18, 1.048976e-18, 
    1.048478e-18, 1.050392e-18, 1.044788e-18, 1.046942e-18, 1.0307e-18, 
    1.030795e-18, 1.031242e-18, 1.029278e-18, 1.029158e-18, 1.027358e-18, 
    1.02896e-18, 1.029642e-18, 1.031373e-18, 1.032395e-18, 1.033367e-18, 
    1.035503e-18, 1.037886e-18, 1.041215e-18, 1.043604e-18, 1.045204e-18, 
    1.044223e-18, 1.045089e-18, 1.044121e-18, 1.043667e-18, 1.048703e-18, 
    1.045876e-18, 1.050117e-18, 1.049882e-18, 1.047964e-18, 1.049909e-18, 
    1.030863e-18, 1.030311e-18, 1.028395e-18, 1.029895e-18, 1.027162e-18, 
    1.028692e-18, 1.029571e-18, 1.032961e-18, 1.033706e-18, 1.034395e-18, 
    1.035758e-18, 1.037504e-18, 1.040565e-18, 1.043226e-18, 1.045653e-18, 
    1.045475e-18, 1.045538e-18, 1.046079e-18, 1.044737e-18, 1.046299e-18, 
    1.046561e-18, 1.045876e-18, 1.049851e-18, 1.048716e-18, 1.049877e-18, 
    1.049139e-18, 1.030491e-18, 1.031419e-18, 1.030917e-18, 1.03186e-18, 
    1.031196e-18, 1.034147e-18, 1.035031e-18, 1.039165e-18, 1.03747e-18, 
    1.040168e-18, 1.037744e-18, 1.038174e-18, 1.040254e-18, 1.037875e-18, 
    1.043079e-18, 1.039551e-18, 1.0461e-18, 1.042581e-18, 1.046321e-18, 
    1.045642e-18, 1.046765e-18, 1.047771e-18, 1.049035e-18, 1.051365e-18, 
    1.050826e-18, 1.052774e-18, 1.032801e-18, 1.034003e-18, 1.033898e-18, 
    1.035156e-18, 1.036085e-18, 1.0381e-18, 1.041326e-18, 1.040114e-18, 
    1.04234e-18, 1.042787e-18, 1.039404e-18, 1.041481e-18, 1.034808e-18, 
    1.035887e-18, 1.035245e-18, 1.032896e-18, 1.040392e-18, 1.036548e-18, 
    1.043643e-18, 1.041564e-18, 1.047627e-18, 1.044613e-18, 1.050529e-18, 
    1.053052e-18, 1.055427e-18, 1.058196e-18, 1.03466e-18, 1.033843e-18, 
    1.035305e-18, 1.037326e-18, 1.039201e-18, 1.041691e-18, 1.041945e-18, 
    1.042411e-18, 1.043619e-18, 1.044633e-18, 1.042558e-18, 1.044887e-18, 
    1.036136e-18, 1.040726e-18, 1.033534e-18, 1.035701e-18, 1.037207e-18, 
    1.036547e-18, 1.039975e-18, 1.040782e-18, 1.044059e-18, 1.042366e-18, 
    1.052429e-18, 1.047982e-18, 1.060304e-18, 1.056867e-18, 1.033558e-18, 
    1.034657e-18, 1.038479e-18, 1.036661e-18, 1.041857e-18, 1.043134e-18, 
    1.044172e-18, 1.045498e-18, 1.045641e-18, 1.046426e-18, 1.045139e-18, 
    1.046376e-18, 1.041696e-18, 1.043788e-18, 1.038043e-18, 1.039442e-18, 
    1.038799e-18, 1.038092e-18, 1.040272e-18, 1.042591e-18, 1.042641e-18, 
    1.043384e-18, 1.045475e-18, 1.041878e-18, 1.053001e-18, 1.046136e-18, 
    1.035855e-18, 1.037969e-18, 1.038272e-18, 1.037453e-18, 1.043006e-18, 
    1.040995e-18, 1.046407e-18, 1.044946e-18, 1.04734e-18, 1.046151e-18, 
    1.045975e-18, 1.044447e-18, 1.043495e-18, 1.041087e-18, 1.039127e-18, 
    1.037572e-18, 1.037934e-18, 1.039642e-18, 1.042733e-18, 1.045654e-18, 
    1.045014e-18, 1.047158e-18, 1.041481e-18, 1.043862e-18, 1.042942e-18, 
    1.045342e-18, 1.040081e-18, 1.044559e-18, 1.038935e-18, 1.039429e-18, 
    1.040956e-18, 1.044023e-18, 1.044703e-18, 1.045427e-18, 1.04498e-18, 
    1.042811e-18, 1.042456e-18, 1.040919e-18, 1.040494e-18, 1.039321e-18, 
    1.03835e-18, 1.039237e-18, 1.040168e-18, 1.042813e-18, 1.045192e-18, 
    1.047785e-18, 1.048419e-18, 1.051441e-18, 1.04898e-18, 1.053039e-18, 
    1.049587e-18, 1.05556e-18, 1.044819e-18, 1.049487e-18, 1.041025e-18, 
    1.041939e-18, 1.043589e-18, 1.047371e-18, 1.04533e-18, 1.047717e-18, 
    1.042442e-18, 1.0397e-18, 1.038991e-18, 1.037667e-18, 1.039022e-18, 
    1.038912e-18, 1.040208e-18, 1.039791e-18, 1.0429e-18, 1.041231e-18, 
    1.045971e-18, 1.047698e-18, 1.05257e-18, 1.055551e-18, 1.058583e-18, 
    1.05992e-18, 1.060326e-18, 1.060496e-18 ;

 CWDN_TO_LITR3N =
  3.244996e-19, 3.253771e-19, 3.252066e-19, 3.259136e-19, 3.255216e-19, 
    3.259844e-19, 3.246777e-19, 3.254118e-19, 3.249433e-19, 3.245788e-19, 
    3.272836e-19, 3.259452e-19, 3.286726e-19, 3.278206e-19, 3.299595e-19, 
    3.285399e-19, 3.302454e-19, 3.299188e-19, 3.309021e-19, 3.306205e-19, 
    3.318762e-19, 3.31032e-19, 3.325267e-19, 3.316748e-19, 3.318081e-19, 
    3.310041e-19, 3.26215e-19, 3.27117e-19, 3.261615e-19, 3.262902e-19, 
    3.262325e-19, 3.255296e-19, 3.25175e-19, 3.244327e-19, 3.245676e-19, 
    3.251129e-19, 3.26348e-19, 3.259291e-19, 3.26985e-19, 3.269611e-19, 
    3.281348e-19, 3.276058e-19, 3.295761e-19, 3.290167e-19, 3.306323e-19, 
    3.302263e-19, 3.306132e-19, 3.304959e-19, 3.306147e-19, 3.300192e-19, 
    3.302744e-19, 3.297502e-19, 3.277049e-19, 3.283065e-19, 3.265108e-19, 
    3.254288e-19, 3.247099e-19, 3.241992e-19, 3.242714e-19, 3.24409e-19, 
    3.251161e-19, 3.257805e-19, 3.262864e-19, 3.266246e-19, 3.269577e-19, 
    3.279645e-19, 3.284975e-19, 3.29689e-19, 3.294743e-19, 3.298382e-19, 
    3.301859e-19, 3.30769e-19, 3.306731e-19, 3.309299e-19, 3.298287e-19, 
    3.305606e-19, 3.29352e-19, 3.296827e-19, 3.270474e-19, 3.260422e-19, 
    3.256138e-19, 3.252394e-19, 3.243269e-19, 3.249571e-19, 3.247087e-19, 
    3.252997e-19, 3.256749e-19, 3.254894e-19, 3.266338e-19, 3.261891e-19, 
    3.28529e-19, 3.27522e-19, 3.301453e-19, 3.295184e-19, 3.302955e-19, 
    3.298991e-19, 3.305782e-19, 3.299671e-19, 3.310255e-19, 3.312556e-19, 
    3.310983e-19, 3.317027e-19, 3.299332e-19, 3.306131e-19, 3.254841e-19, 
    3.255144e-19, 3.256554e-19, 3.250353e-19, 3.249974e-19, 3.24429e-19, 
    3.249348e-19, 3.251501e-19, 3.256967e-19, 3.260196e-19, 3.263266e-19, 
    3.27001e-19, 3.277534e-19, 3.288046e-19, 3.295591e-19, 3.300643e-19, 
    3.297546e-19, 3.300281e-19, 3.297223e-19, 3.295791e-19, 3.311693e-19, 
    3.302767e-19, 3.316158e-19, 3.315418e-19, 3.309359e-19, 3.315501e-19, 
    3.255356e-19, 3.253615e-19, 3.247564e-19, 3.2523e-19, 3.243671e-19, 
    3.248501e-19, 3.251276e-19, 3.261982e-19, 3.264334e-19, 3.266512e-19, 
    3.270813e-19, 3.276329e-19, 3.285996e-19, 3.294398e-19, 3.302062e-19, 
    3.3015e-19, 3.301698e-19, 3.303408e-19, 3.29917e-19, 3.304104e-19, 
    3.30493e-19, 3.302767e-19, 3.315319e-19, 3.311735e-19, 3.315402e-19, 
    3.313069e-19, 3.254181e-19, 3.257111e-19, 3.255528e-19, 3.258504e-19, 
    3.256407e-19, 3.265726e-19, 3.268519e-19, 3.281573e-19, 3.27622e-19, 
    3.28474e-19, 3.277087e-19, 3.278443e-19, 3.285014e-19, 3.277501e-19, 
    3.293933e-19, 3.282793e-19, 3.303475e-19, 3.29236e-19, 3.30417e-19, 
    3.302028e-19, 3.305575e-19, 3.308749e-19, 3.312742e-19, 3.320102e-19, 
    3.318398e-19, 3.32455e-19, 3.261478e-19, 3.265273e-19, 3.264941e-19, 
    3.268912e-19, 3.271848e-19, 3.278209e-19, 3.288399e-19, 3.284569e-19, 
    3.2916e-19, 3.29301e-19, 3.282329e-19, 3.288887e-19, 3.267814e-19, 
    3.271221e-19, 3.269194e-19, 3.261776e-19, 3.28545e-19, 3.273308e-19, 
    3.295715e-19, 3.289149e-19, 3.308296e-19, 3.298778e-19, 3.31746e-19, 
    3.325428e-19, 3.332927e-19, 3.341671e-19, 3.267346e-19, 3.264767e-19, 
    3.269385e-19, 3.275766e-19, 3.281687e-19, 3.289549e-19, 3.290354e-19, 
    3.291825e-19, 3.295637e-19, 3.29884e-19, 3.292289e-19, 3.299643e-19, 
    3.272007e-19, 3.286503e-19, 3.263791e-19, 3.270635e-19, 3.275391e-19, 
    3.273307e-19, 3.284132e-19, 3.28668e-19, 3.297028e-19, 3.291681e-19, 
    3.323461e-19, 3.309417e-19, 3.348327e-19, 3.337474e-19, 3.263866e-19, 
    3.267338e-19, 3.279407e-19, 3.273667e-19, 3.290075e-19, 3.294107e-19, 
    3.297386e-19, 3.301571e-19, 3.302025e-19, 3.304504e-19, 3.300441e-19, 
    3.304344e-19, 3.289566e-19, 3.296174e-19, 3.27803e-19, 3.282449e-19, 
    3.280417e-19, 3.278186e-19, 3.285069e-19, 3.292392e-19, 3.292551e-19, 
    3.294897e-19, 3.3015e-19, 3.290141e-19, 3.325267e-19, 3.303589e-19, 
    3.271122e-19, 3.277798e-19, 3.278754e-19, 3.276168e-19, 3.293703e-19, 
    3.287354e-19, 3.304444e-19, 3.299829e-19, 3.307389e-19, 3.303633e-19, 
    3.30308e-19, 3.298254e-19, 3.295247e-19, 3.287645e-19, 3.281455e-19, 
    3.276544e-19, 3.277686e-19, 3.28308e-19, 3.29284e-19, 3.302064e-19, 
    3.300044e-19, 3.306815e-19, 3.288886e-19, 3.296408e-19, 3.293501e-19, 
    3.301079e-19, 3.284467e-19, 3.298607e-19, 3.280847e-19, 3.282407e-19, 
    3.287228e-19, 3.296916e-19, 3.299061e-19, 3.301347e-19, 3.299937e-19, 
    3.293088e-19, 3.291967e-19, 3.287111e-19, 3.285769e-19, 3.282067e-19, 
    3.279e-19, 3.281802e-19, 3.284743e-19, 3.293092e-19, 3.300608e-19, 
    3.308794e-19, 3.310797e-19, 3.320341e-19, 3.312569e-19, 3.325387e-19, 
    3.314485e-19, 3.333349e-19, 3.29943e-19, 3.31417e-19, 3.287448e-19, 
    3.290332e-19, 3.295543e-19, 3.307486e-19, 3.301043e-19, 3.308579e-19, 
    3.291923e-19, 3.283264e-19, 3.281026e-19, 3.276842e-19, 3.281122e-19, 
    3.280774e-19, 3.284866e-19, 3.283551e-19, 3.293369e-19, 3.288097e-19, 
    3.303066e-19, 3.30852e-19, 3.323905e-19, 3.333319e-19, 3.342893e-19, 
    3.347114e-19, 3.348399e-19, 3.348936e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.100726e-43, 5.605194e-45, 
    3.498145e-40, 2.53635e-43, 1.405053e-39, 2.860358e-40, 3.155876e-38, 
    8.419162e-39, 2.624818e-36, 5.766906e-38, 4.399989e-35, 1.071883e-36, 
    1.939966e-36, 5.068994e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.942727e-44, 1.401298e-45, 5.228945e-41, 3.049225e-42, 8.900133e-39, 
    1.278835e-39, 8.133579e-39, 4.660608e-39, 8.192598e-39, 4.676525e-40, 
    1.613396e-39, 1.244143e-40, 2.802597e-45, 7.286752e-44, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.121039e-44, 2.031883e-43, 9.19462e-41, 3.137227e-41, 
    1.924305e-40, 1.051815e-39, 1.695091e-38, 1.079296e-38, 3.593701e-38, 
    1.834622e-40, 6.345298e-39, 1.690947e-41, 8.899506e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.39622e-43, 1.401298e-45, 8.642228e-40, 3.915788e-41, 
    1.785855e-39, 2.594924e-40, 6.893387e-39, 3.6223e-40, 5.59756e-38, 
    1.61379e-37, 7.839023e-38, 1.212262e-36, 3.067653e-40, 8.134899e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.203895e-45, 1.017343e-42, 
    4.801269e-41, 5.826459e-40, 1.27116e-40, 4.881381e-40, 1.083344e-40, 
    5.302794e-41, 1.08715e-37, 1.632183e-39, 8.222793e-37, 5.898124e-37, 
    3.697471e-38, 6.123528e-37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.401298e-45, 3.47522e-43, 2.638505e-41, 1.15981e-39, 8.837471e-40, 
    9.726132e-40, 2.220196e-39, 2.83372e-40, 3.098589e-39, 4.600644e-39, 
    1.630998e-39, 5.640851e-37, 1.106896e-37, 5.856523e-37, 2.036912e-37, 0, 
    0, 0, 0, 0, 0, 0, 3.222986e-44, 1.401298e-45, 1.793662e-43, 2.802597e-45, 
    5.605194e-45, 2.073922e-43, 4.203895e-45, 2.089476e-41, 6.305843e-44, 
    2.292201e-39, 9.419528e-42, 3.198822e-39, 1.14138e-39, 6.244441e-39, 
    2.781966e-38, 1.755172e-37, 4.722894e-36, 2.230228e-36, 3.237457e-35, 0, 
    0, 0, 0, 0, 5.605194e-45, 1.221932e-42, 1.625506e-43, 6.366099e-42, 
    1.306851e-41, 4.904545e-44, 1.575059e-42, 0, 0, 0, 0, 2.606415e-43, 0, 
    5.110676e-41, 1.80207e-42, 2.251942e-38, 2.340813e-40, 1.471128e-36, 
    4.718157e-35, 1.069506e-33, 3.474821e-32, 0, 0, 0, 1.401298e-45, 
    3.503246e-44, 2.218255e-42, 3.358912e-42, 7.146622e-42, 4.912392e-41, 
    2.409084e-40, 9.066401e-42, 3.573101e-40, 0, 4.540207e-43, 0, 0, 
    1.401298e-45, 0, 1.289195e-43, 4.97461e-43, 9.84216e-41, 6.63655e-42, 
    2.034721e-35, 3.803153e-38, 4.371386e-31, 6.681893e-33, 0, 0, 
    9.809089e-45, 0, 2.907694e-42, 2.277671e-41, 1.173952e-40, 9.156785e-40, 
    1.139511e-39, 3.752387e-39, 5.277444e-40, 3.475073e-39, 2.237874e-42, 
    6.425234e-41, 4.203895e-45, 5.324934e-44, 1.821688e-44, 5.605194e-45, 
    2.129974e-43, 9.555454e-42, 1.034298e-41, 3.392263e-41, 8.898455e-40, 
    3.009989e-42, 4.420301e-35, 2.435304e-39, 0, 4.203895e-45, 7.006492e-45, 
    1.401298e-45, 1.856861e-41, 7.076557e-43, 3.645385e-39, 3.914247e-40, 
    1.470874e-38, 2.473112e-39, 1.896537e-39, 1.804298e-40, 4.040644e-41, 
    8.239635e-43, 3.082857e-44, 1.401298e-45, 4.203895e-45, 7.426882e-44, 
    1.200072e-41, 1.162563e-39, 4.354619e-40, 1.122507e-38, 1.572257e-42, 
    7.226917e-41, 1.677214e-41, 7.204426e-40, 1.541428e-43, 2.160732e-40, 
    2.242078e-44, 5.184804e-44, 6.628142e-43, 9.319896e-41, 2.685967e-40, 
    8.211385e-40, 4.12688e-40, 1.360801e-41, 7.683319e-42, 6.235778e-43, 
    3.082857e-43, 4.344025e-44, 8.407791e-45, 3.643376e-44, 1.793662e-43, 
    1.362482e-41, 5.731339e-40, 2.841443e-38, 7.189204e-38, 5.260623e-36, 
    1.626792e-37, 4.653514e-35, 3.901921e-37, 1.275646e-33, 3.229811e-40, 
    3.37117e-37, 7.426882e-43, 3.319676e-42, 4.69449e-41, 1.543183e-38, 
    7.080719e-40, 2.572929e-38, 7.512361e-42, 8.127531e-44, 2.382207e-44, 
    2.802597e-45, 2.522337e-44, 2.101948e-44, 1.905766e-43, 9.52883e-44, 
    1.568053e-41, 1.042566e-42, 1.884194e-39, 2.502087e-38, 2.457097e-35, 
    1.256787e-33, 5.56119e-32, 2.773154e-31, 4.486484e-31, 5.4801e-31 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  22.1825, 22.24694, 22.23443, 22.28639, 22.25759, 22.2916, 22.1956, 
    22.24946, 22.21509, 22.18835, 22.3872, 22.28872, 22.49, 22.42704, 
    22.58541, 22.48015, 22.60666, 22.58246, 22.65555, 22.63461, 22.72797, 
    22.66522, 22.77655, 22.71303, 22.72293, 22.66313, 22.30861, 22.37491, 
    22.30466, 22.31412, 22.3099, 22.25816, 22.23204, 22.17764, 22.18753, 
    22.22752, 22.31837, 22.28758, 22.36539, 22.36363, 22.45027, 22.4112, 
    22.55702, 22.51557, 22.63549, 22.6053, 22.63405, 22.62534, 22.63416, 
    22.5899, 22.60886, 22.56995, 22.4185, 22.46295, 22.33039, 22.25064, 
    22.19794, 22.16051, 22.1658, 22.17587, 22.22775, 22.27664, 22.31389, 
    22.33881, 22.36337, 22.43756, 22.47704, 22.56536, 22.54949, 22.57644, 
    22.6023, 22.64563, 22.63851, 22.65759, 22.57579, 22.63011, 22.54044, 
    22.56495, 22.36975, 22.2959, 22.26427, 22.23682, 22.16986, 22.21608, 
    22.19785, 22.24129, 22.26887, 22.25524, 22.33949, 22.30671, 22.47938, 
    22.40496, 22.59929, 22.55276, 22.61045, 22.58102, 22.63143, 22.58606, 
    22.66471, 22.68181, 22.67012, 22.71515, 22.58354, 22.63402, 22.25484, 
    22.25706, 22.26744, 22.22182, 22.21904, 22.17735, 22.21447, 22.23027, 
    22.27049, 22.29423, 22.31683, 22.36654, 22.42205, 22.49981, 22.55577, 
    22.59329, 22.5703, 22.59059, 22.5679, 22.55728, 22.67538, 22.60902, 
    22.70867, 22.70316, 22.65803, 22.70378, 22.25863, 22.24584, 22.20136, 
    22.23617, 22.17282, 22.20823, 22.22858, 22.30733, 22.32472, 22.34075, 
    22.37248, 22.41319, 22.48464, 22.5469, 22.60382, 22.59965, 22.60112, 
    22.61381, 22.58234, 22.61897, 22.6251, 22.60905, 22.70242, 22.67574, 
    22.70304, 22.68568, 22.25, 22.27154, 22.2599, 22.28177, 22.26633, 
    22.33491, 22.35547, 22.45188, 22.41237, 22.47533, 22.41879, 22.42879, 
    22.47726, 22.42187, 22.54341, 22.46087, 22.6143, 22.53169, 22.61947, 
    22.60357, 22.62993, 22.65351, 22.68323, 22.73802, 22.72534, 22.77123, 
    22.30367, 22.3316, 22.32919, 22.35846, 22.3801, 22.4271, 22.50245, 
    22.47412, 22.5262, 22.53664, 22.45756, 22.50605, 22.35033, 22.37541, 
    22.36052, 22.30584, 22.48057, 22.39082, 22.55668, 22.50802, 22.65014, 
    22.57937, 22.71835, 22.77768, 22.83382, 22.89915, 22.3469, 22.32792, 
    22.36196, 22.40898, 22.45279, 22.51098, 22.51696, 22.52785, 22.55614, 
    22.5799, 22.53124, 22.58586, 22.38111, 22.4884, 22.32069, 22.37108, 
    22.40623, 22.39087, 22.4709, 22.48976, 22.5664, 22.5268, 22.76298, 
    22.65841, 22.94911, 22.86775, 22.32127, 22.34686, 22.4359, 22.39353, 
    22.51489, 22.54477, 22.56911, 22.60014, 22.60354, 22.62194, 22.59178, 
    22.62077, 22.5111, 22.5601, 22.42578, 22.45842, 22.44343, 22.42694, 
    22.47783, 22.53199, 22.53324, 22.5506, 22.59937, 22.51539, 22.77631, 
    22.61492, 22.37477, 22.42397, 22.43111, 22.41203, 22.54177, 22.49472, 
    22.6215, 22.58724, 22.64341, 22.61548, 22.61137, 22.57554, 22.55322, 
    22.49686, 22.45106, 22.41481, 22.42324, 22.46307, 22.53533, 22.6038, 
    22.58879, 22.63914, 22.50608, 22.5618, 22.54023, 22.59651, 22.47335, 
    22.57793, 22.44661, 22.45813, 22.49379, 22.56552, 22.58154, 22.59847, 
    22.58804, 22.53718, 22.52889, 22.49295, 22.48298, 22.45563, 22.43295, 
    22.45365, 22.47537, 22.53724, 22.59298, 22.65383, 22.66876, 22.73968, 
    22.68182, 22.77719, 22.69591, 22.83676, 22.58413, 22.6937, 22.49545, 
    22.5168, 22.55535, 22.64403, 22.59624, 22.65218, 22.52857, 22.4644, 
    22.44792, 22.41699, 22.44863, 22.44606, 22.47634, 22.46661, 22.5393, 
    22.50025, 22.61124, 22.65176, 22.76638, 22.83666, 22.90841, 22.94004, 
    22.94968, 22.95371 ;

 EFLX_LH_TOT_R =
  22.1825, 22.24694, 22.23443, 22.28639, 22.25759, 22.2916, 22.1956, 
    22.24946, 22.21509, 22.18835, 22.3872, 22.28872, 22.49, 22.42704, 
    22.58541, 22.48015, 22.60666, 22.58246, 22.65555, 22.63461, 22.72797, 
    22.66522, 22.77655, 22.71303, 22.72293, 22.66313, 22.30861, 22.37491, 
    22.30466, 22.31412, 22.3099, 22.25816, 22.23204, 22.17764, 22.18753, 
    22.22752, 22.31837, 22.28758, 22.36539, 22.36363, 22.45027, 22.4112, 
    22.55702, 22.51557, 22.63549, 22.6053, 22.63405, 22.62534, 22.63416, 
    22.5899, 22.60886, 22.56995, 22.4185, 22.46295, 22.33039, 22.25064, 
    22.19794, 22.16051, 22.1658, 22.17587, 22.22775, 22.27664, 22.31389, 
    22.33881, 22.36337, 22.43756, 22.47704, 22.56536, 22.54949, 22.57644, 
    22.6023, 22.64563, 22.63851, 22.65759, 22.57579, 22.63011, 22.54044, 
    22.56495, 22.36975, 22.2959, 22.26427, 22.23682, 22.16986, 22.21608, 
    22.19785, 22.24129, 22.26887, 22.25524, 22.33949, 22.30671, 22.47938, 
    22.40496, 22.59929, 22.55276, 22.61045, 22.58102, 22.63143, 22.58606, 
    22.66471, 22.68181, 22.67012, 22.71515, 22.58354, 22.63402, 22.25484, 
    22.25706, 22.26744, 22.22182, 22.21904, 22.17735, 22.21447, 22.23027, 
    22.27049, 22.29423, 22.31683, 22.36654, 22.42205, 22.49981, 22.55577, 
    22.59329, 22.5703, 22.59059, 22.5679, 22.55728, 22.67538, 22.60902, 
    22.70867, 22.70316, 22.65803, 22.70378, 22.25863, 22.24584, 22.20136, 
    22.23617, 22.17282, 22.20823, 22.22858, 22.30733, 22.32472, 22.34075, 
    22.37248, 22.41319, 22.48464, 22.5469, 22.60382, 22.59965, 22.60112, 
    22.61381, 22.58234, 22.61897, 22.6251, 22.60905, 22.70242, 22.67574, 
    22.70304, 22.68568, 22.25, 22.27154, 22.2599, 22.28177, 22.26633, 
    22.33491, 22.35547, 22.45188, 22.41237, 22.47533, 22.41879, 22.42879, 
    22.47726, 22.42187, 22.54341, 22.46087, 22.6143, 22.53169, 22.61947, 
    22.60357, 22.62993, 22.65351, 22.68323, 22.73802, 22.72534, 22.77123, 
    22.30367, 22.3316, 22.32919, 22.35846, 22.3801, 22.4271, 22.50245, 
    22.47412, 22.5262, 22.53664, 22.45756, 22.50605, 22.35033, 22.37541, 
    22.36052, 22.30584, 22.48057, 22.39082, 22.55668, 22.50802, 22.65014, 
    22.57937, 22.71835, 22.77768, 22.83382, 22.89915, 22.3469, 22.32792, 
    22.36196, 22.40898, 22.45279, 22.51098, 22.51696, 22.52785, 22.55614, 
    22.5799, 22.53124, 22.58586, 22.38111, 22.4884, 22.32069, 22.37108, 
    22.40623, 22.39087, 22.4709, 22.48976, 22.5664, 22.5268, 22.76298, 
    22.65841, 22.94911, 22.86775, 22.32127, 22.34686, 22.4359, 22.39353, 
    22.51489, 22.54477, 22.56911, 22.60014, 22.60354, 22.62194, 22.59178, 
    22.62077, 22.5111, 22.5601, 22.42578, 22.45842, 22.44343, 22.42694, 
    22.47783, 22.53199, 22.53324, 22.5506, 22.59937, 22.51539, 22.77631, 
    22.61492, 22.37477, 22.42397, 22.43111, 22.41203, 22.54177, 22.49472, 
    22.6215, 22.58724, 22.64341, 22.61548, 22.61137, 22.57554, 22.55322, 
    22.49686, 22.45106, 22.41481, 22.42324, 22.46307, 22.53533, 22.6038, 
    22.58879, 22.63914, 22.50608, 22.5618, 22.54023, 22.59651, 22.47335, 
    22.57793, 22.44661, 22.45813, 22.49379, 22.56552, 22.58154, 22.59847, 
    22.58804, 22.53718, 22.52889, 22.49295, 22.48298, 22.45563, 22.43295, 
    22.45365, 22.47537, 22.53724, 22.59298, 22.65383, 22.66876, 22.73968, 
    22.68182, 22.77719, 22.69591, 22.83676, 22.58413, 22.6937, 22.49545, 
    22.5168, 22.55535, 22.64403, 22.59624, 22.65218, 22.52857, 22.4644, 
    22.44792, 22.41699, 22.44863, 22.44606, 22.47634, 22.46661, 22.5393, 
    22.50025, 22.61124, 22.65176, 22.76638, 22.83666, 22.90841, 22.94004, 
    22.94968, 22.95371 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 ERRH2O =
  -22916.25, -22950.76, -22944, -22972.22, -22956.51, -22975.07, -22923.19, 
    -22952.15, -22933.6, -22919.32, -23028.23, -22973.49, -23086.8, -23050.6, 
    -23142.21, -23081.12, -23154.76, -23140.42, -23183.97, -23171.37, 
    -23228.43, -23189.82, -23258.83, -23219.12, -23225.26, -23188.56, 
    -22984.39, -23021.34, -22982.22, -22987.45, -22985.1, -22956.84, 
    -22942.76, -22913.64, -22918.89, -22940.29, -22989.8, -22972.84, 
    -23015.86, -23014.88, -23063.85, -23041.59, -23125.52, -23101.51, 
    -23171.89, -23153.9, -23171.04, -23165.83, -23171.11, -23144.8, 
    -23156.02, -23133.07, -23045.74, -23071.14, -22996.44, -22952.84, 
    -22924.45, -22904.58, -22907.38, -22912.72, -22940.42, -22966.86, 
    -22987.28, -23001.08, -23014.74, -23056.68, -23079.3, -23130.42, 
    -23121.12, -23136.9, -23152.12, -23178, -23173.71, -23185.22, -23136.48, 
    -23168.71, -23115.85, -23130.14, -23018.47, -22977.4, -22960.21, 
    -22945.29, -22909.54, -22934.15, -22924.4, -22947.68, -22962.63, 
    -22955.22, -23001.46, -22983.34, -23080.64, -23038.1, -23150.34, 
    -23123.03, -23156.95, -23139.55, -23169.49, -23142.52, -23189.53, 
    -23199.95, -23192.82, -23220.39, -23141.04, -23171.04, -22955.02, 
    -22956.22, -22961.85, -22937.23, -22935.74, -22913.49, -22933.27, 
    -22941.76, -22963.5, -22976.48, -22988.92, -23016.52, -23047.78, 
    -23092.47, -23124.79, -23146.78, -23133.26, -23145.19, -23131.86, 
    -23125.64, -23196.04, -23156.13, -23216.39, -23213, -23185.5, -23213.38, 
    -22957.07, -22950.13, -22926.27, -22944.92, -22911.09, -22929.94, 
    -22940.88, -22983.72, -22993.27, -23002.18, -23019.83, -23042.72, 
    -23083.65, -23119.64, -23153.01, -23150.54, -23151.41, -23158.96, 
    -23140.33, -23162.03, -23165.71, -23156.12, -23212.54, -23196.22, 
    -23212.92, -23202.27, -22952.38, -22964.08, -22957.75, -22969.67, 
    -22961.27, -22998.97, -23010.42, -23064.82, -23042.27, -23078.29, 
    -23045.89, -23051.59, -23079.48, -23047.63, -23117.65, -23070.01, 
    -23159.25, -23110.91, -23162.33, -23152.86, -23168.56, -23182.75, 
    -23200.79, -23234.62, -23226.72, -23255.44, -22981.66, -22997.11, 
    -22995.74, -23012.01, -23024.1, -23050.6, -23093.98, -23077.54, 
    -23107.63, -23113.67, -23068.01, -23096.09, -23007.52, -23021.52, 
    -23013.17, -22982.88, -23081.32, -23030.16, -23125.32, -23097.19, 
    -23180.72, -23138.64, -23222.39, -23259.6, -23295.41, -23337.94, 
    -23005.6, -22995.04, -23013.95, -23040.38, -23065.29, -23098.89, 
    -23102.31, -23108.6, -23124.98, -23138.89, -23110.59, -23142.4, 
    -23024.79, -23085.83, -22991.06, -23019.11, -23038.81, -23030.14, 
    -23075.68, -23086.58, -23131.02, -23107.97, -23250.34, -23185.77, 
    -23370.65, -23317.54, -22991.36, -23005.56, -23055.65, -23031.63, 
    -23101.12, -23118.39, -23132.56, -23150.86, -23152.85, -23163.81, 
    -23145.89, -23163.1, -23098.96, -23127.3, -23049.85, -23068.53, 
    -23059.91, -23050.5, -23079.68, -23111.03, -23111.7, -23121.79, -23150.6, 
    -23101.41, -23258.88, -23159.8, -23021.1, -23048.89, -23052.9, -23042.05, 
    -23116.65, -23089.48, -23163.54, -23143.21, -23176.65, -23159.95, 
    -23157.51, -23136.34, -23123.3, -23090.73, -23064.3, -23043.62, -23048.4, 
    -23071.21, -23112.95, -23153.03, -23144.17, -23174.09, -23096.07, 
    -23128.33, -23115.79, -23148.69, -23077.11, -23137.93, -23061.72, 
    -23068.34, -23088.94, -23130.54, -23139.86, -23149.88, -23143.69, 
    -23114.01, -23109.2, -23088.43, -23082.68, -23066.9, -23053.93, 
    -23065.78, -23078.29, -23114.02, -23146.63, -23182.96, -23191.97, 
    -23235.76, -23200.03, -23259.45, -23208.8, -23297.5, -23141.5, -23207.33, 
    -23089.88, -23102.22, -23124.59, -23177.11, -23148.54, -23182, -23109.01, 
    -23072, -23062.48, -23044.87, -23062.89, -23061.41, -23078.81, -23073.2, 
    -23115.21, -23092.68, -23157.45, -23181.73, -23252.4, -23297.32, 
    -23343.88, -23364.63, -23370.99, -23373.66 ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -1.679149e-14, -1.512313e-14, -1.570194e-14, -1.30169e-14, -1.375613e-14, 
    -1.676952e-14, -4.667439e-15, -1.041734e-14, -1.794265e-14, 
    -5.000467e-15, -1.114673e-14, -8.200681e-15, -1.917863e-14, 
    -1.536179e-14, -1.254234e-14, -1.918165e-14, -1.038964e-14, 
    -1.429787e-14, -1.542285e-14, -1.702438e-14, -5.229788e-15, 
    -1.055971e-14, -2.264654e-14, -8.881592e-15, -1.286745e-14, 
    -1.097316e-14, -1.376368e-14, -1.080667e-14, -1.273685e-14, 
    -8.353599e-15, -1.019064e-14, -1.343993e-14, -1.097886e-14, -1.12208e-14, 
    -1.554847e-14, -1.503838e-14, -1.597861e-14, -9.71335e-16, -2.209131e-15, 
    -1.350411e-14, -1.314523e-14, -1.072632e-14, -1.176109e-14, 
    -1.347109e-14, -6.030571e-15, -1.63121e-14, -1.333918e-14, -4.015277e-15, 
    -1.177409e-14, -1.716802e-14, -2.456201e-14, -1.128145e-14, 
    -1.363252e-14, -1.669326e-14, -5.708582e-15, -1.582731e-14, 
    -1.147882e-14, -1.380824e-14, -7.101675e-15, -2.358649e-14, 
    -1.043944e-14, -1.532288e-14, -1.797237e-14, -7.097895e-15, 
    -1.914224e-14, -1.346462e-14, -1.095813e-14, -2.411633e-14, 
    -1.301019e-14, -1.469757e-14, -1.561223e-14, -9.834689e-15, 
    -1.107121e-14, -8.543468e-15, -2.469282e-15, -1.74924e-14, -1.902458e-14, 
    -1.688924e-14, -8.402156e-15, -3.666899e-15, -1.592395e-14, 
    -1.997602e-14, -7.657771e-15, -1.136573e-14, -1.868986e-14, 
    -1.660133e-14, -1.257806e-14, -1.94658e-14, -1.078958e-14, -9.433651e-15, 
    -8.622258e-15, -1.385284e-14, -1.57277e-14, -1.446108e-14, -1.135725e-14, 
    -1.433309e-14, -1.245253e-14, -7.916366e-15, -1.615862e-14, 
    -1.491824e-14, -2.202424e-14, -1.942806e-14, -5.543745e-15, 
    -5.710568e-15, -1.278948e-14, -1.682998e-14, -1.638045e-14, -1.67352e-14, 
    -1.509105e-14, -1.664821e-14, -1.873423e-14, -1.565135e-14, 
    -1.579048e-14, -1.744741e-14, -1.880135e-14, -1.290754e-14, 
    -1.188672e-14, -8.961637e-15, -1.012136e-14, -1.1115e-14, -1.403707e-14, 
    -5.923478e-15, -1.724889e-14, -1.332661e-14, -1.668771e-14, 
    -9.254179e-15, -1.203664e-14, -8.326679e-15, -1.372904e-14, 
    -1.414031e-14, -1.535147e-14, -1.71694e-14, -1.370432e-14, -1.804217e-14, 
    -1.064633e-14, -5.370426e-15, -1.321267e-14, -1.315733e-14, 
    -1.404091e-14, -1.266755e-14, -1.526015e-14, -9.521131e-15, 
    -1.155903e-14, -9.480489e-15, -1.370843e-14, -5.99829e-15, -2.130532e-14, 
    -1.668777e-14, -8.605368e-15, -1.284111e-14, -1.875565e-14, 
    -1.364095e-14, -1.160295e-14, -9.275428e-15, -1.630892e-14, -8.27742e-15, 
    -1.763948e-14, -9.619065e-15, -1.656799e-16, -1.007854e-14, 
    -1.478542e-14, -5.410892e-15, -1.515335e-14, -1.511668e-14, -5.51176e-15, 
    -1.323109e-14, -1.896725e-14, -1.657101e-14, -6.991847e-15, 
    -1.884381e-14, -1.500221e-14, -1.563252e-14, -1.351499e-14, 
    -1.928904e-14, -5.609719e-15, -6.776522e-15, -2.446602e-15, 
    -1.374712e-14, -1.513088e-14, -1.346329e-14, -8.154452e-15, 
    -8.725317e-15, -1.158259e-14, -5.855388e-15, -1.561973e-14, 
    -1.898835e-14, -1.60644e-14, -9.991446e-15, -2.080875e-14, -1.905751e-14, 
    -1.163331e-14, -1.08516e-14, -7.155557e-15, -1.70222e-14, -1.443284e-14, 
    -1.449862e-14, -1.500535e-14, -1.695827e-14, -2.091054e-14, 
    -1.259649e-14, -9.416486e-15, -8.002509e-15, -9.867958e-15, 
    -8.500705e-15, -1.929022e-14, -7.980582e-15, -1.259321e-14, 
    -1.517272e-14, -1.711347e-14, -1.17136e-14, -9.997227e-15, -9.352282e-15, 
    -7.965474e-15, -6.44286e-15, -1.372282e-14, -1.431436e-14, -1.626112e-14, 
    -2.701224e-14, -1.039601e-14, -1.696808e-14, -1.878525e-14, 
    -1.416395e-14, -1.327291e-14, -7.897517e-15, 3.22583e-15, -1.076847e-14, 
    -1.238857e-14, -1.080477e-14, -7.20564e-15, -1.085466e-14, -9.388928e-15, 
    -1.358821e-14, -1.901994e-14, -1.268985e-14, -1.73024e-14, -1.169788e-14, 
    -1.796733e-14, -8.93127e-15, -8.046328e-15, -2.20216e-15, -6.756777e-15, 
    -1.051892e-14, -1.546484e-14, -5.665602e-15, -2.021421e-14, 
    -3.610932e-15, -1.761386e-15, 1.329122e-15, -1.133683e-14, -1.811706e-14, 
    -1.253524e-14, -1.845293e-14, -1.664673e-14, -1.151648e-14, 
    -1.629285e-14, -7.008494e-15, -2.1111e-14, -1.51735e-14, -1.575758e-14, 
    -2.424826e-14, -8.038741e-15, -4.175435e-15, -1.103964e-14, 
    -1.316633e-14, -1.273506e-14, -7.900929e-15, -1.207931e-14, 
    -1.235604e-14, -1.570425e-14, -1.025983e-14, -7.924739e-15, -2.71597e-14, 
    -4.48352e-15, -1.433737e-14, -1.362853e-14, -1.324306e-14, -1.773298e-14, 
    -1.024274e-14, -1.060815e-14, -1.5941e-14, -1.689181e-14, -1.216724e-14, 
    -9.500951e-15, -1.063934e-14, -1.607468e-14, -9.014562e-15, 
    -2.110638e-14, -1.00732e-14, -8.676653e-15, -1.716093e-14, -2.143712e-14, 
    -6.547892e-15, -1.648397e-14, -1.875596e-14, -1.388175e-14, 
    -1.084457e-14, -1.413552e-14, -7.843857e-15, -1.842909e-14, 
    -1.109723e-14, -1.422838e-14, -1.358882e-14, -1.222101e-14, 
    -1.258731e-14, -1.011394e-14, -1.46052e-14, -1.107221e-14, -1.265772e-14, 
    -1.431956e-14, -1.03401e-14, -2.240629e-14, -8.584313e-15, -8.685785e-15, 
    -1.94242e-14, -1.316562e-14, -1.178656e-14, -1.176421e-14, -1.851979e-14, 
    -2.142306e-14, -1.392568e-14, -2.601077e-14, -7.692838e-15, 
    -2.274409e-14, -7.878546e-15, -1.135702e-14, -7.510214e-15, 
    -1.844369e-14, -9.69561e-15, -2.065427e-14, -7.865608e-15, -1.870697e-14, 
    -1.831833e-14, -1.699152e-14, -4.518573e-15, -1.693727e-14, 
    -1.908026e-14, -1.010691e-14, -1.279921e-14 ;

 ERRSOI =
  -2.55794e-10, -3.872515e-10, -2.37985e-10, -4.882458e-10, -2.551985e-10, 
    -3.700595e-10, -2.860796e-10, -3.784759e-10, -2.296937e-10, 
    -4.980246e-10, -2.888184e-10, -4.051415e-10, -3.201044e-10, -3.64494e-10, 
    -2.411286e-10, -1.806006e-10, -3.882622e-10, -4.4857e-10, -4.34935e-10, 
    -1.649585e-10, -3.07225e-10, -4.800906e-10, -2.989412e-10, -3.098435e-10, 
    -6.714542e-10, -3.65532e-10, -3.546631e-10, -3.210593e-10, -4.234866e-10, 
    -4.217774e-10, -5.458975e-10, -2.780982e-10, -3.297003e-10, 
    -3.349148e-10, -3.472138e-10, -3.243898e-10, -2.788594e-10, 
    -2.138915e-10, -5.275601e-10, -3.825739e-10, -4.09106e-10, -3.577535e-10, 
    -3.379395e-10, -3.125125e-10, -2.348639e-10, -3.537506e-10, 
    -2.663126e-10, -3.139496e-10, -1.230342e-10, -3.51039e-10, -3.716767e-10, 
    -3.451943e-10, -4.011486e-10, -3.425655e-10, -4.549624e-10, 
    -3.357211e-10, -3.393028e-10, -1.74857e-10, -3.569237e-10, -3.291482e-10, 
    -3.568707e-10, -3.768742e-10, -2.303819e-10, -4.139493e-10, 
    -3.990697e-10, -4.542028e-10, -3.163996e-10, -3.397516e-10, 
    -4.619939e-10, -3.680898e-10, -4.332808e-10, -3.648435e-10, -2.50212e-10, 
    -3.616189e-10, -5.045985e-10, -3.193966e-10, -4.166982e-10, 
    -3.125541e-10, -3.747784e-10, -4.420379e-10, -2.788123e-10, 
    -4.018803e-10, -2.044054e-10, -3.372795e-10, -4.350432e-10, 
    -1.833512e-10, -2.8212e-10, -5.232875e-10, -4.124328e-10, -3.144127e-10, 
    -4.147474e-10, -4.901408e-10, -4.086207e-10, -4.447513e-10, 
    -2.536997e-10, -3.308468e-10, -3.173776e-10, -2.108933e-10, 
    -4.872056e-10, -2.497974e-10, -2.961421e-10, -4.92312e-10, -3.582837e-10, 
    -2.818402e-10, -4.38655e-10, -3.983656e-10, -2.313541e-10, -4.709537e-10, 
    -2.996736e-10, -2.689384e-10, -4.108727e-10, -6.230886e-10, -3.37462e-10, 
    -4.885416e-10, -3.881741e-10, -5.311789e-10, -4.134232e-10, 
    -4.024692e-10, -1.817821e-10, -3.943284e-10, -2.933275e-10, 
    -4.494596e-10, -5.23777e-10, -4.116235e-10, -4.576773e-10, -3.260541e-10, 
    -4.790318e-10, -5.273171e-10, -6.252497e-10, -3.325229e-10, 
    -1.386551e-10, -4.748222e-10, -3.808207e-10, -4.719433e-10, 
    -3.654267e-10, -5.364849e-10, -5.351049e-10, -3.203562e-10, 
    -3.570607e-10, -4.419924e-10, -3.202227e-10, -3.304013e-10, 
    -4.324669e-10, -5.260332e-10, -3.120607e-10, -4.569912e-10, 
    -3.547005e-10, -3.545807e-10, -3.171738e-10, -5.137306e-10, 
    -3.087456e-10, -4.189064e-10, -3.544425e-10, -4.25429e-10, -2.844097e-10, 
    -2.654752e-10, -1.102529e-10, -3.279e-10, -2.19299e-10, -3.495582e-10, 
    -3.794819e-10, -4.128478e-10, -2.754864e-10, -4.939071e-10, 
    -5.916117e-10, -5.527282e-10, -3.114363e-10, -4.619502e-10, 
    -1.961977e-10, -5.881349e-10, -3.874997e-10, -3.738936e-10, 
    -3.496516e-10, -3.404358e-10, -2.352859e-10, -3.307715e-10, 
    -3.017642e-10, -3.263664e-10, -3.23256e-10, -4.909149e-10, -6.297231e-10, 
    -4.48544e-10, -3.81973e-10, -3.704245e-10, -4.336906e-10, -3.949806e-10, 
    -4.878264e-10, -4.197453e-10, -3.434458e-10, -3.936471e-10, 
    -3.616519e-10, -2.368557e-10, -3.939072e-10, -3.241001e-10, 
    -3.568738e-10, -1.872979e-10, -4.066921e-10, -4.664683e-10, 
    -3.044306e-10, -5.415154e-10, -1.647437e-10, -4.076154e-10, 
    -3.345396e-10, -3.350476e-10, -2.665697e-10, -2.944124e-10, 
    -3.720061e-10, -9.702626e-11, -2.574704e-10, -1.999101e-10, 
    -3.754403e-10, -4.151927e-10, -3.774618e-10, -4.084128e-10, 
    -4.314679e-10, -5.285207e-10, -3.029004e-10, -2.156447e-10, 
    -3.250044e-10, -3.359008e-10, -3.149883e-10, -6.0139e-10, -4.218026e-10, 
    -1.229783e-10, -3.718808e-10, -4.012415e-10, -3.311218e-10, 
    -4.296056e-10, -2.357873e-10, -4.094882e-10, -1.874222e-10, 
    -3.643226e-10, -3.496844e-10, -2.287769e-10, -4.019188e-10, 
    -5.538466e-10, -3.925097e-10, -4.055668e-10, -3.571948e-10, 
    -4.687146e-10, -2.405624e-10, -3.662522e-10, -3.4035e-10, -3.05694e-10, 
    -4.956612e-10, -2.435898e-10, -4.065887e-10, -3.287504e-10, 
    -3.921643e-10, -1.300362e-10, -4.008781e-10, -5.079189e-10, 
    -2.721173e-10, -2.757715e-10, -3.922159e-10, -3.656921e-10, 
    -5.456062e-10, -3.327493e-10, -2.96679e-10, -3.097302e-10, -4.501604e-10, 
    -5.871115e-10, -5.696658e-10, -4.436278e-10, -4.116573e-10, 
    -3.213528e-10, -3.542123e-10, -1.90547e-10, -2.058452e-10, -2.947567e-10, 
    -3.504112e-10, -3.556554e-10, -2.858954e-10, -3.249253e-10, 
    -3.483523e-10, -3.393494e-10, -4.085698e-10, -3.631264e-10, -4.53994e-10, 
    -2.312421e-10, -5.02995e-10, -2.608443e-10, -2.886423e-10, -3.14417e-10, 
    -2.911621e-10, -2.217975e-10, -4.49298e-10, -3.223572e-10, -3.566987e-10, 
    -4.007628e-10, -5.429732e-10, -2.088541e-10, -4.080998e-10, 
    -3.269929e-10, -5.189577e-10, -3.62624e-10, -4.195168e-10, -3.655721e-10, 
    -4.077992e-10, -2.502028e-10, -3.45798e-10, -3.744954e-10, -3.763097e-10, 
    -4.294994e-10, -5.792561e-10, -4.634256e-10, -3.396314e-10, 
    -2.995005e-10, -1.775338e-10, -3.553186e-10, -5.129904e-10, 
    -3.634137e-10, -3.345064e-10, -2.860818e-10, -4.158165e-10, 
    -3.388813e-10, -3.697278e-10, -3.744479e-10, -3.821206e-10, -3.8303e-10, 
    -2.863613e-10, -4.160548e-10, -3.496754e-10, -4.094401e-10, 
    -5.008222e-10, -2.301304e-10, -4.15862e-10, -3.629379e-10, -5.354867e-10, 
    -3.872639e-10, -5.411662e-10, -4.095855e-10, -2.671027e-10, 
    -2.495106e-10, -3.521864e-10, -2.042493e-10, -2.420156e-10, -2.456282e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  1.77948e-16, 1.72803e-16, 1.738034e-16, 1.696532e-16, 1.719556e-16, 
    1.692379e-16, 1.769052e-16, 1.725985e-16, 1.75348e-16, 1.774852e-16, 
    1.615979e-16, 1.694681e-16, 1.534244e-16, 1.584442e-16, 1.45834e-16, 
    1.542052e-16, 1.441459e-16, 1.460762e-16, 1.402678e-16, 1.419319e-16, 
    1.344998e-16, 1.394997e-16, 1.306474e-16, 1.356943e-16, 1.349046e-16, 
    1.396645e-16, 1.67885e-16, 1.625775e-16, 1.681992e-16, 1.674425e-16, 
    1.677822e-16, 1.719078e-16, 1.739864e-16, 1.783416e-16, 1.775511e-16, 
    1.743526e-16, 1.671022e-16, 1.695638e-16, 1.633611e-16, 1.635011e-16, 
    1.565945e-16, 1.597087e-16, 1.480991e-16, 1.513993e-16, 1.418625e-16, 
    1.44261e-16, 1.41975e-16, 1.426683e-16, 1.41966e-16, 1.454837e-16, 
    1.439766e-16, 1.47072e-16, 1.591253e-16, 1.555831e-16, 1.661467e-16, 
    1.724969e-16, 1.767162e-16, 1.797097e-16, 1.792865e-16, 1.784796e-16, 
    1.743338e-16, 1.704365e-16, 1.674662e-16, 1.654791e-16, 1.635213e-16, 
    1.57593e-16, 1.544564e-16, 1.474314e-16, 1.486999e-16, 1.465515e-16, 
    1.444997e-16, 1.410538e-16, 1.416211e-16, 1.401027e-16, 1.466086e-16, 
    1.422847e-16, 1.494223e-16, 1.474702e-16, 1.629867e-16, 1.688999e-16, 
    1.714111e-16, 1.73611e-16, 1.789611e-16, 1.752663e-16, 1.767228e-16, 
    1.732582e-16, 1.710564e-16, 1.721455e-16, 1.654248e-16, 1.680376e-16, 
    1.542705e-16, 1.602009e-16, 1.44739e-16, 1.484396e-16, 1.43852e-16, 
    1.461932e-16, 1.421815e-16, 1.45792e-16, 1.395378e-16, 1.381755e-16, 
    1.391064e-16, 1.35531e-16, 1.459921e-16, 1.419748e-16, 1.721759e-16, 
    1.719983e-16, 1.71171e-16, 1.748075e-16, 1.750301e-16, 1.783632e-16, 
    1.753976e-16, 1.741345e-16, 1.70929e-16, 1.690325e-16, 1.672298e-16, 
    1.632661e-16, 1.588387e-16, 1.526477e-16, 1.481997e-16, 1.452177e-16, 
    1.470464e-16, 1.454319e-16, 1.472366e-16, 1.480826e-16, 1.386858e-16, 
    1.439624e-16, 1.360453e-16, 1.364835e-16, 1.400665e-16, 1.364341e-16, 
    1.718736e-16, 1.728957e-16, 1.764437e-16, 1.736671e-16, 1.787262e-16, 
    1.758941e-16, 1.742654e-16, 1.679825e-16, 1.666025e-16, 1.653223e-16, 
    1.627942e-16, 1.595493e-16, 1.538563e-16, 1.489027e-16, 1.443804e-16, 
    1.447118e-16, 1.445951e-16, 1.435846e-16, 1.460874e-16, 1.431736e-16, 
    1.426844e-16, 1.439633e-16, 1.365422e-16, 1.386626e-16, 1.364928e-16, 
    1.378735e-16, 1.725635e-16, 1.708437e-16, 1.71773e-16, 1.700255e-16, 
    1.712564e-16, 1.65782e-16, 1.641406e-16, 1.564603e-16, 1.59613e-16, 
    1.545959e-16, 1.591036e-16, 1.583047e-16, 1.544313e-16, 1.588601e-16, 
    1.491754e-16, 1.557407e-16, 1.435453e-16, 1.501015e-16, 1.431343e-16, 
    1.444e-16, 1.423047e-16, 1.404277e-16, 1.380667e-16, 1.337089e-16, 
    1.347182e-16, 1.310737e-16, 1.682801e-16, 1.660492e-16, 1.66246e-16, 
    1.639116e-16, 1.621851e-16, 1.584432e-16, 1.524406e-16, 1.546981e-16, 
    1.505541e-16, 1.49722e-16, 1.560179e-16, 1.52152e-16, 1.645565e-16, 
    1.625521e-16, 1.637458e-16, 1.681039e-16, 1.541773e-16, 1.613246e-16, 
    1.481261e-16, 1.519988e-16, 1.406953e-16, 1.463168e-16, 1.352736e-16, 
    1.305501e-16, 1.261058e-16, 1.209084e-16, 1.648321e-16, 1.663479e-16, 
    1.636342e-16, 1.598785e-16, 1.563949e-16, 1.517625e-16, 1.512888e-16, 
    1.504207e-16, 1.481727e-16, 1.462823e-16, 1.501459e-16, 1.458085e-16, 
    1.620864e-16, 1.53557e-16, 1.669206e-16, 1.628963e-16, 1.601001e-16, 
    1.613272e-16, 1.549562e-16, 1.534543e-16, 1.473506e-16, 1.505063e-16, 
    1.317157e-16, 1.400306e-16, 1.169516e-16, 1.234034e-16, 1.668774e-16, 
    1.648375e-16, 1.577368e-16, 1.611155e-16, 1.514535e-16, 1.490747e-16, 
    1.471411e-16, 1.446686e-16, 1.44402e-16, 1.429369e-16, 1.453375e-16, 
    1.430319e-16, 1.517527e-16, 1.478559e-16, 1.58549e-16, 1.559464e-16, 
    1.571438e-16, 1.58457e-16, 1.54404e-16, 1.500849e-16, 1.499933e-16, 
    1.486082e-16, 1.447034e-16, 1.514144e-16, 1.306409e-16, 1.434707e-16, 
    1.62613e-16, 1.586825e-16, 1.58122e-16, 1.596444e-16, 1.493131e-16, 
    1.530567e-16, 1.429728e-16, 1.456985e-16, 1.412324e-16, 1.434518e-16, 
    1.437782e-16, 1.466285e-16, 1.484027e-16, 1.52885e-16, 1.565317e-16, 
    1.594237e-16, 1.587513e-16, 1.555745e-16, 1.498209e-16, 1.443775e-16, 
    1.455699e-16, 1.415719e-16, 1.521541e-16, 1.477168e-16, 1.494317e-16, 
    1.449602e-16, 1.547579e-16, 1.464126e-16, 1.568905e-16, 1.559721e-16, 
    1.53131e-16, 1.474154e-16, 1.461517e-16, 1.448012e-16, 1.456347e-16, 
    1.496749e-16, 1.503371e-16, 1.532003e-16, 1.539904e-16, 1.561721e-16, 
    1.579779e-16, 1.563278e-16, 1.545947e-16, 1.496735e-16, 1.452376e-16, 
    1.404009e-16, 1.392174e-16, 1.33563e-16, 1.38165e-16, 1.305693e-16, 
    1.370258e-16, 1.258488e-16, 1.459301e-16, 1.372171e-16, 1.53002e-16, 
    1.51302e-16, 1.482262e-16, 1.41172e-16, 1.449813e-16, 1.405267e-16, 
    1.503631e-16, 1.554646e-16, 1.567852e-16, 1.592478e-16, 1.567289e-16, 
    1.569338e-16, 1.545235e-16, 1.552981e-16, 1.495101e-16, 1.526193e-16, 
    1.437862e-16, 1.40562e-16, 1.314555e-16, 1.258706e-16, 1.201853e-16, 
    1.176744e-16, 1.169102e-16, 1.165906e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  22.1825, 22.24694, 22.23443, 22.28639, 22.25759, 22.2916, 22.1956, 
    22.24946, 22.21509, 22.18835, 22.3872, 22.28872, 22.49, 22.42704, 
    22.58541, 22.48015, 22.60666, 22.58246, 22.65555, 22.63461, 22.72797, 
    22.66522, 22.77655, 22.71303, 22.72293, 22.66313, 22.30861, 22.37491, 
    22.30466, 22.31412, 22.3099, 22.25816, 22.23204, 22.17764, 22.18753, 
    22.22752, 22.31837, 22.28758, 22.36539, 22.36363, 22.45027, 22.4112, 
    22.55702, 22.51557, 22.63549, 22.6053, 22.63405, 22.62534, 22.63416, 
    22.5899, 22.60886, 22.56995, 22.4185, 22.46295, 22.33039, 22.25064, 
    22.19794, 22.16051, 22.1658, 22.17587, 22.22775, 22.27664, 22.31389, 
    22.33881, 22.36337, 22.43756, 22.47704, 22.56536, 22.54949, 22.57644, 
    22.6023, 22.64563, 22.63851, 22.65759, 22.57579, 22.63011, 22.54044, 
    22.56495, 22.36975, 22.2959, 22.26427, 22.23682, 22.16986, 22.21608, 
    22.19785, 22.24129, 22.26887, 22.25524, 22.33949, 22.30671, 22.47938, 
    22.40496, 22.59929, 22.55276, 22.61045, 22.58102, 22.63143, 22.58606, 
    22.66471, 22.68181, 22.67012, 22.71515, 22.58354, 22.63402, 22.25484, 
    22.25706, 22.26744, 22.22182, 22.21904, 22.17735, 22.21447, 22.23027, 
    22.27049, 22.29423, 22.31683, 22.36654, 22.42205, 22.49981, 22.55577, 
    22.59329, 22.5703, 22.59059, 22.5679, 22.55728, 22.67538, 22.60902, 
    22.70867, 22.70316, 22.65803, 22.70378, 22.25863, 22.24584, 22.20136, 
    22.23617, 22.17282, 22.20823, 22.22858, 22.30733, 22.32472, 22.34075, 
    22.37248, 22.41319, 22.48464, 22.5469, 22.60382, 22.59965, 22.60112, 
    22.61381, 22.58234, 22.61897, 22.6251, 22.60905, 22.70242, 22.67574, 
    22.70304, 22.68568, 22.25, 22.27154, 22.2599, 22.28177, 22.26633, 
    22.33491, 22.35547, 22.45188, 22.41237, 22.47533, 22.41879, 22.42879, 
    22.47726, 22.42187, 22.54341, 22.46087, 22.6143, 22.53169, 22.61947, 
    22.60357, 22.62993, 22.65351, 22.68323, 22.73802, 22.72534, 22.77123, 
    22.30367, 22.3316, 22.32919, 22.35846, 22.3801, 22.4271, 22.50245, 
    22.47412, 22.5262, 22.53664, 22.45756, 22.50605, 22.35033, 22.37541, 
    22.36052, 22.30584, 22.48057, 22.39082, 22.55668, 22.50802, 22.65014, 
    22.57937, 22.71835, 22.77768, 22.83382, 22.89915, 22.3469, 22.32792, 
    22.36196, 22.40898, 22.45279, 22.51098, 22.51696, 22.52785, 22.55614, 
    22.5799, 22.53124, 22.58586, 22.38111, 22.4884, 22.32069, 22.37108, 
    22.40623, 22.39087, 22.4709, 22.48976, 22.5664, 22.5268, 22.76298, 
    22.65841, 22.94911, 22.86775, 22.32127, 22.34686, 22.4359, 22.39353, 
    22.51489, 22.54477, 22.56911, 22.60014, 22.60354, 22.62194, 22.59178, 
    22.62077, 22.5111, 22.5601, 22.42578, 22.45842, 22.44343, 22.42694, 
    22.47783, 22.53199, 22.53324, 22.5506, 22.59937, 22.51539, 22.77631, 
    22.61492, 22.37477, 22.42397, 22.43111, 22.41203, 22.54177, 22.49472, 
    22.6215, 22.58724, 22.64341, 22.61548, 22.61137, 22.57554, 22.55322, 
    22.49686, 22.45106, 22.41481, 22.42324, 22.46307, 22.53533, 22.6038, 
    22.58879, 22.63914, 22.50608, 22.5618, 22.54023, 22.59651, 22.47335, 
    22.57793, 22.44661, 22.45813, 22.49379, 22.56552, 22.58154, 22.59847, 
    22.58804, 22.53718, 22.52889, 22.49295, 22.48298, 22.45563, 22.43295, 
    22.45365, 22.47537, 22.53724, 22.59298, 22.65383, 22.66876, 22.73968, 
    22.68182, 22.77719, 22.69591, 22.83676, 22.58413, 22.6937, 22.49545, 
    22.5168, 22.55535, 22.64403, 22.59624, 22.65218, 22.52857, 22.4644, 
    22.44792, 22.41699, 22.44863, 22.44606, 22.47634, 22.46661, 22.5393, 
    22.50025, 22.61124, 22.65176, 22.76638, 22.83666, 22.90841, 22.94004, 
    22.94968, 22.95371 ;

 FGR =
  -389.0773, -390.1737, -389.9607, -390.8445, -390.3545, -390.933, -389.2999, 
    -390.2169, -389.6317, -389.1764, -392.5582, -390.884, -394.299, 
    -393.2315, -395.9133, -394.1325, -396.2723, -395.8625, -397.0972, 
    -396.7436, -398.3208, -397.2604, -399.1391, -398.068, -398.2353, 
    -397.2253, -391.2216, -392.3496, -391.1546, -391.3155, -391.2434, 
    -390.3644, -389.9209, -388.994, -389.1624, -389.8434, -391.3879, 
    -390.8641, -392.1852, -392.1554, -393.6252, -392.9626, -395.4324, 
    -394.7308, -396.7584, -396.2485, -396.7343, -396.5871, -396.7362, 
    -395.9885, -396.3088, -395.6509, -393.0866, -393.8402, -391.5916, 
    -390.2379, -389.34, -388.7023, -388.7924, -388.9642, -389.8474, 
    -390.6782, -391.311, -391.7342, -392.1512, -393.4113, -394.0795, 
    -395.574, -395.3049, -395.7612, -396.1978, -396.93, -396.8096, -397.132, 
    -395.7495, -396.6682, -395.1514, -395.5663, -392.2623, -391.0055, 
    -390.4693, -390.0016, -388.8617, -389.6488, -389.3385, -390.0771, 
    -390.5461, -390.3142, -391.7457, -391.1892, -394.119, -392.8574, 
    -396.1469, -395.3601, -396.3355, -395.838, -396.6902, -395.9232, 
    -397.2521, -397.5411, -397.3436, -398.1031, -395.8806, -396.7341, 
    -390.3076, -390.3455, -390.5218, -389.7465, -389.6992, -388.9892, 
    -389.6212, -389.89, -390.5735, -390.9772, -391.3612, -392.2052, 
    -393.1472, -394.4647, -395.4111, -396.0453, -395.6566, -395.9998, 
    -395.6161, -395.4363, -397.4327, -396.3117, -397.9939, -397.9009, 
    -397.1395, -397.9114, -390.372, -390.1544, -389.3982, -389.99, -388.9119, 
    -389.5152, -389.8618, -391.2003, -391.4949, -391.7673, -392.3058, 
    -392.9965, -394.2076, -395.2614, -396.2233, -396.1529, -396.1776, 
    -396.3923, -395.8603, -396.4796, -396.5833, -396.3118, -397.8885, 
    -397.4381, -397.8989, -397.6058, -390.2252, -390.5915, -390.3935, 
    -390.7656, -390.5033, -391.6688, -392.0182, -393.6531, -392.9828, 
    -394.0502, -393.0914, -393.2612, -394.084, -393.1434, -395.2029, 
    -393.8059, -396.4006, -395.0053, -396.488, -396.2191, -396.6645, 
    -397.063, -397.5647, -398.4895, -398.2755, -399.049, -391.1376, 
    -391.6123, -391.5709, -392.0679, -392.4353, -393.2321, -394.509, 
    -394.029, -394.9106, -395.0874, -393.7483, -394.5702, -391.9302, 
    -392.3565, -392.103, -391.1748, -394.1391, -392.6179, -395.4267, 
    -394.6031, -397.0061, -395.8109, -398.1575, -399.159, -400.103, 
    -401.2035, -391.8718, -391.5492, -392.1271, -392.9258, -393.6678, 
    -394.6533, -394.7543, -394.9388, -395.4171, -395.8189, -394.9967, 
    -395.9197, -392.4545, -394.2713, -391.4269, -392.2831, -392.8789, 
    -392.618, -393.9743, -394.2937, -395.5913, -394.9208, -398.9115, 
    -397.1466, -402.0424, -400.675, -391.4364, -391.8708, -393.3819, 
    -392.6631, -394.7193, -395.225, -395.6365, -396.1616, -396.2186, 
    -396.5298, -396.0198, -396.5098, -394.6554, -395.4843, -393.2097, 
    -393.7632, -393.5087, -393.2292, -394.0917, -395.0096, -395.0298, 
    -395.324, -396.1516, -394.7276, -399.1379, -396.4139, -392.3445, 
    -393.1801, -393.3003, -392.9765, -395.1743, -394.3781, -396.5223, 
    -395.9431, -396.8922, -396.4206, -396.3511, -395.7454, -395.368, 
    -394.4144, -393.6386, -393.0235, -393.1666, -393.8422, -395.0659, 
    -396.2235, -395.9698, -396.8201, -394.5702, -395.5135, -395.1487, 
    -396.0999, -394.0161, -395.7887, -393.5627, -393.758, -394.3622, 
    -395.577, -395.8467, -396.1334, -395.9567, -395.097, -394.9565, 
    -394.3477, -394.1793, -393.7155, -393.3312, -393.6822, -394.0506, 
    -395.0977, -396.0406, -397.0685, -397.3203, -398.519, -397.5424, 
    -399.153, -397.7823, -400.1552, -395.8923, -397.7433, -394.39, -394.7516, 
    -395.4048, -396.9039, -396.0954, -397.0413, -394.951, -393.8652, 
    -393.585, -393.0608, -393.597, -393.5534, -394.0663, -393.9016, 
    -395.1324, -394.4713, -396.3492, -397.034, -398.9677, -400.1519, 
    -401.3578, -401.8897, -402.0516, -402.1192 ;

 FGR12 =
  -50.36827, -50.43694, -50.42362, -50.47903, -50.44832, -50.4846, -50.38223, 
    -50.43963, -50.403, -50.3745, -50.58674, -50.48154, -50.69683, -50.6294, 
    -50.79919, -50.68629, -50.82204, -50.79605, -50.8746, -50.85209, 
    -50.95255, -50.88501, -51.0049, -50.93647, -50.94711, -50.88276, 
    -50.50278, -50.57359, -50.49856, -50.50865, -50.50414, -50.44892, 
    -50.42105, -50.36309, -50.37363, -50.41624, -50.5132, -50.48032, 
    -50.56344, -50.56157, -50.65427, -50.61245, -50.76873, -50.72427, 
    -50.85302, -50.82058, -50.85149, -50.84212, -50.8516, -50.80405, 
    -50.8244, -50.78262, -50.62025, -50.66784, -50.52602, -50.4409, 
    -50.38472, -50.34484, -50.35048, -50.3612, -50.41649, -50.46864, 
    -50.50842, -50.53503, -50.5613, -50.64064, -50.68295, -50.77768, 
    -50.76066, -50.78958, -50.81736, -50.86393, -50.85628, -50.87679, 
    -50.78889, -50.84724, -50.75094, -50.77724, -50.56808, -50.4892, 
    -50.45543, -50.42616, -50.35481, -50.40404, -50.38462, -50.43092, 
    -50.46035, -50.44581, -50.53576, -50.50075, -50.68544, -50.60578, 
    -50.81411, -50.76416, -50.82611, -50.79451, -50.84866, -50.79992, 
    -50.88446, -50.90285, -50.89028, -50.93874, -50.79721, -50.85145, 
    -50.44539, -50.44775, -50.45882, -50.41017, -50.4072, -50.36279, 
    -50.40234, -50.41917, -50.46208, -50.48742, -50.51156, -50.56467, 
    -50.62406, -50.70735, -50.76739, -50.80767, -50.78299, -50.80478, 
    -50.78041, -50.76901, -50.89593, -50.82458, -50.93177, -50.92584, 
    -50.87727, -50.9265, -50.44942, -50.43579, -50.38837, -50.42547, 
    -50.35796, -50.39568, -50.41739, -50.5014, -50.51998, -50.5371, 
    -50.57103, -50.61457, -50.6911, -50.75786, -50.81899, -50.81451, 
    -50.81609, -50.82972, -50.79592, -50.83527, -50.84185, -50.82461, 
    -50.92504, -50.89632, -50.92571, -50.90702, -50.44023, -50.4632, 
    -50.45078, -50.47411, -50.45765, -50.53085, -50.55285, -50.65598, 
    -50.6137, -50.68111, -50.62057, -50.63127, -50.68317, -50.62386, 
    -50.75411, -50.66563, -50.83024, -50.74155, -50.83581, -50.81873, 
    -50.84705, -50.8724, -50.90439, -50.96338, -50.94973, -50.99918, 
    -50.49751, -50.52732, -50.52476, -50.55603, -50.57918, -50.62946, 
    -50.71019, -50.67983, -50.73566, -50.74686, -50.66208, -50.71404, 
    -50.54735, -50.57415, -50.55824, -50.49983, -50.68673, -50.59064, 
    -50.76837, -50.71616, -50.86877, -50.79273, -50.9422, -51.00613, 
    -51.06661, -51.13707, -50.54367, -50.5234, -50.55978, -50.61006, 
    -50.65697, -50.71932, -50.72575, -50.73743, -50.76778, -50.79329, 
    -50.74107, -50.79969, -50.58026, -50.69511, -50.51568, -50.56952, 
    -50.60712, -50.59069, -50.67638, -50.69658, -50.7788, -50.73631, 
    -50.99028, -50.87767, -51.19102, -51.10319, -50.5163, -50.54364, 
    -50.63888, -50.59354, -50.72353, -50.75558, -50.78171, -50.81504, 
    -50.81869, -50.83846, -50.80606, -50.8372, -50.71947, -50.77203, 
    -50.62806, -50.663, -50.64694, -50.62929, -50.68381, -50.74186, 
    -50.74322, -50.76184, -50.81419, -50.72408, -51.00464, -50.83092, 
    -50.57348, -50.6261, -50.63375, -50.61333, -50.75236, -50.70191, 
    -50.83799, -50.80118, -50.86154, -50.83153, -50.8271, -50.78862, 
    -50.76465, -50.7042, -50.65512, -50.61631, -50.62534, -50.66798, 
    -50.74545, -50.81896, -50.80284, -50.85695, -50.7141, -50.77387, 
    -50.75072, -50.81113, -50.67901, -50.79116, -50.65036, -50.6627, 
    -50.70091, -50.77784, -50.79506, -50.81324, -50.80204, -50.74744, 
    -50.73854, -50.7, -50.68931, -50.66002, -50.63573, -50.65789, -50.68117, 
    -50.7475, -50.80735, -50.87274, -50.88882, -50.96516, -50.90287, 
    -51.0056, -50.91803, -51.06977, -50.79785, -50.91564, -50.70269, 
    -50.72558, -50.76694, -50.86219, -50.81085, -50.87096, -50.7382, 
    -50.66941, -50.65176, -50.61865, -50.65252, -50.64977, -50.6822, 
    -50.67178, -50.74971, -50.70784, -50.82697, -50.87052, -50.99396, 
    -51.06967, -51.14706, -51.18123, -51.19165, -51.196 ;

 FGR_R =
  -389.0773, -390.1737, -389.9607, -390.8445, -390.3545, -390.933, -389.2999, 
    -390.2169, -389.6317, -389.1764, -392.5582, -390.884, -394.299, 
    -393.2315, -395.9133, -394.1325, -396.2723, -395.8625, -397.0972, 
    -396.7436, -398.3208, -397.2604, -399.1391, -398.068, -398.2353, 
    -397.2253, -391.2216, -392.3496, -391.1546, -391.3155, -391.2434, 
    -390.3644, -389.9209, -388.994, -389.1624, -389.8434, -391.3879, 
    -390.8641, -392.1852, -392.1554, -393.6252, -392.9626, -395.4324, 
    -394.7308, -396.7584, -396.2485, -396.7343, -396.5871, -396.7362, 
    -395.9885, -396.3088, -395.6509, -393.0866, -393.8402, -391.5916, 
    -390.2379, -389.34, -388.7023, -388.7924, -388.9642, -389.8474, 
    -390.6782, -391.311, -391.7342, -392.1512, -393.4113, -394.0795, 
    -395.574, -395.3049, -395.7612, -396.1978, -396.93, -396.8096, -397.132, 
    -395.7495, -396.6682, -395.1514, -395.5663, -392.2623, -391.0055, 
    -390.4693, -390.0016, -388.8617, -389.6488, -389.3385, -390.0771, 
    -390.5461, -390.3142, -391.7457, -391.1892, -394.119, -392.8574, 
    -396.1469, -395.3601, -396.3355, -395.838, -396.6902, -395.9232, 
    -397.2521, -397.5411, -397.3436, -398.1031, -395.8806, -396.7341, 
    -390.3076, -390.3455, -390.5218, -389.7465, -389.6992, -388.9892, 
    -389.6212, -389.89, -390.5735, -390.9772, -391.3612, -392.2052, 
    -393.1472, -394.4647, -395.4111, -396.0453, -395.6566, -395.9998, 
    -395.6161, -395.4363, -397.4327, -396.3117, -397.9939, -397.9009, 
    -397.1395, -397.9114, -390.372, -390.1544, -389.3982, -389.99, -388.9119, 
    -389.5152, -389.8618, -391.2003, -391.4949, -391.7673, -392.3058, 
    -392.9965, -394.2076, -395.2614, -396.2233, -396.1529, -396.1776, 
    -396.3923, -395.8603, -396.4796, -396.5833, -396.3118, -397.8885, 
    -397.4381, -397.8989, -397.6058, -390.2252, -390.5915, -390.3935, 
    -390.7656, -390.5033, -391.6688, -392.0182, -393.6531, -392.9828, 
    -394.0502, -393.0914, -393.2612, -394.084, -393.1434, -395.2029, 
    -393.8059, -396.4006, -395.0053, -396.488, -396.2191, -396.6645, 
    -397.063, -397.5647, -398.4895, -398.2755, -399.049, -391.1376, 
    -391.6123, -391.5709, -392.0679, -392.4353, -393.2321, -394.509, 
    -394.029, -394.9106, -395.0874, -393.7483, -394.5702, -391.9302, 
    -392.3565, -392.103, -391.1748, -394.1391, -392.6179, -395.4267, 
    -394.6031, -397.0061, -395.8109, -398.1575, -399.159, -400.103, 
    -401.2035, -391.8718, -391.5492, -392.1271, -392.9258, -393.6678, 
    -394.6533, -394.7543, -394.9388, -395.4171, -395.8189, -394.9967, 
    -395.9197, -392.4545, -394.2713, -391.4269, -392.2831, -392.8789, 
    -392.618, -393.9743, -394.2937, -395.5913, -394.9208, -398.9115, 
    -397.1466, -402.0424, -400.675, -391.4364, -391.8708, -393.3819, 
    -392.6631, -394.7193, -395.225, -395.6365, -396.1616, -396.2186, 
    -396.5298, -396.0198, -396.5098, -394.6554, -395.4843, -393.2097, 
    -393.7632, -393.5087, -393.2292, -394.0917, -395.0096, -395.0298, 
    -395.324, -396.1516, -394.7276, -399.1379, -396.4139, -392.3445, 
    -393.1801, -393.3003, -392.9765, -395.1743, -394.3781, -396.5223, 
    -395.9431, -396.8922, -396.4206, -396.3511, -395.7454, -395.368, 
    -394.4144, -393.6386, -393.0235, -393.1666, -393.8422, -395.0659, 
    -396.2235, -395.9698, -396.8201, -394.5702, -395.5135, -395.1487, 
    -396.0999, -394.0161, -395.7887, -393.5627, -393.758, -394.3622, 
    -395.577, -395.8467, -396.1334, -395.9567, -395.097, -394.9565, 
    -394.3477, -394.1793, -393.7155, -393.3312, -393.6822, -394.0506, 
    -395.0977, -396.0406, -397.0685, -397.3203, -398.519, -397.5424, 
    -399.153, -397.7823, -400.1552, -395.8923, -397.7433, -394.39, -394.7516, 
    -395.4048, -396.9039, -396.0954, -397.0413, -394.951, -393.8652, 
    -393.585, -393.0608, -393.597, -393.5534, -394.0663, -393.9016, 
    -395.1324, -394.4713, -396.3492, -397.034, -398.9677, -400.1519, 
    -401.3578, -401.8897, -402.0516, -402.1192 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  46.42476, 46.50126, 46.4864, 46.54806, 46.51388, 46.55423, 46.4403, 
    46.50428, 46.46345, 46.43168, 46.6676, 46.55082, 46.78905, 46.71459, 
    46.90166, 46.77744, 46.92671, 46.89813, 46.98426, 46.95959, 47.0696, 
    46.99564, 47.12669, 47.05197, 47.06364, 46.99319, 46.57437, 46.65305, 
    46.5697, 46.58092, 46.5759, 46.51457, 46.48362, 46.41895, 46.4307, 
    46.47822, 46.58597, 46.54943, 46.6416, 46.63952, 46.74205, 46.69583, 
    46.86813, 46.81918, 46.96062, 46.92506, 46.95894, 46.94867, 46.95908, 
    46.90691, 46.92926, 46.88337, 46.70448, 46.75705, 46.60018, 46.50573, 
    46.4431, 46.3986, 46.40489, 46.41687, 46.4785, 46.53646, 46.58061, 
    46.61013, 46.63922, 46.72712, 46.77374, 46.878, 46.85923, 46.89106, 
    46.92152, 46.97259, 46.96419, 46.98668, 46.89025, 46.95433, 46.84853, 
    46.87746, 46.64696, 46.5593, 46.52188, 46.48925, 46.40972, 46.46464, 
    46.44299, 46.49453, 46.52725, 46.51107, 46.61094, 46.57211, 46.7765, 
    46.68849, 46.91796, 46.86308, 46.93112, 46.89642, 46.95587, 46.90236, 
    46.99506, 47.01522, 47.00144, 47.05443, 46.89939, 46.95893, 46.51061, 
    46.51325, 46.52555, 46.47146, 46.46815, 46.41862, 46.46271, 46.48147, 
    46.52916, 46.55732, 46.58411, 46.64299, 46.70871, 46.80061, 46.86664, 
    46.91088, 46.88377, 46.9077, 46.88094, 46.8684, 47.00766, 46.92946, 
    47.04681, 47.04032, 46.98721, 47.04105, 46.5151, 46.49992, 46.44715, 
    46.48845, 46.41322, 46.45531, 46.4795, 46.57289, 46.59344, 46.61245, 
    46.65001, 46.6982, 46.78268, 46.85619, 46.9233, 46.91838, 46.92011, 
    46.93508, 46.89798, 46.94118, 46.94841, 46.92947, 47.03945, 47.00804, 
    47.04018, 47.01974, 46.50486, 46.53041, 46.5166, 46.54256, 46.52426, 
    46.60557, 46.62994, 46.744, 46.69724, 46.77169, 46.70481, 46.71666, 
    46.77405, 46.70844, 46.85211, 46.75465, 46.93567, 46.83832, 46.94176, 
    46.92301, 46.95407, 46.98187, 47.01687, 47.08138, 47.06645, 47.12041, 
    46.56851, 46.60162, 46.59874, 46.63341, 46.65904, 46.71463, 46.80371, 
    46.77023, 46.83173, 46.84406, 46.75064, 46.80798, 46.62381, 46.65354, 
    46.63586, 46.57111, 46.7779, 46.67178, 46.86773, 46.81028, 46.9779, 
    46.89452, 47.05822, 47.12807, 47.19393, 47.27068, 46.61973, 46.59723, 
    46.63755, 46.69325, 46.74502, 46.81377, 46.82082, 46.83369, 46.86706, 
    46.89509, 46.83773, 46.90212, 46.66037, 46.78712, 46.58869, 46.64842, 
    46.68998, 46.67178, 46.76641, 46.78869, 46.87921, 46.83244, 47.11081, 
    46.9877, 47.32921, 47.23382, 46.58936, 46.61967, 46.72507, 46.67493, 
    46.81838, 46.85366, 46.88236, 46.91899, 46.92297, 46.94468, 46.9091, 
    46.94328, 46.81392, 46.87175, 46.71307, 46.75168, 46.73393, 46.71443, 
    46.7746, 46.83862, 46.84004, 46.86056, 46.91827, 46.81896, 47.12659, 
    46.93658, 46.65271, 46.711, 46.71939, 46.6968, 46.85012, 46.79457, 
    46.94415, 46.90375, 46.96996, 46.93706, 46.93221, 46.88996, 46.86363, 
    46.79711, 46.74298, 46.70008, 46.71006, 46.75719, 46.84255, 46.92331, 
    46.90561, 46.96493, 46.80798, 46.87378, 46.84834, 46.91469, 46.76933, 
    46.89296, 46.73769, 46.75132, 46.79347, 46.87821, 46.89703, 46.91703, 
    46.9047, 46.84473, 46.83492, 46.79246, 46.78071, 46.74836, 46.72155, 
    46.74603, 46.77173, 46.84477, 46.91055, 46.98226, 46.99982, 47.08343, 
    47.0153, 47.12764, 47.03203, 47.19755, 46.9002, 47.02932, 46.79541, 
    46.82063, 46.8662, 46.97077, 46.91438, 46.98035, 46.83455, 46.75879, 
    46.73925, 46.70268, 46.74009, 46.73705, 46.77283, 46.76133, 46.8472, 
    46.80108, 46.93208, 46.97984, 47.11473, 47.19734, 47.28146, 47.31855, 
    47.32985, 47.33457 ;

 FIRA_R =
  46.42476, 46.50126, 46.4864, 46.54806, 46.51388, 46.55423, 46.4403, 
    46.50428, 46.46345, 46.43168, 46.6676, 46.55082, 46.78905, 46.71459, 
    46.90166, 46.77744, 46.92671, 46.89813, 46.98426, 46.95959, 47.0696, 
    46.99564, 47.12669, 47.05197, 47.06364, 46.99319, 46.57437, 46.65305, 
    46.5697, 46.58092, 46.5759, 46.51457, 46.48362, 46.41895, 46.4307, 
    46.47822, 46.58597, 46.54943, 46.6416, 46.63952, 46.74205, 46.69583, 
    46.86813, 46.81918, 46.96062, 46.92506, 46.95894, 46.94867, 46.95908, 
    46.90691, 46.92926, 46.88337, 46.70448, 46.75705, 46.60018, 46.50573, 
    46.4431, 46.3986, 46.40489, 46.41687, 46.4785, 46.53646, 46.58061, 
    46.61013, 46.63922, 46.72712, 46.77374, 46.878, 46.85923, 46.89106, 
    46.92152, 46.97259, 46.96419, 46.98668, 46.89025, 46.95433, 46.84853, 
    46.87746, 46.64696, 46.5593, 46.52188, 46.48925, 46.40972, 46.46464, 
    46.44299, 46.49453, 46.52725, 46.51107, 46.61094, 46.57211, 46.7765, 
    46.68849, 46.91796, 46.86308, 46.93112, 46.89642, 46.95587, 46.90236, 
    46.99506, 47.01522, 47.00144, 47.05443, 46.89939, 46.95893, 46.51061, 
    46.51325, 46.52555, 46.47146, 46.46815, 46.41862, 46.46271, 46.48147, 
    46.52916, 46.55732, 46.58411, 46.64299, 46.70871, 46.80061, 46.86664, 
    46.91088, 46.88377, 46.9077, 46.88094, 46.8684, 47.00766, 46.92946, 
    47.04681, 47.04032, 46.98721, 47.04105, 46.5151, 46.49992, 46.44715, 
    46.48845, 46.41322, 46.45531, 46.4795, 46.57289, 46.59344, 46.61245, 
    46.65001, 46.6982, 46.78268, 46.85619, 46.9233, 46.91838, 46.92011, 
    46.93508, 46.89798, 46.94118, 46.94841, 46.92947, 47.03945, 47.00804, 
    47.04018, 47.01974, 46.50486, 46.53041, 46.5166, 46.54256, 46.52426, 
    46.60557, 46.62994, 46.744, 46.69724, 46.77169, 46.70481, 46.71666, 
    46.77405, 46.70844, 46.85211, 46.75465, 46.93567, 46.83832, 46.94176, 
    46.92301, 46.95407, 46.98187, 47.01687, 47.08138, 47.06645, 47.12041, 
    46.56851, 46.60162, 46.59874, 46.63341, 46.65904, 46.71463, 46.80371, 
    46.77023, 46.83173, 46.84406, 46.75064, 46.80798, 46.62381, 46.65354, 
    46.63586, 46.57111, 46.7779, 46.67178, 46.86773, 46.81028, 46.9779, 
    46.89452, 47.05822, 47.12807, 47.19393, 47.27068, 46.61973, 46.59723, 
    46.63755, 46.69325, 46.74502, 46.81377, 46.82082, 46.83369, 46.86706, 
    46.89509, 46.83773, 46.90212, 46.66037, 46.78712, 46.58869, 46.64842, 
    46.68998, 46.67178, 46.76641, 46.78869, 46.87921, 46.83244, 47.11081, 
    46.9877, 47.32921, 47.23382, 46.58936, 46.61967, 46.72507, 46.67493, 
    46.81838, 46.85366, 46.88236, 46.91899, 46.92297, 46.94468, 46.9091, 
    46.94328, 46.81392, 46.87175, 46.71307, 46.75168, 46.73393, 46.71443, 
    46.7746, 46.83862, 46.84004, 46.86056, 46.91827, 46.81896, 47.12659, 
    46.93658, 46.65271, 46.711, 46.71939, 46.6968, 46.85012, 46.79457, 
    46.94415, 46.90375, 46.96996, 46.93706, 46.93221, 46.88996, 46.86363, 
    46.79711, 46.74298, 46.70008, 46.71006, 46.75719, 46.84255, 46.92331, 
    46.90561, 46.96493, 46.80798, 46.87378, 46.84834, 46.91469, 46.76933, 
    46.89296, 46.73769, 46.75132, 46.79347, 46.87821, 46.89703, 46.91703, 
    46.9047, 46.84473, 46.83492, 46.79246, 46.78071, 46.74836, 46.72155, 
    46.74603, 46.77173, 46.84477, 46.91055, 46.98226, 46.99982, 47.08343, 
    47.0153, 47.12764, 47.03203, 47.19755, 46.9002, 47.02932, 46.79541, 
    46.82063, 46.8662, 46.97077, 46.91438, 46.98035, 46.83455, 46.75879, 
    46.73925, 46.70268, 46.74009, 46.73705, 46.77283, 46.76133, 46.8472, 
    46.80108, 46.93208, 46.97984, 47.11473, 47.19734, 47.28146, 47.31855, 
    47.32985, 47.33457 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  260.7709, 260.8474, 260.8326, 260.8942, 260.86, 260.9004, 260.7864, 
    260.8504, 260.8096, 260.7778, 261.0137, 260.897, 261.1352, 261.0607, 
    261.2478, 261.1236, 261.2729, 261.2443, 261.3304, 261.3057, 261.4157, 
    261.3418, 261.4728, 261.3981, 261.4098, 261.3393, 260.9205, 260.9992, 
    260.9158, 260.9271, 260.922, 260.8607, 260.8298, 260.7651, 260.7769, 
    260.8244, 260.9321, 260.8956, 260.9877, 260.9857, 261.0882, 261.042, 
    261.2143, 261.1653, 261.3068, 261.2712, 261.3051, 261.2948, 261.3052, 
    261.2531, 261.2754, 261.2295, 261.0506, 261.1032, 260.9463, 260.8519, 
    260.7892, 260.7448, 260.751, 260.763, 260.8246, 260.8826, 260.9268, 
    260.9563, 260.9854, 261.0733, 261.1199, 261.2242, 261.2054, 261.2372, 
    261.2677, 261.3187, 261.3103, 261.3328, 261.2364, 261.3005, 261.1947, 
    261.2236, 260.9931, 260.9055, 260.868, 260.8354, 260.7559, 260.8108, 
    260.7891, 260.8407, 260.8734, 260.8572, 260.9571, 260.9182, 261.1227, 
    261.0346, 261.2641, 261.2092, 261.2773, 261.2426, 261.302, 261.2485, 
    261.3412, 261.3614, 261.3476, 261.4006, 261.2455, 261.3051, 260.8568, 
    260.8594, 260.8717, 260.8176, 260.8143, 260.7648, 260.8089, 260.8276, 
    260.8753, 260.9035, 260.9303, 260.9891, 261.0548, 261.1468, 261.2128, 
    261.257, 261.2299, 261.2538, 261.2271, 261.2145, 261.3538, 261.2756, 
    261.3929, 261.3865, 261.3333, 261.3872, 260.8612, 260.8461, 260.7933, 
    260.8346, 260.7594, 260.8015, 260.8257, 260.919, 260.9396, 260.9586, 
    260.9962, 261.0443, 261.1288, 261.2023, 261.2694, 261.2645, 261.2663, 
    261.2812, 261.2441, 261.2873, 261.2946, 261.2756, 261.3856, 261.3542, 
    261.3863, 261.3659, 260.851, 260.8766, 260.8627, 260.8887, 260.8704, 
    260.9517, 260.9761, 261.0901, 261.0434, 261.1178, 261.051, 261.0628, 
    261.1202, 261.0546, 261.1982, 261.1008, 261.2818, 261.1845, 261.2879, 
    261.2692, 261.3002, 261.328, 261.363, 261.4275, 261.4126, 261.4666, 
    260.9146, 260.9478, 260.9449, 260.9796, 261.0052, 261.0608, 261.1498, 
    261.1164, 261.1779, 261.1902, 261.0968, 261.1541, 260.9699, 260.9997, 
    260.982, 260.9172, 261.1241, 261.0179, 261.2139, 261.1564, 261.324, 
    261.2407, 261.4044, 261.4742, 261.5401, 261.6168, 260.9659, 260.9434, 
    260.9837, 261.0394, 261.0912, 261.1599, 261.167, 261.1798, 261.2132, 
    261.2412, 261.1839, 261.2483, 261.0065, 261.1333, 260.9348, 260.9946, 
    261.0361, 261.0179, 261.1125, 261.1348, 261.2253, 261.1786, 261.4569, 
    261.3338, 261.6754, 261.58, 260.9355, 260.9658, 261.0712, 261.0211, 
    261.1645, 261.1998, 261.2285, 261.2651, 261.2691, 261.2908, 261.2552, 
    261.2894, 261.1601, 261.2179, 261.0592, 261.0978, 261.0801, 261.0606, 
    261.1207, 261.1848, 261.1862, 261.2067, 261.2644, 261.1651, 261.4727, 
    261.2827, 260.9988, 261.0571, 261.0655, 261.0429, 261.1963, 261.1407, 
    261.2903, 261.2499, 261.3161, 261.2832, 261.2784, 261.2361, 261.2098, 
    261.1432, 261.0891, 261.0462, 261.0562, 261.1033, 261.1887, 261.2694, 
    261.2518, 261.3111, 261.1541, 261.2199, 261.1945, 261.2608, 261.1155, 
    261.2391, 261.0838, 261.0975, 261.1396, 261.2244, 261.2432, 261.2632, 
    261.2509, 261.1909, 261.1811, 261.1386, 261.1269, 261.0945, 261.0677, 
    261.0922, 261.1179, 261.1909, 261.2567, 261.3284, 261.346, 261.4296, 
    261.3615, 261.4738, 261.3782, 261.5437, 261.2463, 261.3755, 261.1415, 
    261.1668, 261.2123, 261.3169, 261.2605, 261.3265, 261.1807, 261.1049, 
    261.0854, 261.0488, 261.0862, 261.0832, 261.119, 261.1075, 261.1933, 
    261.1472, 261.2782, 261.326, 261.4609, 261.5435, 261.6276, 261.6647, 
    261.676, 261.6807 ;

 FIRE_R =
  260.7709, 260.8474, 260.8326, 260.8942, 260.86, 260.9004, 260.7864, 
    260.8504, 260.8096, 260.7778, 261.0137, 260.897, 261.1352, 261.0607, 
    261.2478, 261.1236, 261.2729, 261.2443, 261.3304, 261.3057, 261.4157, 
    261.3418, 261.4728, 261.3981, 261.4098, 261.3393, 260.9205, 260.9992, 
    260.9158, 260.9271, 260.922, 260.8607, 260.8298, 260.7651, 260.7769, 
    260.8244, 260.9321, 260.8956, 260.9877, 260.9857, 261.0882, 261.042, 
    261.2143, 261.1653, 261.3068, 261.2712, 261.3051, 261.2948, 261.3052, 
    261.2531, 261.2754, 261.2295, 261.0506, 261.1032, 260.9463, 260.8519, 
    260.7892, 260.7448, 260.751, 260.763, 260.8246, 260.8826, 260.9268, 
    260.9563, 260.9854, 261.0733, 261.1199, 261.2242, 261.2054, 261.2372, 
    261.2677, 261.3187, 261.3103, 261.3328, 261.2364, 261.3005, 261.1947, 
    261.2236, 260.9931, 260.9055, 260.868, 260.8354, 260.7559, 260.8108, 
    260.7891, 260.8407, 260.8734, 260.8572, 260.9571, 260.9182, 261.1227, 
    261.0346, 261.2641, 261.2092, 261.2773, 261.2426, 261.302, 261.2485, 
    261.3412, 261.3614, 261.3476, 261.4006, 261.2455, 261.3051, 260.8568, 
    260.8594, 260.8717, 260.8176, 260.8143, 260.7648, 260.8089, 260.8276, 
    260.8753, 260.9035, 260.9303, 260.9891, 261.0548, 261.1468, 261.2128, 
    261.257, 261.2299, 261.2538, 261.2271, 261.2145, 261.3538, 261.2756, 
    261.3929, 261.3865, 261.3333, 261.3872, 260.8612, 260.8461, 260.7933, 
    260.8346, 260.7594, 260.8015, 260.8257, 260.919, 260.9396, 260.9586, 
    260.9962, 261.0443, 261.1288, 261.2023, 261.2694, 261.2645, 261.2663, 
    261.2812, 261.2441, 261.2873, 261.2946, 261.2756, 261.3856, 261.3542, 
    261.3863, 261.3659, 260.851, 260.8766, 260.8627, 260.8887, 260.8704, 
    260.9517, 260.9761, 261.0901, 261.0434, 261.1178, 261.051, 261.0628, 
    261.1202, 261.0546, 261.1982, 261.1008, 261.2818, 261.1845, 261.2879, 
    261.2692, 261.3002, 261.328, 261.363, 261.4275, 261.4126, 261.4666, 
    260.9146, 260.9478, 260.9449, 260.9796, 261.0052, 261.0608, 261.1498, 
    261.1164, 261.1779, 261.1902, 261.0968, 261.1541, 260.9699, 260.9997, 
    260.982, 260.9172, 261.1241, 261.0179, 261.2139, 261.1564, 261.324, 
    261.2407, 261.4044, 261.4742, 261.5401, 261.6168, 260.9659, 260.9434, 
    260.9837, 261.0394, 261.0912, 261.1599, 261.167, 261.1798, 261.2132, 
    261.2412, 261.1839, 261.2483, 261.0065, 261.1333, 260.9348, 260.9946, 
    261.0361, 261.0179, 261.1125, 261.1348, 261.2253, 261.1786, 261.4569, 
    261.3338, 261.6754, 261.58, 260.9355, 260.9658, 261.0712, 261.0211, 
    261.1645, 261.1998, 261.2285, 261.2651, 261.2691, 261.2908, 261.2552, 
    261.2894, 261.1601, 261.2179, 261.0592, 261.0978, 261.0801, 261.0606, 
    261.1207, 261.1848, 261.1862, 261.2067, 261.2644, 261.1651, 261.4727, 
    261.2827, 260.9988, 261.0571, 261.0655, 261.0429, 261.1963, 261.1407, 
    261.2903, 261.2499, 261.3161, 261.2832, 261.2784, 261.2361, 261.2098, 
    261.1432, 261.0891, 261.0462, 261.0562, 261.1033, 261.1887, 261.2694, 
    261.2518, 261.3111, 261.1541, 261.2199, 261.1945, 261.2608, 261.1155, 
    261.2391, 261.0838, 261.0975, 261.1396, 261.2244, 261.2432, 261.2632, 
    261.2509, 261.1909, 261.1811, 261.1386, 261.1269, 261.0945, 261.0677, 
    261.0922, 261.1179, 261.1909, 261.2567, 261.3284, 261.346, 261.4296, 
    261.3615, 261.4738, 261.3782, 261.5437, 261.2463, 261.3755, 261.1415, 
    261.1668, 261.2123, 261.3169, 261.2605, 261.3265, 261.1807, 261.1049, 
    261.0854, 261.0488, 261.0862, 261.0832, 261.119, 261.1075, 261.1933, 
    261.1472, 261.2782, 261.326, 261.4609, 261.5435, 261.6276, 261.6647, 
    261.676, 261.6807 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  320.5223, 321.4778, 321.2922, 322.0623, 321.6353, 322.1394, 320.7163, 
    321.5155, 321.0055, 320.6087, 323.5557, 322.0967, 325.0722, 324.1422, 
    326.4785, 324.9272, 326.7912, 326.4343, 327.5097, 327.2017, 328.5755, 
    327.6518, 329.2881, 328.3553, 328.501, 327.6213, 322.3909, 323.3739, 
    322.3325, 322.4727, 322.4099, 321.644, 321.2576, 320.4496, 320.5964, 
    321.19, 322.5358, 322.0794, 323.2306, 323.2046, 324.4852, 323.9079, 
    326.0596, 325.4484, 327.2145, 326.7704, 327.1936, 327.0654, 327.1953, 
    326.5439, 326.823, 326.2499, 324.0159, 324.6725, 322.7133, 321.5338, 
    320.7513, 320.1955, 320.274, 320.4237, 321.1935, 321.9174, 322.4688, 
    322.8375, 323.2008, 324.2989, 324.881, 326.1829, 325.9484, 326.3459, 
    326.7263, 327.364, 327.2592, 327.54, 326.3358, 327.136, 325.8148, 
    326.1762, 323.2979, 322.2026, 321.7355, 321.3278, 320.3344, 321.0204, 
    320.7499, 321.3936, 321.8023, 321.6002, 322.8476, 322.3627, 324.9155, 
    323.8163, 326.6819, 325.9966, 326.8462, 326.4128, 327.1552, 326.4871, 
    327.6446, 327.8964, 327.7243, 328.3859, 326.45, 327.1935, 321.5945, 
    321.6274, 321.7811, 321.1055, 321.0643, 320.4456, 320.9963, 321.2306, 
    321.8261, 322.178, 322.5125, 323.248, 324.0688, 325.2165, 326.041, 
    326.5934, 326.2548, 326.5537, 326.2195, 326.0629, 327.8019, 326.8255, 
    328.2907, 328.2097, 327.5466, 328.2188, 321.6506, 321.461, 320.8019, 
    321.3177, 320.3782, 320.9039, 321.206, 322.3724, 322.6291, 322.8664, 
    323.3356, 323.9374, 324.9926, 325.9106, 326.7485, 326.6871, 326.7087, 
    326.8957, 326.4323, 326.9717, 327.0621, 326.8256, 328.1989, 327.8066, 
    328.208, 327.9527, 321.5226, 321.8418, 321.6693, 321.9936, 321.765, 
    322.7806, 323.0851, 324.5096, 323.9255, 324.8554, 324.0201, 324.168, 
    324.885, 324.0653, 325.8596, 324.6427, 326.9029, 325.6876, 326.979, 
    326.7448, 327.1328, 327.4799, 327.9169, 328.7224, 328.5359, 329.2097, 
    322.3177, 322.7314, 322.6953, 323.1283, 323.4485, 324.1426, 325.2552, 
    324.837, 325.605, 325.759, 324.5924, 325.3084, 323.0084, 323.3798, 
    323.1589, 322.3501, 324.9329, 323.6076, 326.0546, 325.3371, 327.4304, 
    326.3893, 328.4332, 329.3055, 330.1275, 331.0859, 322.9574, 322.6764, 
    323.1799, 323.8758, 324.5222, 325.3808, 325.4688, 325.6295, 326.0462, 
    326.3963, 325.6801, 326.484, 323.4653, 325.048, 322.5698, 323.3159, 
    323.8349, 323.6076, 324.7892, 325.0675, 326.198, 325.6139, 329.09, 
    327.5528, 331.8164, 330.6257, 322.5781, 322.9566, 324.2732, 323.6469, 
    325.4383, 325.8789, 326.2373, 326.6948, 326.7444, 327.0155, 326.5712, 
    326.998, 325.3827, 326.1047, 324.1231, 324.6054, 324.3837, 324.1402, 
    324.8915, 325.6913, 325.7089, 325.9651, 326.6862, 325.4456, 329.2873, 
    326.9147, 323.3693, 324.0975, 324.2021, 323.92, 325.8347, 325.1411, 
    327.0089, 326.5044, 327.3311, 326.9203, 326.8598, 326.3322, 326.0034, 
    325.1728, 324.4968, 323.9609, 324.0856, 324.6742, 325.7403, 326.7487, 
    326.5277, 327.2683, 325.3084, 326.1302, 325.8125, 326.641, 324.8257, 
    326.3701, 324.4306, 324.6009, 325.1273, 326.1856, 326.4204, 326.6702, 
    326.5162, 325.7674, 325.645, 325.1146, 324.9679, 324.5638, 324.229, 
    324.5348, 324.8558, 325.768, 326.5894, 327.4847, 327.704, 328.7482, 
    327.8975, 329.3004, 328.1067, 330.1731, 326.4603, 328.0726, 325.1514, 
    325.4664, 326.0356, 327.3414, 326.6371, 327.4611, 325.6402, 324.6943, 
    324.4501, 323.9934, 324.4605, 324.4226, 324.8694, 324.7259, 325.7982, 
    325.2223, 326.8582, 327.4547, 329.1389, 330.1702, 331.2203, 331.6834, 
    331.8243, 331.8832 ;

 FSH_G =
  327.1818, 328.1378, 327.9521, 328.7227, 328.2954, 328.7998, 327.3759, 
    328.1755, 327.6652, 327.2682, 330.2169, 328.7571, 331.7343, 330.8037, 
    333.1414, 331.5893, 333.4543, 333.0971, 334.1732, 333.865, 335.2396, 
    334.3154, 335.9527, 335.0193, 335.1651, 334.2849, 329.0515, 330.035, 
    328.993, 329.1334, 329.0705, 328.3041, 327.9174, 327.1091, 327.256, 
    327.8499, 329.1965, 328.7397, 329.8916, 329.8656, 331.1469, 330.5693, 
    332.7222, 332.1107, 333.8779, 333.4335, 333.8569, 333.7286, 333.8586, 
    333.2069, 333.4861, 332.9127, 330.6774, 331.3344, 329.3741, 328.1938, 
    327.4109, 326.8548, 326.9334, 327.0832, 327.8533, 328.5777, 329.1294, 
    329.4983, 329.8618, 330.9605, 331.5429, 332.8456, 332.6111, 333.0088, 
    333.3893, 334.0275, 333.9225, 334.2035, 332.9986, 333.7993, 332.4773, 
    332.8389, 329.9589, 328.8631, 328.3956, 327.9877, 326.9938, 327.6801, 
    327.4096, 328.0536, 328.4625, 328.2603, 329.5084, 329.0232, 331.5775, 
    330.4776, 333.3449, 332.6592, 333.5093, 333.0757, 333.8185, 333.15, 
    334.3082, 334.5601, 334.3879, 335.0499, 333.1129, 333.8568, 328.2546, 
    328.2875, 328.4413, 327.7654, 327.7241, 327.105, 327.656, 327.8905, 
    328.4863, 328.8384, 329.1732, 329.909, 330.7303, 331.8787, 332.7037, 
    333.2564, 332.9176, 333.2167, 332.8823, 332.7256, 334.4656, 333.4886, 
    334.9547, 334.8736, 334.2101, 334.8828, 328.3107, 328.121, 327.4616, 
    327.9776, 327.0376, 327.5636, 327.8659, 329.033, 329.2897, 329.5273, 
    329.9967, 330.5988, 331.6547, 332.5732, 333.4115, 333.3502, 333.3717, 
    333.5588, 333.0952, 333.6349, 333.7253, 333.4887, 334.8628, 334.4703, 
    334.8719, 334.6165, 328.1827, 328.502, 328.3295, 328.6539, 328.4252, 
    329.4414, 329.746, 331.1713, 330.5869, 331.5174, 330.6816, 330.8296, 
    331.547, 330.7269, 332.5222, 331.3045, 333.5661, 332.35, 333.6422, 
    333.4079, 333.796, 334.1434, 334.5806, 335.3866, 335.2, 335.8741, 
    328.9782, 329.3921, 329.356, 329.7893, 330.1096, 330.8042, 331.9174, 
    331.4989, 332.2674, 332.4215, 331.2542, 331.9707, 329.6693, 330.0409, 
    329.8199, 329.0107, 331.5949, 330.2688, 332.7172, 331.9994, 334.0938, 
    333.0522, 335.0973, 335.97, 336.7926, 337.7515, 329.6183, 329.3371, 
    329.8409, 330.5372, 331.184, 332.0431, 332.1312, 332.292, 332.7088, 
    333.0591, 332.3425, 333.1469, 330.1265, 331.7101, 329.2304, 329.977, 
    330.4963, 330.2688, 331.4512, 331.7296, 332.8607, 332.2763, 335.7544, 
    334.2163, 338.4824, 337.291, 329.2387, 329.6175, 330.9348, 330.3082, 
    332.1006, 332.5415, 332.9001, 333.3578, 333.4075, 333.6787, 333.2342, 
    333.6613, 332.045, 332.7674, 330.7847, 331.2672, 331.0453, 330.8017, 
    331.5535, 332.3537, 332.3713, 332.6277, 333.3492, 332.1079, 335.9518, 
    333.5779, 330.0304, 330.759, 330.8637, 330.5814, 332.4973, 331.8032, 
    333.6721, 333.1673, 333.9945, 333.5835, 333.5229, 332.995, 332.666, 
    331.8349, 331.1586, 330.6224, 330.7471, 331.3361, 332.4028, 333.4117, 
    333.1907, 333.9317, 331.9707, 332.7929, 332.475, 333.304, 331.4877, 
    333.0329, 331.0924, 331.2627, 331.7894, 332.8483, 333.0833, 333.3333, 
    333.1791, 332.4299, 332.3074, 331.7767, 331.6299, 331.2256, 330.8906, 
    331.1966, 331.5178, 332.4305, 333.2523, 334.1483, 334.3676, 335.4124, 
    334.5612, 335.9649, 334.7705, 336.8382, 333.1232, 334.7364, 331.8135, 
    332.1288, 332.6982, 334.0048, 333.3001, 334.1245, 332.3026, 331.3561, 
    331.1118, 330.6549, 331.1223, 331.0843, 331.5314, 331.3878, 332.4608, 
    331.8845, 333.5213, 334.1181, 335.8033, 336.8353, 337.886, 338.3493, 
    338.4904, 338.5493 ;

 FSH_NODYNLNDUSE =
  320.5223, 321.4778, 321.2922, 322.0623, 321.6353, 322.1394, 320.7163, 
    321.5155, 321.0055, 320.6087, 323.5557, 322.0967, 325.0722, 324.1422, 
    326.4785, 324.9272, 326.7912, 326.4343, 327.5097, 327.2017, 328.5755, 
    327.6518, 329.2881, 328.3553, 328.501, 327.6213, 322.3909, 323.3739, 
    322.3325, 322.4727, 322.4099, 321.644, 321.2576, 320.4496, 320.5964, 
    321.19, 322.5358, 322.0794, 323.2306, 323.2046, 324.4852, 323.9079, 
    326.0596, 325.4484, 327.2145, 326.7704, 327.1936, 327.0654, 327.1953, 
    326.5439, 326.823, 326.2499, 324.0159, 324.6725, 322.7133, 321.5338, 
    320.7513, 320.1955, 320.274, 320.4237, 321.1935, 321.9174, 322.4688, 
    322.8375, 323.2008, 324.2989, 324.881, 326.1829, 325.9484, 326.3459, 
    326.7263, 327.364, 327.2592, 327.54, 326.3358, 327.136, 325.8148, 
    326.1762, 323.2979, 322.2026, 321.7355, 321.3278, 320.3344, 321.0204, 
    320.7499, 321.3936, 321.8023, 321.6002, 322.8476, 322.3627, 324.9155, 
    323.8163, 326.6819, 325.9966, 326.8462, 326.4128, 327.1552, 326.4871, 
    327.6446, 327.8964, 327.7243, 328.3859, 326.45, 327.1935, 321.5945, 
    321.6274, 321.7811, 321.1055, 321.0643, 320.4456, 320.9963, 321.2306, 
    321.8261, 322.178, 322.5125, 323.248, 324.0688, 325.2165, 326.041, 
    326.5934, 326.2548, 326.5537, 326.2195, 326.0629, 327.8019, 326.8255, 
    328.2907, 328.2097, 327.5466, 328.2188, 321.6506, 321.461, 320.8019, 
    321.3177, 320.3782, 320.9039, 321.206, 322.3724, 322.6291, 322.8664, 
    323.3356, 323.9374, 324.9926, 325.9106, 326.7485, 326.6871, 326.7087, 
    326.8957, 326.4323, 326.9717, 327.0621, 326.8256, 328.1989, 327.8066, 
    328.208, 327.9527, 321.5226, 321.8418, 321.6693, 321.9936, 321.765, 
    322.7806, 323.0851, 324.5096, 323.9255, 324.8554, 324.0201, 324.168, 
    324.885, 324.0653, 325.8596, 324.6427, 326.9029, 325.6876, 326.979, 
    326.7448, 327.1328, 327.4799, 327.9169, 328.7224, 328.5359, 329.2097, 
    322.3177, 322.7314, 322.6953, 323.1283, 323.4485, 324.1426, 325.2552, 
    324.837, 325.605, 325.759, 324.5924, 325.3084, 323.0084, 323.3798, 
    323.1589, 322.3501, 324.9329, 323.6076, 326.0546, 325.3371, 327.4304, 
    326.3893, 328.4332, 329.3055, 330.1275, 331.0859, 322.9574, 322.6764, 
    323.1799, 323.8758, 324.5222, 325.3808, 325.4688, 325.6295, 326.0462, 
    326.3963, 325.6801, 326.484, 323.4653, 325.048, 322.5698, 323.3159, 
    323.8349, 323.6076, 324.7892, 325.0675, 326.198, 325.6139, 329.09, 
    327.5528, 331.8164, 330.6257, 322.5781, 322.9566, 324.2732, 323.6469, 
    325.4383, 325.8789, 326.2373, 326.6948, 326.7444, 327.0155, 326.5712, 
    326.998, 325.3827, 326.1047, 324.1231, 324.6054, 324.3837, 324.1402, 
    324.8915, 325.6913, 325.7089, 325.9651, 326.6862, 325.4456, 329.2873, 
    326.9147, 323.3693, 324.0975, 324.2021, 323.92, 325.8347, 325.1411, 
    327.0089, 326.5044, 327.3311, 326.9203, 326.8598, 326.3322, 326.0034, 
    325.1728, 324.4968, 323.9609, 324.0856, 324.6742, 325.7403, 326.7487, 
    326.5277, 327.2683, 325.3084, 326.1302, 325.8125, 326.641, 324.8257, 
    326.3701, 324.4306, 324.6009, 325.1273, 326.1856, 326.4204, 326.6702, 
    326.5162, 325.7674, 325.645, 325.1146, 324.9679, 324.5638, 324.229, 
    324.5348, 324.8558, 325.768, 326.5894, 327.4847, 327.704, 328.7482, 
    327.8975, 329.3004, 328.1067, 330.1731, 326.4603, 328.0726, 325.1514, 
    325.4664, 326.0356, 327.3414, 326.6371, 327.4611, 325.6402, 324.6943, 
    324.4501, 323.9934, 324.4605, 324.4226, 324.8694, 324.7259, 325.7982, 
    325.2223, 326.8582, 327.4547, 329.1389, 330.1702, 331.2203, 331.6834, 
    331.8243, 331.8832 ;

 FSH_R =
  320.5223, 321.4778, 321.2922, 322.0623, 321.6353, 322.1394, 320.7163, 
    321.5155, 321.0055, 320.6087, 323.5557, 322.0967, 325.0722, 324.1422, 
    326.4785, 324.9272, 326.7912, 326.4343, 327.5097, 327.2017, 328.5755, 
    327.6518, 329.2881, 328.3553, 328.501, 327.6213, 322.3909, 323.3739, 
    322.3325, 322.4727, 322.4099, 321.644, 321.2576, 320.4496, 320.5964, 
    321.19, 322.5358, 322.0794, 323.2306, 323.2046, 324.4852, 323.9079, 
    326.0596, 325.4484, 327.2145, 326.7704, 327.1936, 327.0654, 327.1953, 
    326.5439, 326.823, 326.2499, 324.0159, 324.6725, 322.7133, 321.5338, 
    320.7513, 320.1955, 320.274, 320.4237, 321.1935, 321.9174, 322.4688, 
    322.8375, 323.2008, 324.2989, 324.881, 326.1829, 325.9484, 326.3459, 
    326.7263, 327.364, 327.2592, 327.54, 326.3358, 327.136, 325.8148, 
    326.1762, 323.2979, 322.2026, 321.7355, 321.3278, 320.3344, 321.0204, 
    320.7499, 321.3936, 321.8023, 321.6002, 322.8476, 322.3627, 324.9155, 
    323.8163, 326.6819, 325.9966, 326.8462, 326.4128, 327.1552, 326.4871, 
    327.6446, 327.8964, 327.7243, 328.3859, 326.45, 327.1935, 321.5945, 
    321.6274, 321.7811, 321.1055, 321.0643, 320.4456, 320.9963, 321.2306, 
    321.8261, 322.178, 322.5125, 323.248, 324.0688, 325.2165, 326.041, 
    326.5934, 326.2548, 326.5537, 326.2195, 326.0629, 327.8019, 326.8255, 
    328.2907, 328.2097, 327.5466, 328.2188, 321.6506, 321.461, 320.8019, 
    321.3177, 320.3782, 320.9039, 321.206, 322.3724, 322.6291, 322.8664, 
    323.3356, 323.9374, 324.9926, 325.9106, 326.7485, 326.6871, 326.7087, 
    326.8957, 326.4323, 326.9717, 327.0621, 326.8256, 328.1989, 327.8066, 
    328.208, 327.9527, 321.5226, 321.8418, 321.6693, 321.9936, 321.765, 
    322.7806, 323.0851, 324.5096, 323.9255, 324.8554, 324.0201, 324.168, 
    324.885, 324.0653, 325.8596, 324.6427, 326.9029, 325.6876, 326.979, 
    326.7448, 327.1328, 327.4799, 327.9169, 328.7224, 328.5359, 329.2097, 
    322.3177, 322.7314, 322.6953, 323.1283, 323.4485, 324.1426, 325.2552, 
    324.837, 325.605, 325.759, 324.5924, 325.3084, 323.0084, 323.3798, 
    323.1589, 322.3501, 324.9329, 323.6076, 326.0546, 325.3371, 327.4304, 
    326.3893, 328.4332, 329.3055, 330.1275, 331.0859, 322.9574, 322.6764, 
    323.1799, 323.8758, 324.5222, 325.3808, 325.4688, 325.6295, 326.0462, 
    326.3963, 325.6801, 326.484, 323.4653, 325.048, 322.5698, 323.3159, 
    323.8349, 323.6076, 324.7892, 325.0675, 326.198, 325.6139, 329.09, 
    327.5528, 331.8164, 330.6257, 322.5781, 322.9566, 324.2732, 323.6469, 
    325.4383, 325.8789, 326.2373, 326.6948, 326.7444, 327.0155, 326.5712, 
    326.998, 325.3827, 326.1047, 324.1231, 324.6054, 324.3837, 324.1402, 
    324.8915, 325.6913, 325.7089, 325.9651, 326.6862, 325.4456, 329.2873, 
    326.9147, 323.3693, 324.0975, 324.2021, 323.92, 325.8347, 325.1411, 
    327.0089, 326.5044, 327.3311, 326.9203, 326.8598, 326.3322, 326.0034, 
    325.1728, 324.4968, 323.9609, 324.0856, 324.6742, 325.7403, 326.7487, 
    326.5277, 327.2683, 325.3084, 326.1302, 325.8125, 326.641, 324.8257, 
    326.3701, 324.4306, 324.6009, 325.1273, 326.1856, 326.4204, 326.6702, 
    326.5162, 325.7674, 325.645, 325.1146, 324.9679, 324.5638, 324.229, 
    324.5348, 324.8558, 325.768, 326.5894, 327.4847, 327.704, 328.7482, 
    327.8975, 329.3004, 328.1067, 330.1731, 326.4603, 328.0726, 325.1514, 
    325.4664, 326.0356, 327.3414, 326.6371, 327.4611, 325.6402, 324.6943, 
    324.4501, 323.9934, 324.4605, 324.4226, 324.8694, 324.7259, 325.7982, 
    325.2223, 326.8582, 327.4547, 329.1389, 330.1702, 331.2203, 331.6834, 
    331.8243, 331.8832 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.659477, -6.660025, -6.659921, -6.660357, -6.66012, -6.660402, -6.659593, 
    -6.660043, -6.659759, -6.659534, -6.661191, -6.660378, -6.662084, 
    -6.661556, -6.662898, -6.661995, -6.663082, -6.662882, -6.663509, 
    -6.663331, -6.664111, -6.663592, -6.664534, -6.663993, -6.664073, 
    -6.663573, -6.660552, -6.661087, -6.660518, -6.660595, -6.660563, 
    -6.66012, -6.659891, -6.659443, -6.659526, -6.659859, -6.660629, 
    -6.660375, -6.661038, -6.661023, -6.661755, -6.661425, -6.662665, 
    -6.662314, -6.663338, -6.663079, -6.663324, -6.663251, -6.663325, 
    -6.662945, -6.663107, -6.662777, -6.661484, -6.66186, -6.660735, 
    -6.660043, -6.659611, -6.659297, -6.659341, -6.659423, -6.659861, 
    -6.660282, -6.6606, -6.660811, -6.661021, -6.661628, -6.661973, 
    -6.662731, -6.662603, -6.662827, -6.663054, -6.663422, -6.663363, 
    -6.663523, -6.662827, -6.663286, -6.662529, -6.662734, -6.661041, 
    -6.660445, -6.660161, -6.65994, -6.659374, -6.659763, -6.659609, 
    -6.659983, -6.660216, -6.660102, -6.660817, -6.660538, -6.661994, 
    -6.661366, -6.663027, -6.66263, -6.663124, -6.662873, -6.663299, 
    -6.662916, -6.663585, -6.663727, -6.66363, -6.664017, -6.662894, 
    -6.663321, -6.660097, -6.660116, -6.660205, -6.659811, -6.659789, 
    -6.659439, -6.659754, -6.659884, -6.660232, -6.660431, -6.660622, 
    -6.661044, -6.66151, -6.662173, -6.662655, -6.662978, -6.662783, 
    -6.662955, -6.662761, -6.662672, -6.663671, -6.663106, -6.663961, 
    -6.663915, -6.663525, -6.66392, -6.660129, -6.660023, -6.659641, 
    -6.65994, -6.659401, -6.659698, -6.659866, -6.660535, -6.660691, 
    -6.660825, -6.661097, -6.661441, -6.662045, -6.662576, -6.663068, 
    -6.663033, -6.663045, -6.663151, -6.662883, -6.663195, -6.663244, 
    -6.663111, -6.663909, -6.663681, -6.663914, -6.663767, -6.660058, 
    -6.660239, -6.660141, -6.660324, -6.660192, -6.660768, -6.66094, 
    -6.66176, -6.661432, -6.661964, -6.661489, -6.661571, -6.661966, 
    -6.661517, -6.66254, -6.661832, -6.663155, -6.662432, -6.663199, 
    -6.663066, -6.663291, -6.663489, -6.663744, -6.664207, -6.664101, 
    -6.664494, -6.660512, -6.660744, -6.66073, -6.660977, -6.661159, 
    -6.661561, -6.662199, -6.661962, -6.662406, -6.662493, -6.661822, 
    -6.662227, -6.660904, -6.66111, -6.660993, -6.660526, -6.662006, 
    -6.661242, -6.662662, -6.662248, -6.66346, -6.662849, -6.664041, 
    -6.664534, -6.665031, -6.665576, -6.660878, -6.660719, -6.661009, 
    -6.661397, -6.661777, -6.662272, -6.662327, -6.662417, -6.662662, 
    -6.662863, -6.662439, -6.662915, -6.661144, -6.662076, -6.660653, 
    -6.661072, -6.661377, -6.66125, -6.661936, -6.662096, -6.662742, 
    -6.662411, -6.664406, -6.663521, -6.666014, -6.66531, -6.660663, 
    -6.66088, -6.661629, -6.661274, -6.662309, -6.662561, -6.662773, 
    -6.663032, -6.663064, -6.663219, -6.662965, -6.663212, -6.662273, 
    -6.662693, -6.661552, -6.661825, -6.661702, -6.661561, -6.661994, 
    -6.662445, -6.662465, -6.662608, -6.66299, -6.662313, -6.6645, -6.663128, 
    -6.661117, -6.661522, -6.661593, -6.661434, -6.662536, -6.662135, 
    -6.663217, -6.662926, -6.663405, -6.663166, -6.66313, -6.662827, 
    -6.662634, -6.662151, -6.661761, -6.661458, -6.66153, -6.661863, 
    -6.662475, -6.663063, -6.662932, -6.663369, -6.662233, -6.662703, 
    -6.662518, -6.663003, -6.661952, -6.662813, -6.661729, -6.661826, 
    -6.662127, -6.662727, -6.662878, -6.663017, -6.662933, -6.662492, 
    -6.662425, -6.662122, -6.662033, -6.661806, -6.661613, -6.661787, 
    -6.661967, -6.662497, -6.66297, -6.66349, -6.663622, -6.664203, 
    -6.663714, -6.664505, -6.663809, -6.665027, -6.66288, -6.663812, 
    -6.662144, -6.662326, -6.662643, -6.663396, -6.663002, -6.663469, 
    -6.662423, -6.661869, -6.661739, -6.661475, -6.661746, -6.661724, 
    -6.661982, -6.6619, -6.662515, -6.662185, -6.663126, -6.663468, 
    -6.664448, -6.665044, -6.665669, -6.66594, -6.666024, -6.666058 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.100726e-43, 5.605194e-45, 
    3.498145e-40, 2.53635e-43, 1.405053e-39, 2.860358e-40, 3.155876e-38, 
    8.419162e-39, 2.624818e-36, 5.766906e-38, 4.399989e-35, 1.071883e-36, 
    1.939966e-36, 5.068994e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.942727e-44, 1.401298e-45, 5.228945e-41, 3.049225e-42, 8.900133e-39, 
    1.278835e-39, 8.133579e-39, 4.660608e-39, 8.192598e-39, 4.676525e-40, 
    1.613396e-39, 1.244143e-40, 2.802597e-45, 7.286752e-44, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.121039e-44, 2.031883e-43, 9.19462e-41, 3.137227e-41, 
    1.924305e-40, 1.051815e-39, 1.695091e-38, 1.079296e-38, 3.593701e-38, 
    1.834622e-40, 6.345298e-39, 1.690947e-41, 8.899506e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.39622e-43, 1.401298e-45, 8.642228e-40, 3.915788e-41, 
    1.785855e-39, 2.594924e-40, 6.893387e-39, 3.6223e-40, 5.59756e-38, 
    1.61379e-37, 7.839023e-38, 1.212262e-36, 3.067653e-40, 8.134899e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.203895e-45, 1.017343e-42, 
    4.801269e-41, 5.826459e-40, 1.27116e-40, 4.881381e-40, 1.083344e-40, 
    5.302794e-41, 1.08715e-37, 1.632183e-39, 8.222793e-37, 5.898124e-37, 
    3.697471e-38, 6.123528e-37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.401298e-45, 3.47522e-43, 2.638505e-41, 1.15981e-39, 8.837471e-40, 
    9.726132e-40, 2.220196e-39, 2.83372e-40, 3.098589e-39, 4.600644e-39, 
    1.630998e-39, 5.640851e-37, 1.106896e-37, 5.856523e-37, 2.036912e-37, 0, 
    0, 0, 0, 0, 0, 0, 3.222986e-44, 1.401298e-45, 1.793662e-43, 2.802597e-45, 
    5.605194e-45, 2.073922e-43, 4.203895e-45, 2.089476e-41, 6.305843e-44, 
    2.292201e-39, 9.419528e-42, 3.198822e-39, 1.14138e-39, 6.244441e-39, 
    2.781966e-38, 1.755172e-37, 4.722894e-36, 2.230228e-36, 3.237457e-35, 0, 
    0, 0, 0, 0, 5.605194e-45, 1.221932e-42, 1.625506e-43, 6.366099e-42, 
    1.306851e-41, 4.904545e-44, 1.575059e-42, 0, 0, 0, 0, 2.606415e-43, 0, 
    5.110676e-41, 1.80207e-42, 2.251942e-38, 2.340813e-40, 1.471128e-36, 
    4.718157e-35, 1.069506e-33, 3.474821e-32, 0, 0, 0, 1.401298e-45, 
    3.503246e-44, 2.218255e-42, 3.358912e-42, 7.146622e-42, 4.912392e-41, 
    2.409084e-40, 9.066401e-42, 3.573101e-40, 0, 4.540207e-43, 0, 0, 
    1.401298e-45, 0, 1.289195e-43, 4.97461e-43, 9.84216e-41, 6.63655e-42, 
    2.034721e-35, 3.803153e-38, 4.371386e-31, 6.681893e-33, 0, 0, 
    9.809089e-45, 0, 2.907694e-42, 2.277671e-41, 1.173952e-40, 9.156785e-40, 
    1.139511e-39, 3.752387e-39, 5.277444e-40, 3.475073e-39, 2.237874e-42, 
    6.425234e-41, 4.203895e-45, 5.324934e-44, 1.821688e-44, 5.605194e-45, 
    2.129974e-43, 9.555454e-42, 1.034298e-41, 3.392263e-41, 8.898455e-40, 
    3.009989e-42, 4.420301e-35, 2.435304e-39, 0, 4.203895e-45, 7.006492e-45, 
    1.401298e-45, 1.856861e-41, 7.076557e-43, 3.645385e-39, 3.914247e-40, 
    1.470874e-38, 2.473112e-39, 1.896537e-39, 1.804298e-40, 4.040644e-41, 
    8.239635e-43, 3.082857e-44, 1.401298e-45, 4.203895e-45, 7.426882e-44, 
    1.200072e-41, 1.162563e-39, 4.354619e-40, 1.122507e-38, 1.572257e-42, 
    7.226917e-41, 1.677214e-41, 7.204426e-40, 1.541428e-43, 2.160732e-40, 
    2.242078e-44, 5.184804e-44, 6.628142e-43, 9.319896e-41, 2.685967e-40, 
    8.211385e-40, 4.12688e-40, 1.360801e-41, 7.683319e-42, 6.235778e-43, 
    3.082857e-43, 4.344025e-44, 8.407791e-45, 3.643376e-44, 1.793662e-43, 
    1.362482e-41, 5.731339e-40, 2.841443e-38, 7.189204e-38, 5.260623e-36, 
    1.626792e-37, 4.653514e-35, 3.901921e-37, 1.275646e-33, 3.229811e-40, 
    3.37117e-37, 7.426882e-43, 3.319676e-42, 4.69449e-41, 1.543183e-38, 
    7.080719e-40, 2.572929e-38, 7.512361e-42, 8.127531e-44, 2.382207e-44, 
    2.802597e-45, 2.522337e-44, 2.101948e-44, 1.905766e-43, 9.52883e-44, 
    1.568053e-41, 1.042566e-42, 1.884194e-39, 2.502087e-38, 2.457097e-35, 
    1.256787e-33, 5.56119e-32, 2.773154e-31, 4.486484e-31, 5.4801e-31 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 4.129627e-42, 4.203895e-44, 
    2.83021e-39, 2.054304e-42, 1.136771e-38, 2.314201e-39, 2.55329e-37, 
    6.8116e-38, 2.123633e-35, 4.665767e-37, 3.559851e-34, 8.672164e-36, 
    1.569547e-35, 4.101116e-37, 0, 1.401298e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2.354181e-43, 1.261169e-44, 4.230506e-40, 2.467126e-41, 
    7.200734e-38, 1.034653e-38, 6.580546e-38, 3.770708e-38, 6.628295e-38, 
    3.783591e-39, 1.305333e-38, 1.006581e-39, 2.242078e-44, 5.927493e-43, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.3887e-44, 1.639519e-42, 7.438947e-40, 
    2.538186e-40, 1.556882e-39, 8.5098e-39, 1.371429e-37, 8.732142e-38, 
    2.907517e-37, 1.484316e-39, 5.133721e-38, 1.368046e-40, 7.200222e-40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.937996e-42, 8.407791e-45, 
    6.992074e-39, 3.16814e-40, 1.444862e-38, 2.099448e-39, 5.577157e-38, 
    2.93066e-39, 4.528757e-37, 1.305651e-36, 6.342233e-37, 9.807913e-36, 
    2.481914e-39, 6.581614e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.942727e-44, 8.229826e-42, 3.884483e-40, 4.713947e-39, 1.028449e-39, 
    3.949331e-39, 8.76494e-40, 4.290271e-40, 8.795685e-37, 1.320532e-38, 
    6.652725e-36, 4.771931e-36, 2.991472e-37, 4.954296e-36, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.541428e-44, 2.808202e-42, 2.134682e-40, 9.383546e-39, 
    7.150036e-39, 7.869013e-39, 1.796271e-38, 2.292652e-39, 2.506942e-38, 
    3.722192e-38, 1.319574e-38, 4.563781e-36, 8.955444e-37, 4.738273e-36, 
    1.647982e-36, 0, 0, 0, 0, 0, 0, 0, 2.662467e-43, 1.401298e-44, 
    1.44614e-42, 2.242078e-44, 4.904545e-44, 1.677354e-42, 2.942727e-44, 
    1.690484e-40, 5.128752e-43, 1.854526e-38, 7.621242e-41, 2.588036e-38, 
    9.234442e-39, 5.052122e-38, 2.250775e-37, 1.420037e-36, 3.821101e-35, 
    1.804386e-35, 2.619294e-34, 0, 0, 0, 0, 1.401298e-45, 4.203895e-44, 
    9.881957e-42, 1.318622e-42, 5.150753e-41, 1.05728e-40, 3.979688e-43, 
    1.274481e-41, 0, 1.401298e-45, 0, 0, 2.106152e-42, 2.802597e-45, 
    4.134783e-40, 1.458471e-41, 1.821954e-37, 1.893859e-39, 1.190229e-35, 
    3.817268e-34, 8.652934e-33, 2.811335e-31, 0, 0, 0, 1.121039e-44, 
    2.81661e-43, 1.794783e-41, 2.717258e-41, 5.782178e-41, 3.974405e-40, 
    1.949091e-39, 7.334957e-41, 2.890849e-39, 1.401298e-45, 3.668599e-42, 0, 
    0, 8.407791e-45, 2.802597e-45, 1.045369e-42, 4.021727e-42, 7.962879e-40, 
    5.369075e-41, 1.646209e-34, 3.076976e-37, 3.536709e-30, 5.406046e-32, 0, 
    0, 8.267661e-44, 2.802597e-45, 2.35278e-41, 1.84282e-40, 9.497917e-40, 
    7.408381e-39, 9.219309e-39, 3.035903e-38, 4.269769e-39, 2.811539e-38, 
    1.810337e-41, 5.198369e-40, 3.783506e-44, 4.259947e-43, 1.415311e-43, 
    4.203895e-44, 1.717992e-42, 7.731524e-41, 8.367854e-41, 2.744555e-40, 
    7.19938e-39, 2.434756e-41, 3.576285e-34, 1.970305e-38, 1.401298e-45, 
    3.363116e-44, 5.745324e-44, 1.401298e-44, 1.502304e-40, 5.727107e-42, 
    2.949332e-38, 3.166862e-39, 1.190024e-37, 2.000895e-38, 1.53441e-38, 
    1.45978e-39, 3.269075e-40, 6.670181e-42, 2.494311e-43, 1.681558e-44, 
    3.222986e-44, 5.969531e-43, 9.709597e-41, 9.405829e-39, 3.523145e-39, 
    9.081748e-38, 1.272099e-41, 5.846974e-40, 1.357003e-40, 5.828806e-39, 
    1.249958e-42, 1.748155e-39, 1.793662e-43, 4.161856e-43, 5.361368e-42, 
    7.540359e-40, 2.173107e-39, 6.643493e-39, 3.338889e-39, 1.100972e-40, 
    6.21658e-41, 5.041872e-42, 2.491509e-42, 3.461207e-43, 6.586103e-44, 
    2.998779e-43, 1.447541e-42, 1.102317e-40, 4.636986e-39, 2.298896e-37, 
    5.816491e-37, 4.256155e-35, 1.316171e-36, 3.764968e-34, 3.156884e-36, 
    1.032073e-32, 2.613105e-39, 2.727476e-36, 6.012972e-42, 2.686009e-41, 
    3.798121e-40, 1.248526e-37, 5.728718e-39, 2.081652e-37, 6.078132e-41, 
    6.600116e-43, 1.975831e-43, 1.961818e-44, 2.073922e-43, 1.723597e-43, 
    1.544231e-42, 7.665103e-43, 1.26861e-40, 8.438619e-42, 1.524425e-38, 
    2.024336e-37, 1.987936e-34, 1.016815e-32, 4.499332e-31, 2.243645e-30, 
    3.629831e-30, 4.433725e-30,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.121039e-44, 0, 7.557203e-42, 
    5.605194e-45, 3.035493e-41, 6.179726e-42, 6.818074e-40, 1.818913e-40, 
    5.670758e-38, 1.245904e-39, 9.505908e-37, 2.315736e-38, 4.191177e-38, 
    1.095125e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.129447e-42, 6.586103e-44, 1.92282e-40, 2.7628e-41, 1.757214e-40, 
    1.006889e-40, 1.769966e-40, 1.010336e-41, 3.48559e-41, 2.68769e-42, 0, 
    1.401298e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.203895e-45, 
    1.987041e-42, 6.782285e-43, 4.157653e-42, 2.272346e-41, 3.662139e-40, 
    2.331747e-40, 7.763964e-40, 3.964273e-42, 1.370862e-40, 3.657389e-43, 
    1.922581e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.605194e-45, 0, 
    1.86709e-41, 8.463843e-43, 3.858195e-41, 5.606595e-42, 1.489272e-40, 
    7.826252e-42, 1.209318e-39, 3.486492e-39, 1.693573e-39, 2.619017e-38, 
    6.628142e-42, 1.757495e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.242078e-44, 1.036961e-42, 1.258786e-41, 2.746545e-42, 1.054617e-41, 
    2.340168e-42, 1.146262e-42, 2.348721e-39, 3.526227e-41, 1.776484e-38, 
    1.274254e-38, 7.988158e-40, 1.322951e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7.006492e-45, 5.703285e-43, 2.505662e-41, 1.909269e-41, 
    2.101247e-41, 4.796645e-41, 6.122273e-42, 6.694283e-41, 9.93941e-41, 
    3.523705e-41, 1.218671e-38, 2.39138e-39, 1.265266e-38, 4.400621e-39, 0, 
    0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 4.203895e-45, 0, 0, 4.203895e-45, 0, 
    4.512181e-43, 1.401298e-45, 4.952189e-41, 2.031883e-43, 6.910784e-41, 
    2.465865e-41, 1.349072e-40, 6.010267e-40, 3.791939e-39, 1.020352e-37, 
    4.818269e-38, 6.994329e-37, 0, 0, 0, 0, 0, 0, 2.662467e-44, 4.203895e-45, 
    1.373272e-43, 2.81661e-43, 1.401298e-45, 3.363116e-44, 0, 0, 0, 0, 
    5.605194e-45, 0, 1.104223e-42, 3.923636e-44, 4.865182e-40, 5.057286e-42, 
    3.178282e-38, 1.019329e-36, 2.310603e-35, 7.507139e-34, 0, 0, 0, 0, 
    1.401298e-45, 4.764415e-44, 7.286752e-44, 1.541428e-43, 1.060783e-42, 
    5.204422e-42, 1.961818e-43, 7.719753e-42, 0, 9.809089e-45, 0, 0, 0, 0, 
    2.802597e-45, 1.121039e-44, 2.12577e-42, 1.429324e-43, 4.39589e-37, 
    8.216472e-40, 9.444112e-33, 1.443582e-34, 0, 0, 0, 0, 6.305843e-44, 
    4.918558e-43, 2.53635e-42, 1.978213e-41, 2.461801e-41, 8.106792e-41, 
    1.140096e-41, 7.507737e-41, 4.764415e-44, 1.388687e-42, 0, 1.401298e-45, 
    0, 0, 4.203895e-45, 2.059909e-43, 2.228065e-43, 7.328791e-43, 
    1.922441e-41, 6.445973e-44, 9.549791e-37, 5.261315e-41, 0, 0, 0, 0, 
    4.007714e-43, 1.541428e-44, 7.875578e-41, 8.456836e-42, 3.177739e-40, 
    5.343011e-41, 4.097397e-41, 3.898412e-42, 8.730089e-43, 1.821688e-44, 0, 
    0, 0, 1.401298e-45, 2.592402e-43, 2.511687e-41, 9.408318e-42, 
    2.425101e-40, 3.363116e-44, 1.561046e-42, 3.629363e-43, 1.556422e-41, 
    2.802597e-45, 4.667725e-42, 0, 1.401298e-45, 1.401298e-44, 2.013666e-42, 
    5.802777e-42, 1.774044e-41, 8.916462e-42, 2.942727e-43, 1.653532e-43, 
    1.401298e-44, 7.006492e-45, 1.401298e-45, 0, 1.401298e-45, 4.203895e-45, 
    2.942727e-43, 1.238187e-41, 6.138766e-40, 1.553182e-39, 1.136525e-37, 
    3.514583e-39, 1.005363e-36, 8.429858e-39, 2.755955e-35, 6.978466e-42, 
    7.283205e-39, 1.541428e-44, 7.146622e-44, 1.01454e-42, 3.333955e-40, 
    1.529798e-41, 5.558657e-40, 1.625506e-43, 1.401298e-45, 0, 0, 0, 0, 
    4.203895e-45, 1.401298e-45, 3.391142e-43, 2.242078e-44, 4.070632e-41, 
    5.405607e-40, 5.308407e-37, 2.715213e-35, 1.201461e-33, 5.99123e-33, 
    9.692775e-33, 1.183942e-32 ;

 F_N2O_NIT =
  2.302583e-14, 2.322413e-14, 2.31855e-14, 2.334595e-14, 2.325687e-14, 
    2.336203e-14, 2.306595e-14, 2.323199e-14, 2.312592e-14, 2.304362e-14, 
    2.365893e-14, 2.33531e-14, 2.397887e-14, 2.378218e-14, 2.427788e-14, 
    2.394819e-14, 2.434465e-14, 2.426834e-14, 2.449839e-14, 2.443236e-14, 
    2.472783e-14, 2.452888e-14, 2.488173e-14, 2.468024e-14, 2.471169e-14, 
    2.452232e-14, 2.341451e-14, 2.362076e-14, 2.340231e-14, 2.343166e-14, 
    2.341848e-14, 2.32587e-14, 2.317838e-14, 2.301069e-14, 2.304108e-14, 
    2.316428e-14, 2.344484e-14, 2.33494e-14, 2.359032e-14, 2.358487e-14, 
    2.385456e-14, 2.373276e-14, 2.418848e-14, 2.405849e-14, 2.443511e-14, 
    2.43401e-14, 2.443064e-14, 2.440316e-14, 2.443099e-14, 2.429173e-14, 
    2.435134e-14, 2.422899e-14, 2.375558e-14, 2.389421e-14, 2.348197e-14, 
    2.323588e-14, 2.30732e-14, 2.295812e-14, 2.297437e-14, 2.300536e-14, 
    2.316499e-14, 2.331561e-14, 2.343073e-14, 2.35079e-14, 2.358407e-14, 
    2.38154e-14, 2.393834e-14, 2.421479e-14, 2.416479e-14, 2.424954e-14, 
    2.433066e-14, 2.446716e-14, 2.444467e-14, 2.45049e-14, 2.424729e-14, 
    2.441833e-14, 2.41363e-14, 2.421327e-14, 2.36048e-14, 2.337514e-14, 
    2.327786e-14, 2.31929e-14, 2.298686e-14, 2.312904e-14, 2.307293e-14, 
    2.320652e-14, 2.329162e-14, 2.324951e-14, 2.351001e-14, 2.340855e-14, 
    2.394563e-14, 2.371351e-14, 2.432119e-14, 2.417504e-14, 2.435628e-14, 
    2.426371e-14, 2.442243e-14, 2.427956e-14, 2.452734e-14, 2.458146e-14, 
    2.454446e-14, 2.468675e-14, 2.427163e-14, 2.443061e-14, 2.324834e-14, 
    2.325521e-14, 2.32872e-14, 2.314672e-14, 2.313814e-14, 2.300984e-14, 
    2.312398e-14, 2.317268e-14, 2.329655e-14, 2.336997e-14, 2.343988e-14, 
    2.359399e-14, 2.376672e-14, 2.400936e-14, 2.41845e-14, 2.430226e-14, 
    2.423001e-14, 2.429378e-14, 2.422249e-14, 2.418911e-14, 2.456117e-14, 
    2.435188e-14, 2.466625e-14, 2.46488e-14, 2.450631e-14, 2.465076e-14, 
    2.326002e-14, 2.322053e-14, 2.308368e-14, 2.319074e-14, 2.299588e-14, 
    2.310484e-14, 2.316761e-14, 2.341065e-14, 2.346424e-14, 2.351398e-14, 
    2.361237e-14, 2.373896e-14, 2.39619e-14, 2.415676e-14, 2.433537e-14, 
    2.432226e-14, 2.432687e-14, 2.436685e-14, 2.426786e-14, 2.438312e-14, 
    2.440248e-14, 2.435185e-14, 2.464645e-14, 2.45621e-14, 2.464842e-14, 
    2.459347e-14, 2.323336e-14, 2.329984e-14, 2.32639e-14, 2.33315e-14, 
    2.328386e-14, 2.349608e-14, 2.35599e-14, 2.385977e-14, 2.373647e-14, 
    2.393287e-14, 2.375638e-14, 2.37876e-14, 2.393927e-14, 2.376589e-14, 
    2.414598e-14, 2.388793e-14, 2.43684e-14, 2.410946e-14, 2.438467e-14, 
    2.433458e-14, 2.441754e-14, 2.449197e-14, 2.458578e-14, 2.475937e-14, 
    2.471911e-14, 2.486465e-14, 2.339914e-14, 2.348572e-14, 2.347809e-14, 
    2.356886e-14, 2.36361e-14, 2.378221e-14, 2.401752e-14, 2.392888e-14, 
    2.409173e-14, 2.412449e-14, 2.387713e-14, 2.402884e-14, 2.354373e-14, 
    2.362174e-14, 2.357527e-14, 2.340592e-14, 2.394926e-14, 2.366959e-14, 
    2.418736e-14, 2.403485e-14, 2.448134e-14, 2.425875e-14, 2.469696e-14, 
    2.488553e-14, 2.506373e-14, 2.527277e-14, 2.353304e-14, 2.347413e-14, 
    2.357966e-14, 2.372607e-14, 2.386236e-14, 2.404417e-14, 2.406282e-14, 
    2.409696e-14, 2.418555e-14, 2.426017e-14, 2.410776e-14, 2.427889e-14, 
    2.363984e-14, 2.397362e-14, 2.345184e-14, 2.360831e-14, 2.371739e-14, 
    2.366951e-14, 2.391873e-14, 2.397766e-14, 2.421793e-14, 2.409357e-14, 
    2.483891e-14, 2.450768e-14, 2.543257e-14, 2.517229e-14, 2.345356e-14, 
    2.353283e-14, 2.38098e-14, 2.367781e-14, 2.405633e-14, 2.414999e-14, 
    2.422626e-14, 2.432394e-14, 2.43345e-14, 2.439249e-14, 2.42975e-14, 
    2.438873e-14, 2.404453e-14, 2.419803e-14, 2.377803e-14, 2.387989e-14, 
    2.383301e-14, 2.378162e-14, 2.394038e-14, 2.411012e-14, 2.411376e-14, 
    2.416832e-14, 2.43224e-14, 2.405782e-14, 2.48818e-14, 2.437119e-14, 
    2.361943e-14, 2.377279e-14, 2.379475e-14, 2.373524e-14, 2.414058e-14, 
    2.399329e-14, 2.439107e-14, 2.428323e-14, 2.446006e-14, 2.43721e-14, 
    2.435917e-14, 2.424648e-14, 2.417645e-14, 2.400001e-14, 2.385695e-14, 
    2.374384e-14, 2.377011e-14, 2.389445e-14, 2.412052e-14, 2.433542e-14, 
    2.428825e-14, 2.444656e-14, 2.402872e-14, 2.420346e-14, 2.413584e-14, 
    2.431236e-14, 2.392652e-14, 2.42549e-14, 2.384295e-14, 2.387892e-14, 
    2.399037e-14, 2.421537e-14, 2.426531e-14, 2.431868e-14, 2.428574e-14, 
    2.412629e-14, 2.410022e-14, 2.398764e-14, 2.395659e-14, 2.387106e-14, 
    2.380035e-14, 2.386494e-14, 2.393286e-14, 2.412634e-14, 2.430139e-14, 
    2.4493e-14, 2.454001e-14, 2.476509e-14, 2.458177e-14, 2.488464e-14, 
    2.462699e-14, 2.50739e-14, 2.427401e-14, 2.461951e-14, 2.399545e-14, 
    2.406227e-14, 2.418339e-14, 2.446239e-14, 2.431157e-14, 2.448801e-14, 
    2.40992e-14, 2.389875e-14, 2.384704e-14, 2.37507e-14, 2.384923e-14, 
    2.384121e-14, 2.393568e-14, 2.39053e-14, 2.413277e-14, 2.401044e-14, 
    2.43588e-14, 2.448658e-14, 2.484934e-14, 2.507309e-14, 2.530196e-14, 
    2.540334e-14, 2.543424e-14, 2.544716e-14 ;

 F_NIT =
  3.837638e-11, 3.870687e-11, 3.864251e-11, 3.890991e-11, 3.876146e-11, 
    3.893671e-11, 3.844325e-11, 3.871999e-11, 3.85432e-11, 3.840604e-11, 
    3.943156e-11, 3.892183e-11, 3.996478e-11, 3.963697e-11, 4.046314e-11, 
    3.991366e-11, 4.057441e-11, 4.044724e-11, 4.083065e-11, 4.072061e-11, 
    4.121304e-11, 4.088148e-11, 4.146955e-11, 4.113373e-11, 4.118616e-11, 
    4.087053e-11, 3.902418e-11, 3.936794e-11, 3.900385e-11, 3.905276e-11, 
    3.903081e-11, 3.87645e-11, 3.863064e-11, 3.835115e-11, 3.84018e-11, 
    3.860712e-11, 3.907473e-11, 3.891567e-11, 3.93172e-11, 3.930811e-11, 
    3.97576e-11, 3.95546e-11, 4.031413e-11, 4.009748e-11, 4.072519e-11, 
    4.056684e-11, 4.071773e-11, 4.067194e-11, 4.071832e-11, 4.048622e-11, 
    4.058556e-11, 4.038165e-11, 3.959263e-11, 3.982369e-11, 3.913661e-11, 
    3.872647e-11, 3.845534e-11, 3.826354e-11, 3.829061e-11, 3.834227e-11, 
    3.860832e-11, 3.885935e-11, 3.905122e-11, 3.917984e-11, 3.930679e-11, 
    3.969234e-11, 3.989723e-11, 4.035799e-11, 4.027464e-11, 4.041589e-11, 
    4.05511e-11, 4.077861e-11, 4.074111e-11, 4.08415e-11, 4.041215e-11, 
    4.069722e-11, 4.022717e-11, 4.035544e-11, 3.934133e-11, 3.895857e-11, 
    3.879643e-11, 3.865483e-11, 3.831144e-11, 3.85484e-11, 3.845489e-11, 
    3.867754e-11, 3.881936e-11, 3.874918e-11, 3.918335e-11, 3.901425e-11, 
    3.990938e-11, 3.952251e-11, 4.053532e-11, 4.029174e-11, 4.059381e-11, 
    4.043952e-11, 4.070406e-11, 4.046593e-11, 4.087889e-11, 4.096911e-11, 
    4.090744e-11, 4.114458e-11, 4.045272e-11, 4.071768e-11, 3.874724e-11, 
    3.875868e-11, 3.8812e-11, 3.857787e-11, 3.856357e-11, 3.834973e-11, 
    3.853997e-11, 3.862113e-11, 3.882758e-11, 3.894995e-11, 3.906647e-11, 
    3.932332e-11, 3.96112e-11, 4.001561e-11, 4.030749e-11, 4.050376e-11, 
    4.038335e-11, 4.048964e-11, 4.037082e-11, 4.031519e-11, 4.093528e-11, 
    4.058647e-11, 4.111041e-11, 4.108133e-11, 4.084385e-11, 4.108459e-11, 
    3.87667e-11, 3.870088e-11, 3.847281e-11, 3.865122e-11, 3.832647e-11, 
    3.850806e-11, 3.861268e-11, 3.901776e-11, 3.910706e-11, 3.918996e-11, 
    3.935395e-11, 3.956494e-11, 3.99365e-11, 4.026126e-11, 4.055896e-11, 
    4.053709e-11, 4.054479e-11, 4.061142e-11, 4.044644e-11, 4.063853e-11, 
    4.06708e-11, 4.058642e-11, 4.107742e-11, 4.093683e-11, 4.108069e-11, 
    4.098911e-11, 3.872226e-11, 3.883307e-11, 3.877316e-11, 3.888584e-11, 
    3.880643e-11, 3.916014e-11, 3.926651e-11, 3.976628e-11, 3.956078e-11, 
    3.988811e-11, 3.959396e-11, 3.964599e-11, 3.989878e-11, 3.960982e-11, 
    4.024329e-11, 3.981321e-11, 4.061401e-11, 4.018243e-11, 4.064112e-11, 
    4.055763e-11, 4.06959e-11, 4.081996e-11, 4.09763e-11, 4.126561e-11, 
    4.119851e-11, 4.144108e-11, 3.899858e-11, 3.914286e-11, 3.913015e-11, 
    3.928143e-11, 3.93935e-11, 3.963701e-11, 4.00292e-11, 3.988147e-11, 
    4.015288e-11, 4.020748e-11, 3.979522e-11, 4.004806e-11, 3.923955e-11, 
    3.936957e-11, 3.929213e-11, 3.900987e-11, 3.991543e-11, 3.944932e-11, 
    4.031227e-11, 4.005809e-11, 4.080224e-11, 4.043125e-11, 4.11616e-11, 
    4.147589e-11, 4.177288e-11, 4.212129e-11, 3.922173e-11, 3.912355e-11, 
    3.929944e-11, 3.954346e-11, 3.97706e-11, 4.007362e-11, 4.010469e-11, 
    4.016161e-11, 4.030926e-11, 4.043362e-11, 4.017959e-11, 4.046481e-11, 
    3.939973e-11, 3.995603e-11, 3.908639e-11, 3.934719e-11, 3.952899e-11, 
    3.944919e-11, 3.986455e-11, 3.996277e-11, 4.036321e-11, 4.015595e-11, 
    4.139818e-11, 4.084614e-11, 4.238762e-11, 4.195382e-11, 3.908927e-11, 
    3.922138e-11, 3.968301e-11, 3.946301e-11, 4.009388e-11, 4.024997e-11, 
    4.03771e-11, 4.05399e-11, 4.05575e-11, 4.065415e-11, 4.049583e-11, 
    4.064788e-11, 4.007421e-11, 4.033004e-11, 3.963006e-11, 3.979982e-11, 
    3.972167e-11, 3.963604e-11, 3.990063e-11, 4.018353e-11, 4.018959e-11, 
    4.028053e-11, 4.053733e-11, 4.009636e-11, 4.146967e-11, 4.061865e-11, 
    3.936571e-11, 3.962132e-11, 3.965791e-11, 3.955874e-11, 4.02343e-11, 
    3.998882e-11, 4.065179e-11, 4.047205e-11, 4.076676e-11, 4.062017e-11, 
    4.059861e-11, 4.04108e-11, 4.029408e-11, 4.000002e-11, 3.976158e-11, 
    3.957306e-11, 3.961685e-11, 3.982409e-11, 4.020086e-11, 4.055902e-11, 
    4.048042e-11, 4.074426e-11, 4.004787e-11, 4.03391e-11, 4.02264e-11, 
    4.05206e-11, 3.987753e-11, 4.042483e-11, 3.973825e-11, 3.97982e-11, 
    3.998394e-11, 4.035896e-11, 4.044219e-11, 4.053113e-11, 4.047623e-11, 
    4.021049e-11, 4.016704e-11, 3.997939e-11, 3.992765e-11, 3.97851e-11, 
    3.966726e-11, 3.97749e-11, 3.98881e-11, 4.021057e-11, 4.050232e-11, 
    4.082166e-11, 4.090002e-11, 4.127515e-11, 4.096961e-11, 4.147441e-11, 
    4.104499e-11, 4.178983e-11, 4.045668e-11, 4.103252e-11, 3.999241e-11, 
    4.010379e-11, 4.030565e-11, 4.077065e-11, 4.051928e-11, 4.081335e-11, 
    4.016533e-11, 3.983125e-11, 3.974506e-11, 3.95845e-11, 3.974873e-11, 
    3.973535e-11, 3.989281e-11, 3.984217e-11, 4.022128e-11, 4.00174e-11, 
    4.0598e-11, 4.081097e-11, 4.141557e-11, 4.178849e-11, 4.216993e-11, 
    4.23389e-11, 4.23904e-11, 4.241194e-11 ;

 F_NIT_vr =
  2.454741e-10, 2.465639e-10, 2.463515e-10, 2.47231e-10, 2.467428e-10, 
    2.473182e-10, 2.456938e-10, 2.466052e-10, 2.46023e-10, 2.455701e-10, 
    2.489369e-10, 2.472681e-10, 2.506745e-10, 2.496075e-10, 2.52289e-10, 
    2.505075e-10, 2.526483e-10, 2.522372e-10, 2.534745e-10, 2.531195e-10, 
    2.547023e-10, 2.536375e-10, 2.55524e-10, 2.544477e-10, 2.546155e-10, 
    2.53601e-10, 2.47606e-10, 2.487309e-10, 2.475388e-10, 2.476992e-10, 
    2.47627e-10, 2.467516e-10, 2.463107e-10, 2.453887e-10, 2.455557e-10, 
    2.462327e-10, 2.477693e-10, 2.472472e-10, 2.48563e-10, 2.485333e-10, 
    2.499995e-10, 2.49338e-10, 2.518062e-10, 2.511037e-10, 2.53134e-10, 
    2.526225e-10, 2.531093e-10, 2.529613e-10, 2.531105e-10, 2.523612e-10, 
    2.526816e-10, 2.520227e-10, 2.49465e-10, 2.502172e-10, 2.479736e-10, 
    2.466259e-10, 2.457326e-10, 2.450992e-10, 2.451881e-10, 2.453588e-10, 
    2.462361e-10, 2.47062e-10, 2.476919e-10, 2.48113e-10, 2.485283e-10, 
    2.497862e-10, 2.504531e-10, 2.519475e-10, 2.516778e-10, 2.521343e-10, 
    2.525714e-10, 2.53305e-10, 2.531841e-10, 2.53507e-10, 2.521211e-10, 
    2.530417e-10, 2.515218e-10, 2.519372e-10, 2.486426e-10, 2.473892e-10, 
    2.468558e-10, 2.463899e-10, 2.452567e-10, 2.460389e-10, 2.457301e-10, 
    2.464638e-10, 2.469303e-10, 2.466991e-10, 2.481242e-10, 2.475694e-10, 
    2.504922e-10, 2.492322e-10, 2.525208e-10, 2.517325e-10, 2.52709e-10, 
    2.522106e-10, 2.530641e-10, 2.522954e-10, 2.53627e-10, 2.539171e-10, 
    2.537182e-10, 2.544807e-10, 2.522511e-10, 2.531065e-10, 2.466942e-10, 
    2.467318e-10, 2.469069e-10, 2.461356e-10, 2.460884e-10, 2.453824e-10, 
    2.4601e-10, 2.462774e-10, 2.469567e-10, 2.473582e-10, 2.477402e-10, 
    2.485814e-10, 2.49521e-10, 2.508367e-10, 2.517833e-10, 2.524178e-10, 
    2.520284e-10, 2.523717e-10, 2.519873e-10, 2.518069e-10, 2.538076e-10, 
    2.526835e-10, 2.543702e-10, 2.542769e-10, 2.535125e-10, 2.542866e-10, 
    2.467577e-10, 2.465408e-10, 2.457889e-10, 2.463768e-10, 2.453051e-10, 
    2.459045e-10, 2.462489e-10, 2.475804e-10, 2.478732e-10, 2.481448e-10, 
    2.486811e-10, 2.493698e-10, 2.505794e-10, 2.516329e-10, 2.525958e-10, 
    2.525248e-10, 2.525495e-10, 2.527642e-10, 2.522312e-10, 2.528512e-10, 
    2.529549e-10, 2.526828e-10, 2.542636e-10, 2.538116e-10, 2.542738e-10, 
    2.539791e-10, 2.466109e-10, 2.469749e-10, 2.467776e-10, 2.47148e-10, 
    2.468864e-10, 2.480471e-10, 2.48395e-10, 2.50026e-10, 2.493561e-10, 
    2.504222e-10, 2.494639e-10, 2.496336e-10, 2.504556e-10, 2.49515e-10, 
    2.515736e-10, 2.501765e-10, 2.527723e-10, 2.513752e-10, 2.528593e-10, 
    2.525894e-10, 2.530354e-10, 2.534351e-10, 2.539378e-10, 2.548667e-10, 
    2.54651e-10, 2.554285e-10, 2.475182e-10, 2.479908e-10, 2.479492e-10, 
    2.484442e-10, 2.488103e-10, 2.496053e-10, 2.508808e-10, 2.504005e-10, 
    2.512816e-10, 2.514585e-10, 2.501191e-10, 2.509408e-10, 2.483048e-10, 
    2.487295e-10, 2.484765e-10, 2.475512e-10, 2.505084e-10, 2.489892e-10, 
    2.517956e-10, 2.509712e-10, 2.533773e-10, 2.521797e-10, 2.545324e-10, 
    2.555392e-10, 2.564882e-10, 2.575969e-10, 2.482489e-10, 2.47927e-10, 
    2.485026e-10, 2.492996e-10, 2.500396e-10, 2.510247e-10, 2.511253e-10, 
    2.513094e-10, 2.517876e-10, 2.5219e-10, 2.513669e-10, 2.522902e-10, 
    2.488273e-10, 2.506404e-10, 2.478018e-10, 2.486554e-10, 2.492489e-10, 
    2.489886e-10, 2.503422e-10, 2.506611e-10, 2.51959e-10, 2.512879e-10, 
    2.552896e-10, 2.535172e-10, 2.584422e-10, 2.570637e-10, 2.478144e-10, 
    2.482468e-10, 2.49754e-10, 2.490366e-10, 2.510898e-10, 2.515959e-10, 
    2.52007e-10, 2.525332e-10, 2.525896e-10, 2.529016e-10, 2.523899e-10, 
    2.528809e-10, 2.510238e-10, 2.518532e-10, 2.495789e-10, 2.501314e-10, 
    2.49877e-10, 2.495975e-10, 2.504586e-10, 2.513768e-10, 2.513964e-10, 
    2.516905e-10, 2.525199e-10, 2.510931e-10, 2.555168e-10, 2.527817e-10, 
    2.487187e-10, 2.495524e-10, 2.496717e-10, 2.493485e-10, 2.515443e-10, 
    2.50748e-10, 2.52894e-10, 2.523132e-10, 2.532641e-10, 2.527913e-10, 
    2.527211e-10, 2.521144e-10, 2.51736e-10, 2.507823e-10, 2.500064e-10, 
    2.493922e-10, 2.495344e-10, 2.502093e-10, 2.514322e-10, 2.525913e-10, 
    2.523369e-10, 2.531884e-10, 2.509352e-10, 2.518792e-10, 2.515135e-10, 
    2.524657e-10, 2.503865e-10, 2.521605e-10, 2.499331e-10, 2.501279e-10, 
    2.507314e-10, 2.51947e-10, 2.522161e-10, 2.525035e-10, 2.523257e-10, 
    2.514654e-10, 2.513243e-10, 2.50715e-10, 2.505464e-10, 2.50083e-10, 
    2.496986e-10, 2.500492e-10, 2.504168e-10, 2.514638e-10, 2.524075e-10, 
    2.534374e-10, 2.536897e-10, 2.548935e-10, 2.539125e-10, 2.555306e-10, 
    2.541534e-10, 2.565381e-10, 2.522632e-10, 2.541193e-10, 2.507591e-10, 
    2.511203e-10, 2.51774e-10, 2.532756e-10, 2.524646e-10, 2.53413e-10, 
    2.513187e-10, 2.502329e-10, 2.499523e-10, 2.494291e-10, 2.499638e-10, 
    2.499203e-10, 2.504324e-10, 2.502673e-10, 2.514978e-10, 2.508365e-10, 
    2.527157e-10, 2.534024e-10, 2.553437e-10, 2.565348e-10, 2.577494e-10, 
    2.582854e-10, 2.584487e-10, 2.585166e-10,
  1.247084e-10, 1.256584e-10, 1.254736e-10, 1.262413e-10, 1.258153e-10, 
    1.263183e-10, 1.249009e-10, 1.256961e-10, 1.251883e-10, 1.247939e-10, 
    1.277361e-10, 1.262756e-10, 1.292607e-10, 1.283242e-10, 1.306818e-10, 
    1.291147e-10, 1.309987e-10, 1.306367e-10, 1.317279e-10, 1.31415e-10, 
    1.328139e-10, 1.318724e-10, 1.335415e-10, 1.325889e-10, 1.327377e-10, 
    1.318414e-10, 1.265692e-10, 1.275538e-10, 1.265109e-10, 1.266511e-10, 
    1.265883e-10, 1.25824e-10, 1.254394e-10, 1.24636e-10, 1.247818e-10, 
    1.25372e-10, 1.267142e-10, 1.262581e-10, 1.274092e-10, 1.273832e-10, 
    1.286691e-10, 1.280887e-10, 1.302575e-10, 1.296397e-10, 1.31428e-10, 
    1.309774e-10, 1.314068e-10, 1.312766e-10, 1.314085e-10, 1.307479e-10, 
    1.310308e-10, 1.3045e-10, 1.281973e-10, 1.288577e-10, 1.268916e-10, 
    1.257146e-10, 1.249357e-10, 1.243839e-10, 1.244619e-10, 1.246105e-10, 
    1.253754e-10, 1.260965e-10, 1.26647e-10, 1.270157e-10, 1.273794e-10, 
    1.284823e-10, 1.290679e-10, 1.303824e-10, 1.30145e-10, 1.305475e-10, 
    1.309326e-10, 1.3158e-10, 1.314734e-10, 1.317588e-10, 1.30537e-10, 
    1.313485e-10, 1.300098e-10, 1.303754e-10, 1.274777e-10, 1.263811e-10, 
    1.259155e-10, 1.255091e-10, 1.245218e-10, 1.252032e-10, 1.249344e-10, 
    1.255745e-10, 1.259817e-10, 1.257802e-10, 1.270258e-10, 1.26541e-10, 
    1.291026e-10, 1.279968e-10, 1.308877e-10, 1.301937e-10, 1.310542e-10, 
    1.306149e-10, 1.313679e-10, 1.306902e-10, 1.318652e-10, 1.321215e-10, 
    1.319463e-10, 1.326199e-10, 1.306526e-10, 1.314067e-10, 1.257746e-10, 
    1.258074e-10, 1.259605e-10, 1.252879e-10, 1.252469e-10, 1.24632e-10, 
    1.251791e-10, 1.254123e-10, 1.260054e-10, 1.263565e-10, 1.266907e-10, 
    1.274267e-10, 1.282505e-10, 1.29406e-10, 1.302387e-10, 1.307979e-10, 
    1.304549e-10, 1.307577e-10, 1.304192e-10, 1.302607e-10, 1.320254e-10, 
    1.310334e-10, 1.32523e-10, 1.324404e-10, 1.317656e-10, 1.324497e-10, 
    1.258305e-10, 1.256415e-10, 1.24986e-10, 1.254989e-10, 1.245651e-10, 
    1.250874e-10, 1.25388e-10, 1.265509e-10, 1.268072e-10, 1.270447e-10, 
    1.275145e-10, 1.281184e-10, 1.291802e-10, 1.301069e-10, 1.309551e-10, 
    1.308929e-10, 1.309148e-10, 1.311044e-10, 1.306347e-10, 1.311816e-10, 
    1.312734e-10, 1.310333e-10, 1.324293e-10, 1.320299e-10, 1.324386e-10, 
    1.321786e-10, 1.257029e-10, 1.260211e-10, 1.258491e-10, 1.261725e-10, 
    1.259446e-10, 1.269591e-10, 1.272639e-10, 1.286939e-10, 1.281064e-10, 
    1.29042e-10, 1.282014e-10, 1.283501e-10, 1.290723e-10, 1.282468e-10, 
    1.300556e-10, 1.28828e-10, 1.311118e-10, 1.298819e-10, 1.31189e-10, 
    1.309514e-10, 1.313449e-10, 1.316977e-10, 1.321421e-10, 1.329634e-10, 
    1.327731e-10, 1.334611e-10, 1.26496e-10, 1.269096e-10, 1.268733e-10, 
    1.273068e-10, 1.276277e-10, 1.283245e-10, 1.294449e-10, 1.290232e-10, 
    1.297979e-10, 1.299536e-10, 1.287768e-10, 1.294987e-10, 1.271869e-10, 
    1.275592e-10, 1.273375e-10, 1.265286e-10, 1.291201e-10, 1.277875e-10, 
    1.302524e-10, 1.295275e-10, 1.316474e-10, 1.305914e-10, 1.326683e-10, 
    1.335596e-10, 1.344009e-10, 1.353859e-10, 1.271358e-10, 1.268544e-10, 
    1.273584e-10, 1.280568e-10, 1.287064e-10, 1.295717e-10, 1.296604e-10, 
    1.298228e-10, 1.302438e-10, 1.305982e-10, 1.29874e-10, 1.306871e-10, 
    1.276453e-10, 1.292361e-10, 1.26748e-10, 1.274951e-10, 1.280156e-10, 
    1.277873e-10, 1.28975e-10, 1.292555e-10, 1.303976e-10, 1.298068e-10, 
    1.333393e-10, 1.317721e-10, 1.36138e-10, 1.349127e-10, 1.267562e-10, 
    1.271348e-10, 1.284559e-10, 1.278267e-10, 1.296296e-10, 1.300748e-10, 
    1.304372e-10, 1.309008e-10, 1.30951e-10, 1.31226e-10, 1.307754e-10, 
    1.312083e-10, 1.295735e-10, 1.303031e-10, 1.283048e-10, 1.2879e-10, 
    1.285668e-10, 1.28322e-10, 1.290781e-10, 1.298853e-10, 1.299028e-10, 
    1.30162e-10, 1.308931e-10, 1.296369e-10, 1.335416e-10, 1.311247e-10, 
    1.275482e-10, 1.282795e-10, 1.283843e-10, 1.281007e-10, 1.300301e-10, 
    1.293297e-10, 1.312193e-10, 1.307077e-10, 1.315465e-10, 1.311294e-10, 
    1.310681e-10, 1.305333e-10, 1.302006e-10, 1.293618e-10, 1.286808e-10, 
    1.281419e-10, 1.282671e-10, 1.288594e-10, 1.299348e-10, 1.309554e-10, 
    1.307316e-10, 1.314826e-10, 1.294985e-10, 1.30329e-10, 1.300077e-10, 
    1.308462e-10, 1.290119e-10, 1.305726e-10, 1.28614e-10, 1.287854e-10, 
    1.293158e-10, 1.303853e-10, 1.306227e-10, 1.308759e-10, 1.307197e-10, 
    1.299622e-10, 1.298384e-10, 1.29303e-10, 1.291552e-10, 1.287481e-10, 
    1.284113e-10, 1.287189e-10, 1.290423e-10, 1.299626e-10, 1.30794e-10, 
    1.317027e-10, 1.319255e-10, 1.329903e-10, 1.32123e-10, 1.335551e-10, 
    1.323368e-10, 1.344486e-10, 1.306636e-10, 1.323014e-10, 1.293401e-10, 
    1.29658e-10, 1.302334e-10, 1.315573e-10, 1.308422e-10, 1.316788e-10, 
    1.298335e-10, 1.288797e-10, 1.286337e-10, 1.281746e-10, 1.286442e-10, 
    1.286059e-10, 1.290558e-10, 1.289112e-10, 1.299932e-10, 1.294116e-10, 
    1.310665e-10, 1.316723e-10, 1.333889e-10, 1.344451e-10, 1.355237e-10, 
    1.360008e-10, 1.361461e-10, 1.362069e-10,
  1.174451e-10, 1.184872e-10, 1.182844e-10, 1.191271e-10, 1.186593e-10, 
    1.192116e-10, 1.176561e-10, 1.185286e-10, 1.179714e-10, 1.175389e-10, 
    1.207697e-10, 1.191648e-10, 1.224471e-10, 1.214163e-10, 1.24013e-10, 
    1.222864e-10, 1.243625e-10, 1.239632e-10, 1.251668e-10, 1.248215e-10, 
    1.263661e-10, 1.253263e-10, 1.271701e-10, 1.261175e-10, 1.262819e-10, 
    1.252921e-10, 1.194871e-10, 1.205694e-10, 1.194231e-10, 1.195772e-10, 
    1.195081e-10, 1.186689e-10, 1.18247e-10, 1.173657e-10, 1.175255e-10, 
    1.181729e-10, 1.196465e-10, 1.191455e-10, 1.204101e-10, 1.203815e-10, 
    1.217958e-10, 1.211573e-10, 1.235452e-10, 1.228645e-10, 1.248359e-10, 
    1.243389e-10, 1.248125e-10, 1.246688e-10, 1.248144e-10, 1.240858e-10, 
    1.243977e-10, 1.237574e-10, 1.212767e-10, 1.220035e-10, 1.198413e-10, 
    1.18549e-10, 1.176943e-10, 1.170894e-10, 1.171748e-10, 1.173377e-10, 
    1.181767e-10, 1.18968e-10, 1.195725e-10, 1.199776e-10, 1.203773e-10, 
    1.215904e-10, 1.222349e-10, 1.236829e-10, 1.234212e-10, 1.238648e-10, 
    1.242895e-10, 1.250036e-10, 1.24886e-10, 1.25201e-10, 1.238532e-10, 
    1.247482e-10, 1.232722e-10, 1.236751e-10, 1.204857e-10, 1.192806e-10, 
    1.187695e-10, 1.183233e-10, 1.172405e-10, 1.179878e-10, 1.17693e-10, 
    1.18395e-10, 1.18842e-10, 1.186209e-10, 1.199887e-10, 1.194561e-10, 
    1.222731e-10, 1.210563e-10, 1.242399e-10, 1.234749e-10, 1.244236e-10, 
    1.239391e-10, 1.247697e-10, 1.240221e-10, 1.253184e-10, 1.256013e-10, 
    1.254079e-10, 1.261517e-10, 1.239807e-10, 1.248125e-10, 1.186146e-10, 
    1.186507e-10, 1.188188e-10, 1.180807e-10, 1.180357e-10, 1.173613e-10, 
    1.179613e-10, 1.182172e-10, 1.18868e-10, 1.192536e-10, 1.196206e-10, 
    1.204294e-10, 1.213353e-10, 1.226071e-10, 1.235244e-10, 1.241409e-10, 
    1.237628e-10, 1.240966e-10, 1.237234e-10, 1.235487e-10, 1.254952e-10, 
    1.244006e-10, 1.260446e-10, 1.259534e-10, 1.252085e-10, 1.259637e-10, 
    1.18676e-10, 1.184686e-10, 1.177495e-10, 1.183121e-10, 1.17288e-10, 
    1.178607e-10, 1.181905e-10, 1.194671e-10, 1.197485e-10, 1.200095e-10, 
    1.205259e-10, 1.211899e-10, 1.223585e-10, 1.233792e-10, 1.243142e-10, 
    1.242456e-10, 1.242697e-10, 1.24479e-10, 1.23961e-10, 1.245641e-10, 
    1.246654e-10, 1.244005e-10, 1.259412e-10, 1.255002e-10, 1.259515e-10, 
    1.256643e-10, 1.18536e-10, 1.188852e-10, 1.186965e-10, 1.190515e-10, 
    1.188013e-10, 1.199155e-10, 1.202505e-10, 1.218232e-10, 1.211768e-10, 
    1.222063e-10, 1.212812e-10, 1.214449e-10, 1.222398e-10, 1.213312e-10, 
    1.233227e-10, 1.219709e-10, 1.244871e-10, 1.231315e-10, 1.245722e-10, 
    1.243101e-10, 1.247443e-10, 1.251335e-10, 1.256241e-10, 1.265312e-10, 
    1.263209e-10, 1.270812e-10, 1.194067e-10, 1.198612e-10, 1.198212e-10, 
    1.202975e-10, 1.206504e-10, 1.214166e-10, 1.226499e-10, 1.221855e-10, 
    1.230387e-10, 1.232102e-10, 1.219144e-10, 1.227092e-10, 1.201658e-10, 
    1.205751e-10, 1.203314e-10, 1.194425e-10, 1.222924e-10, 1.208262e-10, 
    1.235396e-10, 1.227409e-10, 1.25078e-10, 1.239133e-10, 1.262052e-10, 
    1.271902e-10, 1.281205e-10, 1.292108e-10, 1.201096e-10, 1.198004e-10, 
    1.203543e-10, 1.211222e-10, 1.218368e-10, 1.227896e-10, 1.228873e-10, 
    1.230661e-10, 1.235301e-10, 1.239207e-10, 1.231226e-10, 1.240187e-10, 
    1.206699e-10, 1.2242e-10, 1.196836e-10, 1.205047e-10, 1.210769e-10, 
    1.208258e-10, 1.221325e-10, 1.224413e-10, 1.236997e-10, 1.230486e-10, 
    1.269467e-10, 1.252157e-10, 1.300439e-10, 1.286869e-10, 1.196925e-10, 
    1.201085e-10, 1.215613e-10, 1.208692e-10, 1.228533e-10, 1.233438e-10, 
    1.237432e-10, 1.242544e-10, 1.243097e-10, 1.246131e-10, 1.241161e-10, 
    1.245935e-10, 1.227916e-10, 1.235954e-10, 1.21395e-10, 1.21929e-10, 
    1.216832e-10, 1.214138e-10, 1.22246e-10, 1.231352e-10, 1.231543e-10, 
    1.2344e-10, 1.242463e-10, 1.228614e-10, 1.271706e-10, 1.245017e-10, 
    1.205629e-10, 1.213672e-10, 1.214825e-10, 1.211705e-10, 1.232946e-10, 
    1.225231e-10, 1.246057e-10, 1.240414e-10, 1.249666e-10, 1.245065e-10, 
    1.244388e-10, 1.238491e-10, 1.234825e-10, 1.225584e-10, 1.218087e-10, 
    1.212157e-10, 1.213535e-10, 1.220053e-10, 1.231897e-10, 1.243147e-10, 
    1.240678e-10, 1.248962e-10, 1.22709e-10, 1.236241e-10, 1.2327e-10, 
    1.241941e-10, 1.221732e-10, 1.238929e-10, 1.217352e-10, 1.219238e-10, 
    1.225078e-10, 1.236861e-10, 1.239477e-10, 1.242269e-10, 1.240546e-10, 
    1.232198e-10, 1.230833e-10, 1.224936e-10, 1.22331e-10, 1.218827e-10, 
    1.215121e-10, 1.218507e-10, 1.222066e-10, 1.232202e-10, 1.241366e-10, 
    1.251391e-10, 1.25385e-10, 1.265612e-10, 1.256032e-10, 1.271855e-10, 
    1.258394e-10, 1.281735e-10, 1.23993e-10, 1.258002e-10, 1.225345e-10, 
    1.228845e-10, 1.235187e-10, 1.249788e-10, 1.241898e-10, 1.251128e-10, 
    1.23078e-10, 1.220277e-10, 1.217568e-10, 1.212517e-10, 1.217684e-10, 
    1.217263e-10, 1.222215e-10, 1.220623e-10, 1.232539e-10, 1.226132e-10, 
    1.244371e-10, 1.251055e-10, 1.270014e-10, 1.281694e-10, 1.293633e-10, 
    1.298917e-10, 1.300528e-10, 1.301201e-10,
  1.205399e-10, 1.216865e-10, 1.214632e-10, 1.22391e-10, 1.218759e-10, 
    1.224841e-10, 1.207719e-10, 1.217321e-10, 1.211187e-10, 1.206429e-10, 
    1.242013e-10, 1.224325e-10, 1.260518e-10, 1.249141e-10, 1.277816e-10, 
    1.258744e-10, 1.281678e-10, 1.277264e-10, 1.290573e-10, 1.286753e-10, 
    1.303848e-10, 1.292338e-10, 1.312752e-10, 1.301095e-10, 1.302915e-10, 
    1.291959e-10, 1.227875e-10, 1.239804e-10, 1.22717e-10, 1.228867e-10, 
    1.228105e-10, 1.218865e-10, 1.214221e-10, 1.204525e-10, 1.206282e-10, 
    1.213406e-10, 1.229631e-10, 1.224112e-10, 1.238045e-10, 1.237729e-10, 
    1.253329e-10, 1.246283e-10, 1.272644e-10, 1.265125e-10, 1.286913e-10, 
    1.281416e-10, 1.286654e-10, 1.285065e-10, 1.286675e-10, 1.278619e-10, 
    1.282067e-10, 1.274989e-10, 1.247601e-10, 1.25562e-10, 1.231777e-10, 
    1.217546e-10, 1.208139e-10, 1.201485e-10, 1.202425e-10, 1.204217e-10, 
    1.213448e-10, 1.222157e-10, 1.228815e-10, 1.233278e-10, 1.237684e-10, 
    1.251064e-10, 1.258175e-10, 1.274167e-10, 1.271274e-10, 1.276177e-10, 
    1.28087e-10, 1.288768e-10, 1.287466e-10, 1.290951e-10, 1.276048e-10, 
    1.285943e-10, 1.269628e-10, 1.27408e-10, 1.238881e-10, 1.225599e-10, 
    1.219974e-10, 1.215061e-10, 1.203148e-10, 1.211369e-10, 1.208125e-10, 
    1.215849e-10, 1.22077e-10, 1.218335e-10, 1.233401e-10, 1.227533e-10, 
    1.258597e-10, 1.245171e-10, 1.280322e-10, 1.271868e-10, 1.282353e-10, 
    1.276998e-10, 1.28618e-10, 1.277914e-10, 1.29225e-10, 1.295381e-10, 
    1.293241e-10, 1.301472e-10, 1.277457e-10, 1.286654e-10, 1.218267e-10, 
    1.218664e-10, 1.220514e-10, 1.212391e-10, 1.211895e-10, 1.204477e-10, 
    1.211077e-10, 1.213893e-10, 1.221056e-10, 1.225302e-10, 1.229345e-10, 
    1.238258e-10, 1.248249e-10, 1.262284e-10, 1.272415e-10, 1.279228e-10, 
    1.275048e-10, 1.278738e-10, 1.274614e-10, 1.272683e-10, 1.294207e-10, 
    1.282099e-10, 1.300287e-10, 1.299277e-10, 1.291034e-10, 1.299391e-10, 
    1.218943e-10, 1.216659e-10, 1.208746e-10, 1.214937e-10, 1.20367e-10, 
    1.20997e-10, 1.2136e-10, 1.227655e-10, 1.230754e-10, 1.233631e-10, 
    1.239322e-10, 1.246644e-10, 1.259539e-10, 1.270811e-10, 1.281144e-10, 
    1.280385e-10, 1.280652e-10, 1.282965e-10, 1.277239e-10, 1.283907e-10, 
    1.285027e-10, 1.282098e-10, 1.299142e-10, 1.294262e-10, 1.299256e-10, 
    1.296077e-10, 1.217401e-10, 1.221246e-10, 1.219168e-10, 1.223077e-10, 
    1.220322e-10, 1.232595e-10, 1.236287e-10, 1.253631e-10, 1.246499e-10, 
    1.257859e-10, 1.247651e-10, 1.249457e-10, 1.25823e-10, 1.248202e-10, 
    1.270188e-10, 1.255261e-10, 1.283055e-10, 1.268076e-10, 1.283997e-10, 
    1.281099e-10, 1.285899e-10, 1.290205e-10, 1.295632e-10, 1.305675e-10, 
    1.303346e-10, 1.311767e-10, 1.226989e-10, 1.231996e-10, 1.231555e-10, 
    1.236805e-10, 1.240694e-10, 1.249145e-10, 1.262756e-10, 1.257629e-10, 
    1.267049e-10, 1.268944e-10, 1.254636e-10, 1.263411e-10, 1.235353e-10, 
    1.239865e-10, 1.237177e-10, 1.227383e-10, 1.258809e-10, 1.242633e-10, 
    1.272583e-10, 1.263761e-10, 1.28959e-10, 1.276713e-10, 1.302065e-10, 
    1.312976e-10, 1.323285e-10, 1.335381e-10, 1.234733e-10, 1.231326e-10, 
    1.23743e-10, 1.245898e-10, 1.253781e-10, 1.264298e-10, 1.265377e-10, 
    1.267352e-10, 1.272477e-10, 1.276794e-10, 1.267977e-10, 1.277877e-10, 
    1.240912e-10, 1.260218e-10, 1.230039e-10, 1.239089e-10, 1.245398e-10, 
    1.242629e-10, 1.257044e-10, 1.260453e-10, 1.274352e-10, 1.267158e-10, 
    1.310278e-10, 1.291115e-10, 1.344628e-10, 1.329568e-10, 1.230137e-10, 
    1.234721e-10, 1.250741e-10, 1.243107e-10, 1.265002e-10, 1.270419e-10, 
    1.274832e-10, 1.280483e-10, 1.281094e-10, 1.284449e-10, 1.278954e-10, 
    1.284231e-10, 1.26432e-10, 1.2732e-10, 1.248906e-10, 1.254798e-10, 
    1.252085e-10, 1.249114e-10, 1.258297e-10, 1.268115e-10, 1.268326e-10, 
    1.271483e-10, 1.280396e-10, 1.265091e-10, 1.312761e-10, 1.28322e-10, 
    1.23973e-10, 1.248601e-10, 1.249871e-10, 1.246429e-10, 1.269876e-10, 
    1.261356e-10, 1.284367e-10, 1.278128e-10, 1.288358e-10, 1.28327e-10, 
    1.282522e-10, 1.276003e-10, 1.271952e-10, 1.261746e-10, 1.253471e-10, 
    1.246928e-10, 1.248448e-10, 1.25564e-10, 1.268717e-10, 1.281149e-10, 
    1.278421e-10, 1.287579e-10, 1.263408e-10, 1.273516e-10, 1.269605e-10, 
    1.279816e-10, 1.257493e-10, 1.276489e-10, 1.252659e-10, 1.25474e-10, 
    1.261187e-10, 1.274203e-10, 1.277092e-10, 1.280179e-10, 1.278274e-10, 
    1.26905e-10, 1.267542e-10, 1.26103e-10, 1.259235e-10, 1.254287e-10, 
    1.250197e-10, 1.253933e-10, 1.257863e-10, 1.269054e-10, 1.279181e-10, 
    1.290266e-10, 1.292986e-10, 1.306008e-10, 1.295402e-10, 1.312926e-10, 
    1.29802e-10, 1.323876e-10, 1.277595e-10, 1.297583e-10, 1.261481e-10, 
    1.265347e-10, 1.272353e-10, 1.288494e-10, 1.279768e-10, 1.289976e-10, 
    1.267483e-10, 1.255888e-10, 1.252897e-10, 1.247325e-10, 1.253025e-10, 
    1.252561e-10, 1.258026e-10, 1.256268e-10, 1.269427e-10, 1.262351e-10, 
    1.282503e-10, 1.289895e-10, 1.310883e-10, 1.323829e-10, 1.337072e-10, 
    1.342938e-10, 1.344726e-10, 1.345473e-10,
  1.315636e-10, 1.327923e-10, 1.325529e-10, 1.335477e-10, 1.329953e-10, 
    1.336475e-10, 1.318122e-10, 1.328412e-10, 1.321838e-10, 1.316739e-10, 
    1.354906e-10, 1.335922e-10, 1.374788e-10, 1.36256e-10, 1.393397e-10, 
    1.372882e-10, 1.397556e-10, 1.392803e-10, 1.407135e-10, 1.403021e-10, 
    1.421447e-10, 1.409037e-10, 1.431054e-10, 1.418478e-10, 1.420441e-10, 
    1.408629e-10, 1.33973e-10, 1.352534e-10, 1.338973e-10, 1.340794e-10, 
    1.339977e-10, 1.330067e-10, 1.32509e-10, 1.314699e-10, 1.316582e-10, 
    1.324215e-10, 1.341614e-10, 1.335693e-10, 1.350643e-10, 1.350304e-10, 
    1.367059e-10, 1.35949e-10, 1.387831e-10, 1.379741e-10, 1.403192e-10, 
    1.397273e-10, 1.402914e-10, 1.401202e-10, 1.402936e-10, 1.394261e-10, 
    1.397974e-10, 1.390354e-10, 1.360906e-10, 1.369523e-10, 1.343916e-10, 
    1.328655e-10, 1.318572e-10, 1.311444e-10, 1.312451e-10, 1.31437e-10, 
    1.32426e-10, 1.333597e-10, 1.340738e-10, 1.345527e-10, 1.350256e-10, 
    1.364627e-10, 1.372269e-10, 1.38947e-10, 1.386356e-10, 1.391633e-10, 
    1.396685e-10, 1.405191e-10, 1.403789e-10, 1.407543e-10, 1.391494e-10, 
    1.402149e-10, 1.384584e-10, 1.389376e-10, 1.351544e-10, 1.337289e-10, 
    1.331257e-10, 1.325989e-10, 1.313225e-10, 1.322032e-10, 1.318556e-10, 
    1.326834e-10, 1.33211e-10, 1.329499e-10, 1.345658e-10, 1.339363e-10, 
    1.372723e-10, 1.358295e-10, 1.396095e-10, 1.386995e-10, 1.398281e-10, 
    1.392515e-10, 1.402404e-10, 1.393503e-10, 1.408942e-10, 1.412318e-10, 
    1.410011e-10, 1.418884e-10, 1.39301e-10, 1.402914e-10, 1.329426e-10, 
    1.329851e-10, 1.331835e-10, 1.323128e-10, 1.322596e-10, 1.314648e-10, 
    1.321719e-10, 1.324737e-10, 1.332416e-10, 1.33697e-10, 1.341307e-10, 
    1.350872e-10, 1.361602e-10, 1.376687e-10, 1.387584e-10, 1.394916e-10, 
    1.390417e-10, 1.394389e-10, 1.38995e-10, 1.387872e-10, 1.411052e-10, 
    1.398009e-10, 1.417606e-10, 1.416517e-10, 1.407633e-10, 1.41664e-10, 
    1.33015e-10, 1.327702e-10, 1.319222e-10, 1.325856e-10, 1.313784e-10, 
    1.320533e-10, 1.324423e-10, 1.339494e-10, 1.342818e-10, 1.345905e-10, 
    1.352014e-10, 1.359877e-10, 1.373734e-10, 1.385858e-10, 1.396979e-10, 
    1.396162e-10, 1.39645e-10, 1.398941e-10, 1.392775e-10, 1.399955e-10, 
    1.401162e-10, 1.398007e-10, 1.416372e-10, 1.411111e-10, 1.416494e-10, 
    1.413067e-10, 1.328497e-10, 1.33262e-10, 1.330391e-10, 1.334584e-10, 
    1.33163e-10, 1.344795e-10, 1.348757e-10, 1.367385e-10, 1.359722e-10, 
    1.371929e-10, 1.360959e-10, 1.362899e-10, 1.372329e-10, 1.36155e-10, 
    1.385188e-10, 1.369137e-10, 1.399038e-10, 1.382917e-10, 1.400052e-10, 
    1.396931e-10, 1.4021e-10, 1.406739e-10, 1.412588e-10, 1.423418e-10, 
    1.420906e-10, 1.42999e-10, 1.338779e-10, 1.344151e-10, 1.343678e-10, 
    1.349312e-10, 1.353488e-10, 1.362563e-10, 1.377193e-10, 1.371681e-10, 
    1.38181e-10, 1.383849e-10, 1.368464e-10, 1.377899e-10, 1.347754e-10, 
    1.352598e-10, 1.349712e-10, 1.339203e-10, 1.372951e-10, 1.355571e-10, 
    1.387764e-10, 1.378274e-10, 1.406077e-10, 1.39221e-10, 1.419524e-10, 
    1.431296e-10, 1.442426e-10, 1.455498e-10, 1.347088e-10, 1.343432e-10, 
    1.349983e-10, 1.359077e-10, 1.367545e-10, 1.378852e-10, 1.380012e-10, 
    1.382137e-10, 1.38765e-10, 1.392296e-10, 1.382809e-10, 1.393462e-10, 
    1.353724e-10, 1.374465e-10, 1.342052e-10, 1.351765e-10, 1.35854e-10, 
    1.355565e-10, 1.371052e-10, 1.374717e-10, 1.389669e-10, 1.381928e-10, 
    1.428385e-10, 1.407721e-10, 1.465497e-10, 1.449214e-10, 1.342156e-10, 
    1.347076e-10, 1.36428e-10, 1.356078e-10, 1.379608e-10, 1.385436e-10, 
    1.390184e-10, 1.396268e-10, 1.396926e-10, 1.400539e-10, 1.394621e-10, 
    1.400304e-10, 1.378876e-10, 1.388428e-10, 1.362306e-10, 1.368638e-10, 
    1.365723e-10, 1.36253e-10, 1.372399e-10, 1.382958e-10, 1.383184e-10, 
    1.386581e-10, 1.396178e-10, 1.379704e-10, 1.431066e-10, 1.399218e-10, 
    1.352452e-10, 1.36198e-10, 1.363344e-10, 1.359646e-10, 1.384851e-10, 
    1.375688e-10, 1.40045e-10, 1.393732e-10, 1.404749e-10, 1.399269e-10, 
    1.398463e-10, 1.391445e-10, 1.387085e-10, 1.376107e-10, 1.367212e-10, 
    1.360182e-10, 1.361815e-10, 1.369544e-10, 1.383606e-10, 1.396985e-10, 
    1.394048e-10, 1.40391e-10, 1.377894e-10, 1.388769e-10, 1.38456e-10, 
    1.39555e-10, 1.371535e-10, 1.391971e-10, 1.36634e-10, 1.368576e-10, 
    1.375506e-10, 1.389509e-10, 1.392617e-10, 1.395941e-10, 1.39389e-10, 
    1.383964e-10, 1.382341e-10, 1.375337e-10, 1.373407e-10, 1.368089e-10, 
    1.363694e-10, 1.367709e-10, 1.371933e-10, 1.383968e-10, 1.394866e-10, 
    1.406805e-10, 1.409736e-10, 1.423779e-10, 1.412342e-10, 1.431245e-10, 
    1.415165e-10, 1.443067e-10, 1.39316e-10, 1.414693e-10, 1.375822e-10, 
    1.379979e-10, 1.387518e-10, 1.404897e-10, 1.395498e-10, 1.406493e-10, 
    1.382278e-10, 1.369811e-10, 1.366596e-10, 1.360609e-10, 1.366733e-10, 
    1.366234e-10, 1.372107e-10, 1.370218e-10, 1.384368e-10, 1.376757e-10, 
    1.398443e-10, 1.406406e-10, 1.429036e-10, 1.443014e-10, 1.457324e-10, 
    1.463669e-10, 1.465603e-10, 1.466412e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24574.34, 24594.61, 24590.64, 24607.23, 24597.99, 24608.9, 24578.41, 
    24595.43, 24584.53, 24576.14, 24640.15, 24607.97, 24674.59, 24653.3, 
    24707.2, 24671.24, 24714.59, 24706.14, 24731.79, 24724.37, 24757.96, 
    24735.23, 24775.87, 24752.48, 24756.1, 24734.49, 24614.38, 24636.1, 
    24613.1, 24616.17, 24614.79, 24598.18, 24589.91, 24572.8, 24575.88, 
    24588.46, 24617.56, 24607.59, 24632.87, 24632.3, 24661.09, 24648, 
    24697.38, 24683.24, 24724.68, 24714.08, 24724.18, 24721.11, 24724.22, 
    24708.73, 24715.33, 24701.82, 24650.44, 24665.38, 24621.46, 24595.83, 
    24579.15, 24567.48, 24569.13, 24572.26, 24588.54, 24604.08, 24616.08, 
    24624.19, 24632.21, 24656.88, 24670.17, 24700.26, 24694.79, 24704.08, 
    24713.04, 24728.28, 24725.75, 24732.53, 24703.83, 24722.8, 24691.68, 
    24700.09, 24634.41, 24610.27, 24600.17, 24591.4, 24570.39, 24584.85, 
    24579.13, 24592.8, 24601.59, 24597.23, 24624.41, 24613.76, 24670.97, 
    24645.95, 24711.99, 24695.91, 24715.88, 24705.64, 24723.26, 24707.38, 
    24735.06, 24741.2, 24737, 24753.23, 24706.51, 24724.18, 24597.11, 
    24597.82, 24601.13, 24586.66, 24585.79, 24572.72, 24584.34, 24589.33, 
    24602.1, 24609.73, 24617.04, 24633.26, 24651.64, 24677.92, 24696.94, 
    24709.89, 24701.93, 24708.96, 24701.11, 24697.45, 24738.89, 24715.4, 
    24750.88, 24748.88, 24732.69, 24749.11, 24598.32, 24594.24, 24580.22, 
    24591.18, 24571.3, 24582.38, 24588.81, 24613.98, 24619.59, 24624.83, 
    24635.21, 24648.67, 24672.74, 24693.91, 24713.56, 24712.11, 24712.62, 
    24717.06, 24706.1, 24718.87, 24721.03, 24715.39, 24748.61, 24739, 
    24748.84, 24742.56, 24595.57, 24602.44, 24598.72, 24605.73, 24600.79, 
    24622.95, 24629.67, 24661.66, 24648.4, 24669.58, 24650.53, 24653.88, 
    24670.28, 24651.55, 24692.74, 24664.71, 24717.23, 24688.78, 24719.04, 
    24713.47, 24722.71, 24731.07, 24741.69, 24761.61, 24756.96, 24773.87, 
    24612.77, 24621.85, 24621.05, 24630.61, 24637.72, 24653.3, 24678.81, 
    24669.14, 24686.84, 24690.4, 24663.54, 24680.05, 24627.97, 24636.2, 
    24631.29, 24613.49, 24671.37, 24641.28, 24697.26, 24680.7, 24729.88, 
    24705.1, 24754.41, 24776.33, 24797.42, 24822.48, 24626.84, 24620.63, 
    24631.75, 24647.29, 24661.94, 24681.7, 24683.71, 24687.41, 24697.06, 
    24705.25, 24688.59, 24707.31, 24638.12, 24674.02, 24618.3, 24634.78, 
    24646.37, 24641.27, 24668.04, 24674.46, 24700.61, 24687.05, 24770.87, 
    24732.85, 24841.78, 24810.46, 24618.47, 24626.82, 24656.27, 24642.15, 
    24683.01, 24693.18, 24701.52, 24712.29, 24713.46, 24719.92, 24709.37, 
    24719.5, 24681.74, 24698.43, 24652.86, 24663.84, 24658.77, 24653.24, 
    24670.4, 24688.85, 24689.24, 24695.18, 24712.14, 24683.18, 24775.9, 
    24717.56, 24635.95, 24652.29, 24654.65, 24648.27, 24692.15, 24676.16, 
    24719.76, 24707.79, 24727.48, 24717.64, 24716.21, 24703.74, 24696.07, 
    24676.9, 24661.36, 24649.19, 24652.01, 24665.42, 24689.98, 24713.57, 
    24708.35, 24725.97, 24680.04, 24699.03, 24691.64, 24711.02, 24668.89, 
    24704.68, 24659.84, 24663.73, 24675.84, 24700.33, 24705.82, 24711.71, 
    24708.07, 24690.6, 24687.77, 24675.55, 24672.16, 24662.88, 24655.26, 
    24662.22, 24669.58, 24690.61, 24709.8, 24731.19, 24736.5, 24762.29, 
    24741.24, 24776.23, 24746.41, 24798.65, 24706.78, 24745.54, 24676.4, 
    24683.66, 24696.83, 24727.75, 24710.93, 24730.63, 24687.66, 24665.88, 
    24660.29, 24649.93, 24660.52, 24659.66, 24669.89, 24666.59, 24691.31, 
    24678.04, 24716.17, 24730.47, 24772.09, 24798.54, 24825.99, 24838.23, 
    24841.98, 24843.55 ;

 GC_ICE1 =
  17683.55, 17716.04, 17709.67, 17736.23, 17721.45, 17738.92, 17690.08, 
    17717.34, 17699.88, 17686.45, 17788.93, 17737.43, 17844.02, 17809.97, 
    17896.08, 17838.68, 17907.87, 17894.4, 17935.31, 17923.47, 17977.06, 
    17940.8, 18005.62, 17968.32, 17974.09, 17939.62, 17747.68, 17782.45, 
    17745.64, 17750.56, 17748.35, 17721.75, 17708.5, 17681.09, 17686.04, 
    17706.18, 17752.78, 17736.81, 17777.29, 17776.37, 17822.44, 17801.5, 
    17880.41, 17857.85, 17923.96, 17907.06, 17923.17, 17918.26, 17923.23, 
    17898.52, 17909.06, 17887.49, 17805.4, 17829.3, 17759.02, 17717.99, 
    17691.27, 17672.57, 17675.21, 17680.23, 17706.3, 17731.19, 17750.41, 
    17763.39, 17776.24, 17815.7, 17836.96, 17885.01, 17876.28, 17891.1, 
    17905.39, 17929.71, 17925.67, 17936.48, 17890.7, 17920.97, 17871.32, 
    17884.74, 17779.76, 17741.1, 17724.93, 17710.89, 17677.23, 17700.4, 
    17691.23, 17713.13, 17727.21, 17720.23, 17763.75, 17746.69, 17838.23, 
    17798.22, 17903.72, 17878.06, 17909.93, 17893.58, 17921.71, 17896.37, 
    17940.53, 17950.32, 17943.62, 17969.51, 17894.98, 17923.17, 17720.04, 
    17721.18, 17726.47, 17703.3, 17701.89, 17680.96, 17699.57, 17707.56, 
    17728.02, 17740.24, 17751.95, 17777.92, 17807.32, 17849.35, 17879.71, 
    17900.38, 17887.67, 17898.88, 17886.36, 17880.52, 17946.64, 17909.16, 
    17965.76, 17962.57, 17936.74, 17962.93, 17721.97, 17715.44, 17692.98, 
    17710.53, 17678.7, 17696.44, 17706.73, 17747.05, 17756.04, 17764.42, 
    17781.03, 17802.56, 17841.06, 17874.88, 17906.23, 17903.91, 17904.72, 
    17911.81, 17894.32, 17914.7, 17918.15, 17909.15, 17962.14, 17946.81, 
    17962.5, 17952.5, 17717.56, 17728.57, 17722.62, 17733.83, 17725.92, 
    17761.41, 17772.17, 17823.35, 17802.14, 17836.01, 17805.55, 17810.91, 
    17837.13, 17807.18, 17873.01, 17828.23, 17912.09, 17866.68, 17914.98, 
    17906.09, 17920.83, 17934.16, 17951.1, 17982.88, 17975.46, 18002.43, 
    17745.12, 17759.66, 17758.37, 17773.68, 17785.05, 17809.98, 17850.78, 
    17835.32, 17863.6, 17869.27, 17826.35, 17852.76, 17769.45, 17782.62, 
    17774.77, 17746.26, 17838.87, 17790.74, 17880.22, 17853.79, 17932.26, 
    17892.73, 17971.39, 18006.34, 18039.97, 18079.88, 17767.65, 17757.7, 
    17775.5, 17800.37, 17823.79, 17855.39, 17858.6, 17864.51, 17879.9, 
    17892.96, 17866.38, 17896.26, 17785.7, 17843.11, 17753.96, 17780.35, 
    17798.89, 17790.73, 17833.56, 17843.82, 17885.57, 17863.92, 17997.64, 
    17937, 18110.54, 18060.75, 17754.24, 17767.61, 17814.73, 17792.13, 
    17857.49, 17873.71, 17887.02, 17904.21, 17906.08, 17916.37, 17899.54, 
    17915.7, 17855.46, 17882.08, 17809.27, 17826.83, 17818.73, 17809.88, 
    17837.32, 17866.79, 17867.42, 17876.9, 17903.96, 17857.75, 18005.66, 
    17912.61, 17782.22, 17808.37, 17812.13, 17801.93, 17872.07, 17846.54, 
    17916.12, 17897.02, 17928.43, 17912.74, 17910.45, 17890.56, 17878.32, 
    17847.72, 17822.87, 17803.4, 17807.91, 17829.36, 17868.6, 17906.25, 
    17897.92, 17926.02, 17852.74, 17883.04, 17871.26, 17902.17, 17834.91, 
    17892.06, 17820.44, 17826.66, 17846.03, 17885.12, 17893.87, 17903.28, 
    17897.47, 17869.6, 17865.08, 17845.56, 17840.15, 17825.3, 17813.1, 
    17824.25, 17836.02, 17869.61, 17900.23, 17934.36, 17942.82, 17983.95, 
    17950.39, 18006.2, 17958.63, 18041.93, 17895.41, 17957.24, 17846.92, 
    17858.51, 17879.53, 17928.86, 17902.03, 17933.46, 17864.9, 17830.1, 
    17821.15, 17804.58, 17821.53, 17820.14, 17836.51, 17831.23, 17870.72, 
    17849.55, 17910.39, 17933.21, 17999.58, 18041.77, 18085.45, 18104.9, 
    18110.87, 18113.37 ;

 GC_LIQ1 =
  5232.713, 5234.742, 5234.344, 5236.006, 5235.081, 5236.174, 5233.121, 
    5234.824, 5233.733, 5232.894, 5239.315, 5236.081, 5242.794, 5240.642, 
    5246.144, 5242.456, 5246.906, 5246.036, 5248.679, 5247.914, 5251.38, 
    5249.034, 5253.229, 5250.814, 5251.188, 5248.958, 5236.723, 5238.906, 
    5236.595, 5236.903, 5236.764, 5235.1, 5234.272, 5232.56, 5232.869, 
    5234.127, 5237.042, 5236.042, 5238.581, 5238.522, 5241.43, 5240.108, 
    5245.132, 5243.676, 5247.946, 5246.854, 5247.894, 5247.578, 5247.898, 
    5246.302, 5246.982, 5245.59, 5240.354, 5241.863, 5237.432, 5234.864, 
    5233.195, 5232.028, 5232.192, 5232.506, 5234.134, 5235.69, 5236.893, 
    5237.706, 5238.514, 5241.004, 5242.348, 5245.429, 5244.865, 5245.822, 
    5246.746, 5248.317, 5248.057, 5248.755, 5245.797, 5247.752, 5244.546, 
    5245.412, 5238.736, 5236.311, 5235.298, 5234.421, 5232.319, 5233.766, 
    5233.193, 5234.561, 5235.441, 5235.005, 5237.729, 5236.66, 5242.428, 
    5239.9, 5246.638, 5244.981, 5247.039, 5245.983, 5247.8, 5246.163, 
    5249.017, 5249.65, 5249.217, 5250.892, 5246.073, 5247.895, 5234.993, 
    5235.063, 5235.395, 5233.947, 5233.859, 5232.552, 5233.714, 5234.213, 
    5235.492, 5236.257, 5236.989, 5238.62, 5240.475, 5243.131, 5245.087, 
    5246.421, 5245.601, 5246.325, 5245.516, 5245.139, 5249.412, 5246.989, 
    5250.649, 5250.442, 5248.772, 5250.466, 5235.113, 5234.706, 5233.302, 
    5234.398, 5232.41, 5233.518, 5234.161, 5236.683, 5237.246, 5237.771, 
    5238.816, 5240.175, 5242.607, 5244.775, 5246.8, 5246.65, 5246.703, 
    5247.16, 5246.03, 5247.347, 5247.57, 5246.988, 5250.415, 5249.423, 
    5250.438, 5249.791, 5234.838, 5235.526, 5235.154, 5235.855, 5235.36, 
    5237.582, 5238.258, 5241.487, 5240.148, 5242.288, 5240.363, 5240.701, 
    5242.358, 5240.466, 5244.655, 5241.795, 5247.178, 5244.246, 5247.365, 
    5246.791, 5247.744, 5248.605, 5249.701, 5251.757, 5251.277, 5253.023, 
    5236.562, 5237.472, 5237.392, 5238.353, 5239.07, 5240.643, 5243.222, 
    5242.244, 5244.047, 5244.414, 5241.676, 5243.348, 5238.086, 5238.917, 
    5238.421, 5236.633, 5242.468, 5239.429, 5245.12, 5243.415, 5248.482, 
    5245.928, 5251.014, 5253.277, 5255.458, 5258.077, 5237.973, 5237.35, 
    5238.467, 5240.036, 5241.515, 5243.518, 5243.725, 5244.105, 5245.099, 
    5245.943, 5244.227, 5246.156, 5239.111, 5242.737, 5237.116, 5238.773, 
    5239.943, 5239.428, 5242.132, 5242.781, 5245.465, 5244.068, 5252.713, 
    5248.789, 5260.122, 5256.811, 5237.133, 5237.97, 5240.942, 5239.517, 
    5243.653, 5244.699, 5245.559, 5246.669, 5246.79, 5247.455, 5246.368, 
    5247.412, 5243.522, 5245.24, 5240.598, 5241.707, 5241.195, 5240.637, 
    5242.371, 5244.253, 5244.294, 5244.906, 5246.653, 5243.67, 5253.232, 
    5247.212, 5238.892, 5240.542, 5240.779, 5240.135, 5244.594, 5242.954, 
    5247.438, 5246.205, 5248.235, 5247.221, 5247.072, 5245.788, 5244.997, 
    5243.028, 5241.457, 5240.228, 5240.512, 5241.867, 5244.37, 5246.801, 
    5246.263, 5248.079, 5243.347, 5245.302, 5244.542, 5246.538, 5242.218, 
    5245.884, 5241.303, 5241.696, 5242.921, 5245.437, 5246.001, 5246.609, 
    5246.234, 5244.434, 5244.143, 5242.892, 5242.549, 5241.61, 5240.84, 
    5241.543, 5242.288, 5244.435, 5246.413, 5248.618, 5249.165, 5251.827, 
    5249.655, 5253.268, 5250.188, 5255.586, 5246.101, 5250.098, 5242.978, 
    5243.719, 5245.076, 5248.263, 5246.528, 5248.56, 5244.131, 5241.914, 
    5241.348, 5240.302, 5241.372, 5241.285, 5242.319, 5241.985, 5244.507, 
    5243.144, 5247.069, 5248.543, 5252.839, 5255.575, 5258.447, 5259.745, 
    5260.144, 5260.311 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.728482e-09, 8.766966e-09, 8.759486e-09, 8.790525e-09, 8.773307e-09, 
    8.793632e-09, 8.736285e-09, 8.768493e-09, 8.747932e-09, 8.731948e-09, 
    8.850763e-09, 8.79191e-09, 8.911909e-09, 8.87437e-09, 8.968676e-09, 
    8.906067e-09, 8.981302e-09, 8.966873e-09, 9.010307e-09, 8.997864e-09, 
    9.053418e-09, 9.016051e-09, 9.082221e-09, 9.044496e-09, 9.050396e-09, 
    9.014817e-09, 8.803755e-09, 8.843435e-09, 8.801404e-09, 8.807063e-09, 
    8.804523e-09, 8.773662e-09, 8.758109e-09, 8.725542e-09, 8.731455e-09, 
    8.755375e-09, 8.809606e-09, 8.791198e-09, 8.837596e-09, 8.836548e-09, 
    8.888205e-09, 8.864914e-09, 8.951743e-09, 8.927064e-09, 8.998383e-09, 
    8.980447e-09, 8.99754e-09, 8.992357e-09, 8.997608e-09, 8.971302e-09, 
    8.982572e-09, 8.959426e-09, 8.869276e-09, 8.895769e-09, 8.816755e-09, 
    8.769247e-09, 8.737697e-09, 8.715308e-09, 8.718474e-09, 8.724507e-09, 
    8.755515e-09, 8.784671e-09, 8.80689e-09, 8.821753e-09, 8.836398e-09, 
    8.880725e-09, 8.90419e-09, 8.956733e-09, 8.947252e-09, 8.963315e-09, 
    8.978662e-09, 9.004427e-09, 9.000187e-09, 9.011539e-09, 8.962892e-09, 
    8.995221e-09, 8.941852e-09, 8.956448e-09, 8.840373e-09, 8.796165e-09, 
    8.777369e-09, 8.760923e-09, 8.720908e-09, 8.748541e-09, 8.737647e-09, 
    8.763565e-09, 8.780034e-09, 8.771889e-09, 8.822159e-09, 8.802615e-09, 
    8.905581e-09, 8.861229e-09, 8.976872e-09, 8.949198e-09, 8.983505e-09, 
    8.965999e-09, 8.995995e-09, 8.969e-09, 9.015764e-09, 9.025946e-09, 
    9.018988e-09, 9.045721e-09, 8.967502e-09, 8.99754e-09, 8.77166e-09, 
    8.772989e-09, 8.779177e-09, 8.751972e-09, 8.750308e-09, 8.72538e-09, 
    8.747562e-09, 8.757008e-09, 8.780988e-09, 8.795173e-09, 8.808657e-09, 
    8.838304e-09, 8.871416e-09, 8.917722e-09, 8.950992e-09, 8.973294e-09, 
    8.959619e-09, 8.971692e-09, 8.958196e-09, 8.95187e-09, 9.022131e-09, 
    8.982678e-09, 9.041876e-09, 9.0386e-09, 9.011808e-09, 9.03897e-09, 
    8.773921e-09, 8.766277e-09, 8.739736e-09, 8.760507e-09, 8.722665e-09, 
    8.743846e-09, 8.756025e-09, 8.803021e-09, 8.813349e-09, 8.822924e-09, 
    8.841836e-09, 8.866106e-09, 8.908684e-09, 8.945732e-09, 8.979556e-09, 
    8.977077e-09, 8.97795e-09, 8.985505e-09, 8.966789e-09, 8.988578e-09, 
    8.992234e-09, 8.982673e-09, 9.038161e-09, 9.022309e-09, 9.038531e-09, 
    9.028209e-09, 8.768763e-09, 8.781624e-09, 8.774674e-09, 8.787744e-09, 
    8.778536e-09, 8.819479e-09, 8.831756e-09, 8.889203e-09, 8.865628e-09, 
    8.90315e-09, 8.86944e-09, 8.875412e-09, 8.904371e-09, 8.871262e-09, 
    8.943688e-09, 8.894583e-09, 8.985799e-09, 8.936757e-09, 8.988872e-09, 
    8.979409e-09, 8.995078e-09, 9.009109e-09, 9.026764e-09, 9.059338e-09, 
    9.051796e-09, 9.079039e-09, 8.800801e-09, 8.817485e-09, 8.816016e-09, 
    8.833477e-09, 8.84639e-09, 8.87438e-09, 8.919273e-09, 8.902392e-09, 
    8.933386e-09, 8.939607e-09, 8.892521e-09, 8.92143e-09, 8.828651e-09, 
    8.843639e-09, 8.834716e-09, 8.802116e-09, 8.90628e-09, 8.852821e-09, 
    8.951542e-09, 8.922579e-09, 9.007108e-09, 8.965069e-09, 9.047643e-09, 
    9.082942e-09, 9.116171e-09, 9.154999e-09, 8.826591e-09, 8.815254e-09, 
    8.835554e-09, 8.863637e-09, 8.889699e-09, 8.924346e-09, 8.927891e-09, 
    8.934381e-09, 8.951195e-09, 8.965332e-09, 8.936433e-09, 8.968876e-09, 
    8.847112e-09, 8.910921e-09, 8.810968e-09, 8.841063e-09, 8.861982e-09, 
    8.852806e-09, 8.900463e-09, 8.911694e-09, 8.957338e-09, 8.933744e-09, 
    9.074228e-09, 9.012071e-09, 9.184567e-09, 9.136357e-09, 8.811294e-09, 
    8.826553e-09, 8.879659e-09, 8.854391e-09, 8.926659e-09, 8.944448e-09, 
    8.958911e-09, 8.977397e-09, 8.979393e-09, 8.990346e-09, 8.972398e-09, 
    8.989638e-09, 8.924419e-09, 8.953564e-09, 8.87359e-09, 8.893053e-09, 
    8.8841e-09, 8.874278e-09, 8.904593e-09, 8.936888e-09, 8.93758e-09, 
    8.947935e-09, 8.977112e-09, 8.926953e-09, 9.082248e-09, 8.986334e-09, 
    8.843192e-09, 8.872581e-09, 8.876782e-09, 8.865396e-09, 8.942664e-09, 
    8.914666e-09, 8.99008e-09, 8.969698e-09, 9.003094e-09, 8.986499e-09, 
    8.984057e-09, 8.962743e-09, 8.949474e-09, 8.91595e-09, 8.888675e-09, 
    8.867048e-09, 8.872076e-09, 8.895833e-09, 8.938863e-09, 8.979574e-09, 
    8.970655e-09, 9.000556e-09, 8.921419e-09, 8.954601e-09, 8.941775e-09, 
    8.975218e-09, 8.901943e-09, 8.964334e-09, 8.885995e-09, 8.892864e-09, 
    8.914111e-09, 8.956849e-09, 8.966309e-09, 8.976405e-09, 8.970176e-09, 
    8.939956e-09, 8.935006e-09, 8.913595e-09, 8.907683e-09, 8.891369e-09, 
    8.877862e-09, 8.890201e-09, 8.903161e-09, 8.93997e-09, 8.973141e-09, 
    9.009308e-09, 9.01816e-09, 9.060416e-09, 9.026015e-09, 9.082782e-09, 
    9.034516e-09, 9.118071e-09, 8.967953e-09, 9.0331e-09, 8.915078e-09, 
    8.927793e-09, 8.950789e-09, 9.003536e-09, 8.975061e-09, 9.008363e-09, 
    8.934812e-09, 8.896652e-09, 8.886782e-09, 8.868362e-09, 8.887203e-09, 
    8.885671e-09, 8.903699e-09, 8.897906e-09, 8.941192e-09, 8.91794e-09, 
    8.983995e-09, 9.008101e-09, 9.076182e-09, 9.11792e-09, 9.160412e-09, 
    9.17917e-09, 9.18488e-09, 9.187267e-09 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.257191, 6.286504, 6.280798, 6.30449, 6.291339, 6.306864, 6.263125, 
    6.287671, 6.271994, 6.259824, 6.350626, 6.305548, 6.39764, 6.368743, 
    6.441475, 6.39314, 6.451246, 6.440074, 6.473725, 6.464074, 6.507236, 
    6.478182, 6.529669, 6.500288, 6.504881, 6.477226, 6.3146, 6.345005, 
    6.312803, 6.317132, 6.315188, 6.291612, 6.279754, 6.254951, 6.259449, 
    6.277667, 6.319079, 6.305001, 6.340511, 6.339708, 6.379382, 6.361476, 
    6.428376, 6.409319, 6.464477, 6.45058, 6.463824, 6.459806, 6.463876, 
    6.443502, 6.452227, 6.434314, 6.364828, 6.385204, 6.324549, 6.28825, 
    6.264201, 6.247172, 6.249578, 6.254167, 6.277773, 6.300014, 6.316997, 
    6.328372, 6.339592, 6.373637, 6.391693, 6.432236, 6.424905, 6.437325, 
    6.449198, 6.469166, 6.465876, 6.474683, 6.436994, 6.462029, 6.420732, 
    6.432012, 6.342657, 6.308796, 6.294447, 6.281895, 6.251429, 6.272459, 
    6.264163, 6.283907, 6.296474, 6.290256, 6.328684, 6.313728, 6.392764, 
    6.358648, 6.447812, 6.426409, 6.452948, 6.439397, 6.462627, 6.441718, 
    6.477962, 6.48587, 6.480465, 6.501238, 6.44056, 6.463825, 6.290082, 
    6.291096, 6.295819, 6.275074, 6.273805, 6.254828, 6.271711, 6.27891, 
    6.297201, 6.308038, 6.318349, 6.341056, 6.366475, 6.402118, 6.427795, 
    6.445041, 6.434462, 6.443802, 6.433362, 6.428472, 6.482907, 6.452309, 
    6.498248, 6.495701, 6.474893, 6.495988, 6.291808, 6.285975, 6.265753, 
    6.281575, 6.252764, 6.268883, 6.278163, 6.314043, 6.321939, 6.329271, 
    6.343763, 6.362391, 6.395151, 6.423733, 6.449889, 6.44797, 6.448645, 
    6.454497, 6.440009, 6.456878, 6.459713, 6.452304, 6.49536, 6.483042, 
    6.495646, 6.487624, 6.28787, 6.297688, 6.292382, 6.302363, 6.295331, 
    6.326637, 6.336041, 6.380155, 6.362025, 6.390889, 6.364953, 6.369545, 
    6.391837, 6.366352, 6.422157, 6.384296, 6.454725, 6.416809, 6.457106, 
    6.449775, 6.461914, 6.472797, 6.486503, 6.511838, 6.505966, 6.527185, 
    6.31234, 6.325107, 6.32398, 6.337355, 6.347257, 6.368749, 6.403312, 
    6.390301, 6.414196, 6.419001, 6.382701, 6.404976, 6.333659, 6.345151, 
    6.338305, 6.313348, 6.393301, 6.352195, 6.42822, 6.40586, 6.471245, 
    6.438682, 6.502735, 6.530236, 6.556168, 6.586561, 6.332079, 6.323397, 
    6.338945, 6.360499, 6.380531, 6.407223, 6.409956, 6.414966, 6.427951, 
    6.438881, 6.416553, 6.441623, 6.347823, 6.396875, 6.320118, 6.343176, 
    6.359227, 6.35218, 6.388814, 6.397468, 6.432703, 6.414473, 6.523444, 
    6.475101, 6.609748, 6.571962, 6.320366, 6.332048, 6.37281, 6.353396, 
    6.409006, 6.42274, 6.433914, 6.44822, 6.449764, 6.458249, 6.444348, 
    6.457699, 6.40728, 6.429782, 6.368141, 6.383112, 6.376222, 6.36867, 
    6.391995, 6.416905, 6.417434, 6.425435, 6.448018, 6.409232, 6.529706, 
    6.455156, 6.344802, 6.367373, 6.370595, 6.361845, 6.421362, 6.399759, 
    6.458042, 6.442259, 6.46813, 6.455267, 6.453376, 6.436879, 6.426622, 
    6.40075, 6.379744, 6.363113, 6.366978, 6.385253, 6.418429, 6.449905, 
    6.443003, 6.466161, 6.404964, 6.430586, 6.420677, 6.446532, 6.389956, 
    6.438127, 6.377679, 6.382965, 6.399331, 6.432329, 6.439637, 6.447452, 
    6.442628, 6.419272, 6.415449, 6.398932, 6.394378, 6.381814, 6.371424, 
    6.380917, 6.390896, 6.419281, 6.444926, 6.472953, 6.479821, 6.512687, 
    6.48593, 6.530124, 6.492548, 6.557668, 6.440919, 6.491437, 6.400075, 
    6.40988, 6.427642, 6.46848, 6.44641, 6.472223, 6.415299, 6.385886, 
    6.378285, 6.364124, 6.378609, 6.377429, 6.391307, 6.386845, 6.420224, 
    6.402282, 6.453329, 6.472018, 6.524961, 6.557541, 6.590796, 6.605509, 
    6.609991, 6.611865,
  3.971761, 3.991221, 3.987432, 4.003165, 3.994431, 4.004741, 3.975699, 
    3.991996, 3.981587, 3.973508, 4.033811, 4.003867, 4.065043, 4.045842, 
    4.094177, 4.062054, 4.100673, 4.093244, 4.115616, 4.109199, 4.137903, 
    4.11858, 4.152823, 4.133281, 4.136336, 4.117944, 4.009878, 4.030077, 
    4.008684, 4.011559, 4.010268, 3.994613, 3.986741, 3.970273, 3.973259, 
    3.985354, 4.012853, 4.003502, 4.027086, 4.026553, 4.05291, 4.041013, 
    4.085469, 4.072803, 4.109467, 4.100228, 4.109033, 4.106361, 4.109068, 
    4.095523, 4.101323, 4.089416, 4.04324, 4.056779, 4.016485, 3.992383, 
    3.976414, 3.96511, 3.966707, 3.969753, 3.985425, 4.000191, 4.011468, 
    4.019024, 4.026476, 4.049097, 4.061091, 4.088035, 4.083161, 4.091417, 
    4.099309, 4.112585, 4.110397, 4.116253, 4.091197, 4.107841, 4.080387, 
    4.087885, 4.028518, 4.006023, 3.996498, 3.988161, 3.967935, 3.981896, 
    3.976389, 3.989496, 3.99784, 3.993711, 4.01923, 4.009298, 4.061803, 
    4.039135, 4.098388, 4.084161, 4.101802, 4.092794, 4.108238, 4.094337, 
    4.118433, 4.123693, 4.120099, 4.133912, 4.093567, 4.109035, 3.993596, 
    3.99427, 3.997406, 3.983632, 3.98279, 3.970192, 3.981399, 3.986179, 
    3.998323, 4.00552, 4.012367, 4.027449, 4.044335, 4.068018, 4.085083, 
    4.096546, 4.089513, 4.095722, 4.088782, 4.085532, 4.121723, 4.101378, 
    4.131923, 4.130229, 4.116393, 4.13042, 3.994742, 3.990869, 3.977444, 
    3.987948, 3.968821, 3.979522, 3.985684, 4.009508, 4.014751, 4.019621, 
    4.029246, 4.041622, 4.063388, 4.082383, 4.099768, 4.098493, 4.098942, 
    4.102833, 4.093201, 4.104415, 4.1063, 4.101374, 4.130002, 4.121811, 
    4.130193, 4.124858, 3.992127, 3.998646, 3.995123, 4.001751, 3.997082, 
    4.017873, 4.02412, 4.053425, 4.041378, 4.060557, 4.043323, 4.046374, 
    4.061189, 4.044252, 4.081337, 4.056177, 4.102984, 4.077784, 4.104567, 
    4.099693, 4.107762, 4.114999, 4.124112, 4.140963, 4.137057, 4.15117, 
    4.008377, 4.016856, 4.016107, 4.02499, 4.031568, 4.045845, 4.068811, 
    4.060164, 4.076044, 4.079237, 4.055114, 4.069918, 4.022535, 4.03017, 
    4.025621, 4.009047, 4.06216, 4.03485, 4.085365, 4.070504, 4.113967, 
    4.09232, 4.134908, 4.153202, 4.169961, 4.189597, 4.021486, 4.015719, 
    4.026046, 4.040366, 4.053673, 4.07141, 4.073226, 4.076556, 4.085186, 
    4.092451, 4.077612, 4.094274, 4.031948, 4.064534, 4.013543, 4.028859, 
    4.03952, 4.034839, 4.059176, 4.064927, 4.088346, 4.076227, 4.148685, 
    4.116533, 4.204576, 4.180165, 4.013706, 4.021465, 4.048544, 4.035645, 
    4.072595, 4.081722, 4.089149, 4.09866, 4.099685, 4.105327, 4.096085, 
    4.104961, 4.071448, 4.086403, 4.04544, 4.055388, 4.050809, 4.045792, 
    4.06129, 4.077846, 4.078196, 4.083514, 4.098531, 4.072744, 4.152853, 
    4.103276, 4.029936, 4.044932, 4.047072, 4.041258, 4.080807, 4.06645, 
    4.105189, 4.094696, 4.111896, 4.103344, 4.102087, 4.09112, 4.084302, 
    4.067109, 4.05315, 4.0421, 4.044668, 4.056811, 4.078859, 4.09978, 
    4.095192, 4.110587, 4.069909, 4.086938, 4.080352, 4.097537, 4.059936, 
    4.091955, 4.051778, 4.05529, 4.066165, 4.088098, 4.092953, 4.098149, 
    4.094942, 4.079419, 4.076877, 4.0659, 4.062874, 4.054524, 4.047622, 
    4.053929, 4.060561, 4.079423, 4.09647, 4.115103, 4.119669, 4.141531, 
    4.123735, 4.153131, 4.12814, 4.170937, 4.093809, 4.127398, 4.066659, 
    4.073175, 4.084982, 4.112131, 4.097456, 4.114619, 4.076777, 4.057233, 
    4.05218, 4.042772, 4.052395, 4.051612, 4.060833, 4.057868, 4.08005, 
    4.068126, 4.102057, 4.114482, 4.149691, 4.170851, 4.19233, 4.201837, 
    4.204732, 4.205943,
  3.282953, 3.30021, 3.29685, 3.310805, 3.303057, 3.312203, 3.286445, 
    3.300898, 3.291666, 3.284502, 3.338, 3.311428, 3.365734, 3.348682, 
    3.391619, 3.363079, 3.397393, 3.39079, 3.410678, 3.404972, 3.430499, 
    3.413313, 3.443773, 3.426387, 3.429105, 3.412747, 3.316761, 3.334685, 
    3.315701, 3.318253, 3.317107, 3.303219, 3.296236, 3.281634, 3.284281, 
    3.295007, 3.319401, 3.311105, 3.332032, 3.331558, 3.354958, 3.344394, 
    3.383881, 3.372627, 3.40521, 3.396997, 3.404825, 3.40245, 3.404856, 
    3.392816, 3.397971, 3.387388, 3.346372, 3.358394, 3.322623, 3.30124, 
    3.287079, 3.277056, 3.278472, 3.281173, 3.295069, 3.308167, 3.318172, 
    3.324877, 3.33149, 3.351571, 3.362224, 3.386161, 3.38183, 3.389167, 
    3.396181, 3.407982, 3.406038, 3.411244, 3.388971, 3.403764, 3.379365, 
    3.386028, 3.333302, 3.313341, 3.30489, 3.297496, 3.279561, 3.29194, 
    3.287057, 3.29868, 3.306081, 3.302419, 3.32506, 3.316246, 3.362856, 
    3.342727, 3.395362, 3.382718, 3.398397, 3.39039, 3.404118, 3.391761, 
    3.413182, 3.41786, 3.414663, 3.426948, 3.391078, 3.404826, 3.302317, 
    3.302914, 3.305696, 3.29348, 3.292733, 3.281562, 3.291499, 3.295738, 
    3.30651, 3.312894, 3.31897, 3.332354, 3.347344, 3.368376, 3.383537, 
    3.393725, 3.387475, 3.392992, 3.386825, 3.383936, 3.416107, 3.39802, 
    3.42518, 3.423673, 3.411369, 3.423842, 3.303333, 3.299898, 3.287992, 
    3.297307, 3.280347, 3.289835, 3.295299, 3.316433, 3.321085, 3.325406, 
    3.333949, 3.344935, 3.364264, 3.381139, 3.396589, 3.395455, 3.395854, 
    3.399313, 3.390752, 3.400719, 3.402395, 3.398016, 3.423471, 3.416186, 
    3.423641, 3.418896, 3.301014, 3.306797, 3.303671, 3.309551, 3.305409, 
    3.323855, 3.329399, 3.355415, 3.344719, 3.361749, 3.346445, 3.349154, 
    3.36231, 3.34727, 3.380209, 3.357859, 3.399447, 3.377052, 3.400854, 
    3.396522, 3.403695, 3.410129, 3.418233, 3.43322, 3.429746, 3.442302, 
    3.315429, 3.322953, 3.322288, 3.330171, 3.33601, 3.348684, 3.369081, 
    3.361401, 3.375506, 3.378343, 3.356916, 3.370064, 3.327993, 3.334769, 
    3.330732, 3.316023, 3.363173, 3.338923, 3.383789, 3.370585, 3.409212, 
    3.389969, 3.427834, 3.44411, 3.459462, 3.47747, 3.327062, 3.321944, 
    3.331109, 3.34382, 3.355636, 3.37139, 3.373003, 3.375961, 3.383629, 
    3.390085, 3.376899, 3.391705, 3.336346, 3.365282, 3.320013, 3.333605, 
    3.343069, 3.338913, 3.360523, 3.36563, 3.386436, 3.375669, 3.44009, 
    3.411493, 3.491214, 3.468819, 3.320158, 3.327043, 3.351081, 3.339629, 
    3.372442, 3.380551, 3.387151, 3.395603, 3.396515, 3.40153, 3.393315, 
    3.401205, 3.371423, 3.384711, 3.348325, 3.357159, 3.353093, 3.348637, 
    3.3624, 3.377107, 3.377418, 3.382143, 3.395489, 3.372575, 3.443799, 
    3.399706, 3.334562, 3.347874, 3.349774, 3.344612, 3.379738, 3.366984, 
    3.401407, 3.392081, 3.40737, 3.399767, 3.39865, 3.388903, 3.382844, 
    3.367568, 3.355171, 3.34536, 3.347639, 3.358423, 3.378007, 3.3966, 
    3.392522, 3.406206, 3.370056, 3.385186, 3.379334, 3.394606, 3.361198, 
    3.389644, 3.353953, 3.357071, 3.366731, 3.386216, 3.390532, 3.39515, 
    3.392299, 3.378505, 3.376246, 3.366495, 3.363807, 3.356392, 3.350262, 
    3.355863, 3.361753, 3.378509, 3.393657, 3.410222, 3.414282, 3.433725, 
    3.417897, 3.444046, 3.421814, 3.460354, 3.391292, 3.421154, 3.367169, 
    3.372958, 3.383448, 3.407579, 3.394534, 3.409791, 3.376158, 3.358797, 
    3.35431, 3.345957, 3.354501, 3.353806, 3.361994, 3.359361, 3.379066, 
    3.368472, 3.398623, 3.409669, 3.440986, 3.460277, 3.479978, 3.4887, 
    3.491358, 3.492469,
  2.997085, 3.014022, 3.010723, 3.024175, 3.016813, 3.025505, 3.000512, 
    3.014697, 3.005635, 2.998605, 3.05004, 3.024768, 3.076446, 3.060208, 
    3.101117, 3.073916, 3.106623, 3.100327, 3.119298, 3.113854, 3.138219, 
    3.121813, 3.1509, 3.134293, 3.136888, 3.121273, 3.029839, 3.046885, 
    3.028831, 3.031257, 3.030168, 3.016965, 3.01012, 2.995791, 2.998389, 
    3.008914, 3.032348, 3.024461, 3.044363, 3.043912, 3.066184, 3.056127, 
    3.093739, 3.083014, 3.114081, 3.106246, 3.113713, 3.111447, 3.113743, 
    3.102258, 3.107175, 3.097083, 3.058009, 3.069455, 3.035414, 3.015032, 
    3.001133, 2.991301, 2.992689, 2.995338, 3.008975, 3.021669, 3.031181, 
    3.037556, 3.043848, 3.062958, 3.073102, 3.095913, 3.091784, 3.098778, 
    3.105468, 3.116726, 3.11487, 3.119838, 3.098592, 3.112701, 3.089436, 
    3.095786, 3.045569, 3.026587, 3.018553, 3.011358, 2.993757, 3.005904, 
    3.001112, 3.012521, 3.019686, 3.016191, 3.037731, 3.029349, 3.073704, 
    3.05454, 3.104687, 3.092631, 3.107581, 3.099946, 3.113039, 3.101253, 
    3.121688, 3.126152, 3.123101, 3.13483, 3.100601, 3.113714, 3.016091, 
    3.016676, 3.01932, 3.007415, 3.006682, 2.99572, 3.005472, 3.009632, 
    3.020094, 3.026162, 3.031939, 3.044669, 3.058934, 3.078964, 3.093412, 
    3.103125, 3.097166, 3.102427, 3.096546, 3.093793, 3.124479, 3.107221, 
    3.133141, 3.131702, 3.119957, 3.131864, 3.017075, 3.013716, 3.00203, 
    3.011173, 2.994528, 3.003838, 3.009201, 3.029526, 3.033951, 3.03806, 
    3.046187, 3.056641, 3.075046, 3.091125, 3.105857, 3.104775, 3.105156, 
    3.108455, 3.10029, 3.109797, 3.111395, 3.107218, 3.131509, 3.124555, 
    3.131671, 3.127142, 3.014812, 3.020366, 3.017396, 3.022984, 3.019047, 
    3.036584, 3.041857, 3.066618, 3.056436, 3.07265, 3.058079, 3.060658, 
    3.073184, 3.058865, 3.090239, 3.068945, 3.108583, 3.087229, 3.109925, 
    3.105793, 3.112636, 3.118774, 3.126508, 3.140819, 3.137501, 3.149495, 
    3.028572, 3.035727, 3.035094, 3.042593, 3.048147, 3.060211, 3.079635, 
    3.072319, 3.085758, 3.088461, 3.068048, 3.080571, 3.04052, 3.046966, 
    3.043126, 3.029137, 3.074006, 3.050919, 3.093651, 3.081068, 3.117899, 
    3.099543, 3.135675, 3.151221, 3.165896, 3.18312, 3.039635, 3.034767, 
    3.043485, 3.05558, 3.066829, 3.081835, 3.083372, 3.086191, 3.093499, 
    3.099655, 3.087084, 3.101199, 3.048466, 3.076016, 3.03293, 3.045859, 
    3.054865, 3.05091, 3.071484, 3.076348, 3.096176, 3.085913, 3.147381, 
    3.120075, 3.196276, 3.174844, 3.033069, 3.039617, 3.062492, 3.051592, 
    3.082838, 3.090566, 3.096858, 3.104917, 3.105787, 3.11057, 3.102735, 
    3.110259, 3.081867, 3.094531, 3.059869, 3.06828, 3.064408, 3.060166, 
    3.073271, 3.087282, 3.087579, 3.092083, 3.104805, 3.082964, 3.150923, 
    3.108828, 3.04677, 3.059438, 3.061248, 3.056334, 3.08979, 3.077637, 
    3.110453, 3.101558, 3.116141, 3.108888, 3.107822, 3.098527, 3.092751, 
    3.078194, 3.066386, 3.057046, 3.059216, 3.069483, 3.08814, 3.105867, 
    3.101978, 3.115031, 3.080564, 3.094984, 3.089405, 3.103965, 3.072126, 
    3.099232, 3.065227, 3.068196, 3.077396, 3.095965, 3.10008, 3.104484, 
    3.101766, 3.088615, 3.086463, 3.077172, 3.074611, 3.067549, 3.061713, 
    3.067046, 3.072654, 3.088619, 3.103061, 3.118862, 3.122737, 3.1413, 
    3.126187, 3.151159, 3.129924, 3.166748, 3.100804, 3.129296, 3.077814, 
    3.083329, 3.093326, 3.11634, 3.103897, 3.118451, 3.086378, 3.069839, 
    3.065567, 3.057614, 3.065749, 3.065086, 3.072885, 3.070377, 3.08915, 
    3.079055, 3.107796, 3.118335, 3.148237, 3.166675, 3.185521, 3.19387, 
    3.196414, 3.197478,
  2.977282, 2.993935, 2.990691, 3.004174, 2.996686, 3.005526, 2.98065, 
    2.994599, 2.985687, 2.978777, 3.030506, 3.004776, 3.057181, 3.040874, 
    3.081588, 3.054681, 3.087042, 3.080806, 3.099605, 3.094208, 3.118379, 
    3.102099, 3.130979, 3.114483, 3.117059, 3.101563, 3.009936, 3.027292, 
    3.008911, 3.011379, 3.010271, 2.996842, 2.990097, 2.976012, 2.978564, 
    2.98891, 3.01249, 3.004465, 3.024724, 3.024266, 3.046971, 3.036714, 
    3.074285, 3.063675, 3.094433, 3.086669, 3.094068, 3.091822, 3.094097, 
    3.082719, 3.087589, 3.077595, 3.038632, 3.050273, 3.01561, 2.994929, 
    2.981261, 2.9716, 2.972964, 2.975566, 2.988971, 3.001625, 3.011302, 
    3.017792, 3.024199, 3.043678, 3.053877, 3.076436, 3.072351, 3.079273, 
    3.085898, 3.097054, 3.095215, 3.100141, 3.079089, 3.093065, 3.070027, 
    3.076311, 3.025951, 3.006627, 2.998455, 2.991314, 2.974013, 2.985951, 
    2.98124, 2.992459, 2.999609, 2.99607, 3.01797, 3.009438, 3.054471, 
    3.035095, 3.085124, 3.073189, 3.087992, 3.080429, 3.093399, 3.081724, 
    3.101975, 3.106403, 3.103376, 3.115015, 3.081078, 3.094069, 2.995971, 
    2.996548, 2.999236, 2.987437, 2.986716, 2.975942, 2.985526, 2.989617, 
    3.000023, 3.006195, 3.012074, 3.025036, 3.039576, 3.05967, 3.073961, 
    3.083578, 3.077677, 3.082886, 3.077064, 3.074338, 3.104743, 3.087635, 
    3.113338, 3.111911, 3.100258, 3.112071, 2.996953, 2.993635, 2.982142, 
    2.991132, 2.974771, 2.98392, 2.989193, 3.009618, 3.014121, 3.018305, 
    3.026582, 3.037238, 3.055798, 3.071698, 3.086283, 3.085212, 3.085589, 
    3.088857, 3.08077, 3.090187, 3.09177, 3.087632, 3.111719, 3.104819, 
    3.11188, 3.107385, 2.994713, 3.0003, 2.99728, 3.002962, 2.998958, 
    3.016802, 3.022171, 3.047414, 3.037028, 3.05343, 3.038704, 3.041334, 
    3.053957, 3.039505, 3.070821, 3.049769, 3.088984, 3.067843, 3.090314, 
    3.08622, 3.093, 3.099086, 3.106757, 3.120963, 3.117667, 3.129583, 
    3.008647, 3.015929, 3.015285, 3.022921, 3.02858, 3.040878, 3.060334, 
    3.053103, 3.066389, 3.069063, 3.048873, 3.061259, 3.02081, 3.027376, 
    3.023464, 3.009222, 3.05477, 3.031404, 3.074198, 3.061751, 3.098217, 
    3.08003, 3.115855, 3.131298, 3.145895, 3.163047, 3.019908, 3.014953, 
    3.02383, 3.036155, 3.047629, 3.062509, 3.064029, 3.066817, 3.074048, 
    3.080142, 3.0677, 3.081671, 3.028903, 3.056756, 3.013083, 3.026248, 
    3.035426, 3.031395, 3.052278, 3.057085, 3.076696, 3.066542, 3.127481, 
    3.100374, 3.176165, 3.154802, 3.013223, 3.01989, 3.043205, 3.03209, 
    3.063501, 3.071145, 3.077372, 3.085352, 3.086214, 3.090953, 3.083191, 
    3.090645, 3.062541, 3.075069, 3.040529, 3.04911, 3.045159, 3.040832, 
    3.054044, 3.067896, 3.068191, 3.072646, 3.085239, 3.063626, 3.131, 
    3.089225, 3.027176, 3.04009, 3.041936, 3.036925, 3.070378, 3.058359, 
    3.090837, 3.082026, 3.096475, 3.089287, 3.088231, 3.079025, 3.073308, 
    3.058909, 3.047178, 3.037651, 3.039863, 3.050301, 3.068745, 3.086293, 
    3.082441, 3.095375, 3.061253, 3.075516, 3.069997, 3.08441, 3.052912, 
    3.079721, 3.045995, 3.049025, 3.058121, 3.076488, 3.080563, 3.084924, 
    3.082232, 3.069214, 3.067086, 3.057899, 3.055368, 3.048365, 3.04241, 
    3.047851, 3.053434, 3.069219, 3.083514, 3.099173, 3.103016, 3.121439, 
    3.106436, 3.131235, 3.110144, 3.146741, 3.081278, 3.109521, 3.058534, 
    3.063987, 3.073876, 3.096671, 3.084342, 3.098764, 3.067002, 3.050652, 
    3.046342, 3.03823, 3.046527, 3.045851, 3.053662, 3.051185, 3.069744, 
    3.059761, 3.088205, 3.09865, 3.128333, 3.146669, 3.165441, 3.173765, 
    3.176302, 3.177364,
  2.975965, 2.994365, 2.990777, 3.005698, 2.997409, 3.007196, 2.979683, 
    2.995099, 2.985246, 2.977615, 3.03492, 3.006365, 3.064928, 3.046456, 
    3.093122, 3.062046, 3.099436, 3.092218, 3.114001, 3.107741, 3.135819, 
    3.116896, 3.150497, 3.131285, 3.134282, 3.116274, 3.012083, 3.031347, 
    3.010947, 3.013683, 3.012455, 2.99758, 2.99012, 2.974563, 2.97738, 
    2.988808, 3.014915, 3.00602, 3.028495, 3.027985, 3.053247, 3.041825, 
    3.084676, 3.07242, 3.108002, 3.099005, 3.107579, 3.104976, 3.107613, 
    3.094431, 3.10007, 3.088503, 3.04396, 3.056968, 3.018376, 2.995463, 
    2.980358, 2.969663, 2.971201, 2.974072, 2.988876, 3.002875, 3.013598, 
    3.020797, 3.027912, 3.049578, 3.061119, 3.087162, 3.08244, 3.090444, 
    3.098112, 3.111042, 3.108909, 3.114623, 3.090231, 3.106416, 3.079755, 
    3.087018, 3.029856, 3.008416, 2.999366, 2.991466, 2.972358, 2.985538, 
    2.980334, 2.992732, 3.000643, 2.996727, 3.020995, 3.011531, 3.061805, 
    3.040024, 3.097216, 3.083409, 3.100537, 3.091782, 3.106803, 3.09328, 
    3.116752, 3.121894, 3.118379, 3.131905, 3.092532, 3.107579, 2.996617, 
    2.997255, 3.000231, 2.98718, 2.986383, 2.974486, 2.985069, 2.98959, 
    3.001101, 3.007938, 3.014453, 3.028841, 3.04501, 3.067799, 3.084301, 
    3.095426, 3.088598, 3.094625, 3.087889, 3.084738, 3.119966, 3.100123, 
    3.129955, 3.128295, 3.114759, 3.128482, 2.997704, 2.994032, 2.981331, 
    2.991265, 2.973194, 2.983294, 2.98912, 3.01173, 3.016724, 3.021366, 
    3.030559, 3.042408, 3.063334, 3.081686, 3.098558, 3.097318, 3.097755, 
    3.101539, 3.092176, 3.10308, 3.104915, 3.10012, 3.128072, 3.120054, 
    3.128259, 3.123035, 2.995225, 3.001408, 2.998065, 3.004356, 2.999923, 
    3.019698, 3.025658, 3.05374, 3.042175, 3.060605, 3.04404, 3.046968, 
    3.061212, 3.044932, 3.080672, 3.056387, 3.101686, 3.077231, 3.103227, 
    3.098485, 3.106341, 3.113399, 3.122305, 3.138826, 3.13499, 3.148869, 
    3.010655, 3.018729, 3.018016, 3.026491, 3.032779, 3.04646, 3.068565, 
    3.060229, 3.075553, 3.078641, 3.055368, 3.069633, 3.024147, 3.03144, 
    3.027095, 3.011292, 3.062149, 3.035918, 3.084575, 3.0702, 3.112391, 
    3.09132, 3.132881, 3.150868, 3.167814, 3.187248, 3.023146, 3.017647, 
    3.027501, 3.041203, 3.053981, 3.071074, 3.072829, 3.076048, 3.084402, 
    3.091449, 3.077067, 3.093218, 3.033138, 3.064439, 3.015572, 3.030186, 
    3.040392, 3.035909, 3.059278, 3.064818, 3.087464, 3.07573, 3.146418, 
    3.114894, 3.202147, 3.177899, 3.015729, 3.023127, 3.049051, 3.036682, 
    3.072219, 3.081047, 3.088245, 3.09748, 3.098478, 3.103968, 3.094978, 
    3.103611, 3.071111, 3.085582, 3.046072, 3.055631, 3.051229, 3.046409, 
    3.061313, 3.077293, 3.077634, 3.082781, 3.097348, 3.072364, 3.15052, 
    3.101965, 3.031219, 3.045582, 3.047638, 3.04206, 3.08016, 3.066287, 
    3.103833, 3.093629, 3.11037, 3.102037, 3.100814, 3.090157, 3.083546, 
    3.066922, 3.053478, 3.042868, 3.045331, 3.056999, 3.078274, 3.098569, 
    3.094109, 3.109094, 3.069625, 3.086099, 3.07972, 3.096389, 3.060008, 
    3.090961, 3.052159, 3.055536, 3.066012, 3.087222, 3.091936, 3.096983, 
    3.093867, 3.078816, 3.076358, 3.065757, 3.062839, 3.054801, 3.048167, 
    3.054228, 3.060609, 3.078821, 3.095351, 3.113499, 3.11796, 3.13938, 
    3.121933, 3.150794, 3.12624, 3.16877, 3.092763, 3.125517, 3.066489, 
    3.07278, 3.084203, 3.110597, 3.09631, 3.113026, 3.076262, 3.057404, 
    3.052546, 3.043512, 3.052753, 3.052, 3.060873, 3.058018, 3.079428, 
    3.067904, 3.100783, 3.112893, 3.147411, 3.168689, 3.189965, 3.199419, 
    3.202303, 3.203511,
  3.255175, 3.278651, 3.274064, 3.293171, 3.282547, 3.295094, 3.25991, 
    3.279591, 3.267002, 3.257275, 3.330354, 3.294028, 3.368129, 3.344838, 
    3.403924, 3.364486, 3.411981, 3.402771, 3.430626, 3.422602, 3.458712, 
    3.434342, 3.477714, 3.452861, 3.456727, 3.433544, 3.301373, 3.325879, 
    3.299912, 3.30343, 3.30185, 3.282767, 3.273225, 3.253392, 3.256976, 
    3.27155, 3.305014, 3.293585, 3.32231, 3.321672, 3.353385, 3.339017, 
    3.393168, 3.377611, 3.422936, 3.41143, 3.422395, 3.419063, 3.422438, 
    3.405593, 3.412791, 3.398038, 3.3417, 3.358076, 3.30947, 3.280057, 
    3.260769, 3.247205, 3.249116, 3.252766, 3.271635, 3.28955, 3.303321, 
    3.312589, 3.32158, 3.348765, 3.363316, 3.396332, 3.390326, 3.40051, 
    3.41029, 3.426832, 3.424098, 3.431424, 3.400239, 3.420905, 3.386915, 
    3.396149, 3.324013, 3.296661, 3.285053, 3.274945, 3.250587, 3.267375, 
    3.260739, 3.276563, 3.286689, 3.281674, 3.312843, 3.300663, 3.364182, 
    3.336756, 3.409146, 3.391557, 3.413387, 3.402215, 3.421402, 3.404124, 
    3.434157, 3.440765, 3.436247, 3.45366, 3.403172, 3.422395, 3.281534, 
    3.282351, 3.286161, 3.26947, 3.268453, 3.253294, 3.266776, 3.272547, 
    3.287277, 3.296046, 3.304421, 3.322742, 3.343019, 3.37176, 3.392692, 
    3.406862, 3.398159, 3.40584, 3.397256, 3.393247, 3.438287, 3.412859, 
    3.451145, 3.449005, 3.431599, 3.449246, 3.282925, 3.278226, 3.262009, 
    3.274688, 3.25165, 3.264512, 3.271948, 3.300919, 3.307343, 3.313323, 
    3.324893, 3.33975, 3.366113, 3.389368, 3.41086, 3.409276, 3.409834, 
    3.414668, 3.402718, 3.416638, 3.418985, 3.412855, 3.448719, 3.4384, 
    3.44896, 3.442233, 3.279752, 3.28767, 3.283387, 3.29145, 3.285767, 
    3.311173, 3.318763, 3.354007, 3.339457, 3.362666, 3.3418, 3.34548, 
    3.363432, 3.342921, 3.388079, 3.357344, 3.414856, 3.383712, 3.416826, 
    3.410766, 3.42081, 3.429853, 3.441294, 3.462598, 3.457642, 3.475602, 
    3.299537, 3.309925, 3.309006, 3.319804, 3.327672, 3.344842, 3.372729, 
    3.362191, 3.381583, 3.385501, 3.356058, 3.37408, 3.316874, 3.325996, 
    3.320558, 3.300355, 3.364616, 3.331606, 3.393041, 3.374799, 3.428561, 
    3.401626, 3.45492, 3.478196, 3.500371, 3.526644, 3.315617, 3.308531, 
    3.321067, 3.338236, 3.35431, 3.375906, 3.37813, 3.38221, 3.39282, 
    3.40179, 3.383504, 3.404046, 3.328122, 3.36751, 3.305861, 3.324426, 
    3.337219, 3.331594, 3.36099, 3.36799, 3.396715, 3.381808, 3.472425, 
    3.431772, 3.54653, 3.513984, 3.306062, 3.315592, 3.348102, 3.332563, 
    3.377357, 3.388556, 3.39771, 3.409482, 3.410757, 3.417773, 3.40629, 
    3.417317, 3.375953, 3.39432, 3.344355, 3.35639, 3.350843, 3.344779, 
    3.363561, 3.38379, 3.384223, 3.39076, 3.409314, 3.37754, 3.477744, 
    3.415212, 3.325719, 3.343738, 3.346324, 3.339313, 3.38743, 3.369847, 
    3.417601, 3.404569, 3.425971, 3.415304, 3.413741, 3.400144, 3.391732, 
    3.37065, 3.353676, 3.340328, 3.343422, 3.358116, 3.385035, 3.410873, 
    3.405182, 3.424335, 3.374071, 3.394979, 3.38687, 3.40809, 3.361913, 
    3.401168, 3.352015, 3.356271, 3.3695, 3.396408, 3.402411, 3.408849, 
    3.404873, 3.385723, 3.382603, 3.369176, 3.365488, 3.355343, 3.346989, 
    3.354621, 3.362672, 3.38573, 3.406766, 3.429983, 3.435709, 3.463314, 
    3.440815, 3.478099, 3.446357, 3.501659, 3.403466, 3.445427, 3.370103, 
    3.378068, 3.392566, 3.426261, 3.40799, 3.429375, 3.382481, 3.358626, 
    3.352502, 3.341137, 3.352763, 3.351815, 3.363004, 3.359401, 3.3865, 
    3.371893, 3.413702, 3.429204, 3.473712, 3.50155, 3.53033, 3.542928, 
    3.546737, 3.548332,
  3.812404, 3.852935, 3.844963, 3.878335, 3.859724, 3.881718, 3.820526, 
    3.85457, 3.832741, 3.816003, 3.945439, 3.879842, 4.016918, 3.9726, 
    4.084901, 4.009933, 4.100402, 4.082692, 4.136672, 4.120995, 4.192386, 
    4.143967, 4.230846, 4.180668, 4.188405, 4.142399, 3.892797, 3.937107, 
    3.890216, 3.896439, 3.893642, 3.860107, 3.843508, 3.809351, 3.81549, 
    3.840605, 3.899246, 3.879063, 3.930481, 3.929299, 3.988772, 3.961649, 
    4.064366, 4.034974, 4.121646, 4.09934, 4.120591, 4.114113, 4.120676, 
    4.088104, 4.101967, 4.073641, 3.966691, 3.997692, 3.907158, 3.855382, 
    3.822003, 3.79879, 3.802049, 3.808282, 3.840753, 3.871976, 3.896244, 
    3.912714, 3.929129, 3.980018, 4.007694, 4.070388, 4.058969, 4.078364, 
    4.097141, 4.129246, 4.12391, 4.138237, 4.077846, 4.117693, 4.052508, 
    4.070038, 3.93364, 3.884479, 3.864102, 3.846492, 3.804559, 3.833384, 
    3.821951, 3.849302, 3.866964, 3.8582, 3.913167, 3.891543, 4.009351, 
    3.957408, 4.094938, 4.061305, 4.103119, 4.081626, 4.118659, 4.085286, 
    4.143604, 4.156631, 4.147717, 4.182266, 4.083459, 4.120593, 3.857956, 
    3.859382, 3.86604, 3.837005, 3.835248, 3.809184, 3.83235, 3.842334, 
    3.867993, 3.883395, 3.898193, 3.931283, 3.969174, 4.0239, 4.063461, 
    4.090542, 4.073873, 4.088579, 4.07215, 4.064516, 4.151737, 4.102098, 
    4.177245, 4.17298, 4.13858, 4.17346, 3.860383, 3.852195, 3.824135, 
    3.846047, 3.806375, 3.828445, 3.841295, 3.891995, 3.903378, 3.914021, 
    3.935274, 3.963025, 4.013051, 4.057152, 4.09824, 4.095188, 4.096262, 
    4.105596, 4.08259, 4.109409, 4.113963, 4.102091, 4.17241, 4.15196, 
    4.172889, 4.159536, 3.854851, 3.868681, 3.861192, 3.87531, 3.86535, 
    3.910189, 3.923914, 3.989952, 3.962475, 4.006453, 3.966879, 3.973813, 
    4.007917, 3.968989, 4.054711, 3.996297, 4.10596, 4.046457, 4.109775, 
    4.09806, 4.117507, 4.135158, 4.157678, 4.200199, 4.190238, 4.22654, 
    3.889553, 3.907968, 3.906334, 3.925841, 3.940442, 3.972609, 4.025767, 
    4.005544, 4.042443, 4.049835, 3.993851, 4.028355, 3.920425, 3.937325, 
    3.927237, 3.890998, 4.010183, 3.947774, 4.064123, 4.0297, 4.132628, 
    4.080499, 4.184785, 4.23183, 4.277549, 4.332258, 3.918117, 3.905489, 
    3.928178, 3.960184, 3.990528, 4.031776, 4.035948, 4.043625, 4.063704, 
    4.080814, 4.046064, 4.085135, 3.941279, 4.01573, 3.900746, 3.934408, 
    3.958276, 3.947753, 4.00325, 4.016651, 4.071118, 4.042867, 4.220077, 
    4.138919, 4.374618, 4.306069, 3.901104, 3.918072, 3.978763, 3.949563, 
    4.034496, 4.055614, 4.073015, 4.095585, 4.098041, 4.11161, 4.089443, 
    4.110727, 4.031862, 4.066557, 3.97169, 3.994482, 3.983951, 3.972489, 
    4.008162, 4.046605, 4.047421, 4.059792, 4.095261, 4.034841, 4.230908, 
    4.106648, 3.93681, 3.970529, 3.975405, 3.962204, 4.053482, 4.020219, 
    4.111277, 4.08614, 4.127563, 4.106827, 4.103803, 4.077665, 4.061636, 
    4.021764, 3.989324, 3.96411, 3.969933, 3.997768, 4.048954, 4.098266, 
    4.087316, 4.124372, 4.028337, 4.067811, 4.052423, 4.092905, 4.005012, 
    4.079624, 3.986172, 3.994256, 4.019552, 4.070532, 4.082003, 4.094365, 
    4.086723, 4.050254, 4.044367, 4.01893, 4.011853, 3.992491, 3.97666, 
    3.991119, 4.006463, 4.050267, 4.090358, 4.135411, 4.146657, 4.201643, 
    4.15673, 4.231632, 4.167714, 4.280233, 4.084023, 4.165866, 4.020712, 
    4.035832, 4.063222, 4.128131, 4.092711, 4.134221, 4.044136, 3.998741, 
    3.987096, 3.965631, 3.987591, 3.985792, 4.007099, 4.000217, 4.051724, 
    4.024157, 4.103728, 4.133887, 4.222694, 4.280007, 4.339907, 4.366786, 
    4.375068, 4.378545,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24856.9, 24877.73, 24873.65, 24890.69, 24881.21, 24892.41, 24861.09, 
    24878.57, 24867.38, 24858.76, 24924.51, 24891.46, 24959.89, 24938.02, 
    24993.41, 24956.46, 25001, 24992.32, 25018.67, 25011.05, 25045.57, 
    25022.21, 25063.97, 25039.94, 25043.66, 25021.45, 24898.04, 24920.35, 
    24896.73, 24899.88, 24898.46, 24881.4, 24872.9, 24855.33, 24858.49, 
    24871.42, 24901.3, 24891.06, 24917.04, 24916.45, 24946.03, 24932.58, 
    24983.31, 24968.79, 25011.37, 25000.48, 25010.85, 25007.7, 25010.89, 
    24994.98, 25001.77, 24987.88, 24935.09, 24950.44, 24905.31, 24878.99, 
    24861.85, 24849.86, 24851.55, 24854.77, 24871.49, 24887.46, 24899.78, 
    24908.12, 24916.36, 24941.7, 24955.36, 24986.28, 24980.65, 24990.2, 
    24999.4, 25015.06, 25012.47, 25019.43, 24989.94, 25009.44, 24977.46, 
    24986.11, 24918.62, 24893.81, 24883.44, 24874.44, 24852.85, 24867.71, 
    24861.82, 24875.88, 24884.9, 24880.43, 24908.35, 24897.4, 24956.18, 
    24930.47, 24998.33, 24981.8, 25002.33, 24991.8, 25009.91, 24993.6, 
    25022.04, 25028.34, 25024.03, 25040.71, 24992.7, 25010.85, 24880.3, 
    24881.03, 24884.43, 24869.57, 24868.66, 24855.24, 24867.18, 24872.3, 
    24885.43, 24893.26, 24900.77, 24917.44, 24936.32, 24963.32, 24982.87, 
    24996.17, 24987.99, 24995.21, 24987.14, 24983.39, 25025.98, 25001.83, 
    25038.29, 25036.24, 25019.6, 25036.47, 24881.54, 24877.36, 24862.95, 
    24874.21, 24853.79, 24865.17, 24871.77, 24897.63, 24903.4, 24908.78, 
    24919.44, 24933.27, 24957.99, 24979.76, 24999.94, 24998.45, 24998.97, 
    25003.54, 24992.27, 25005.4, 25007.62, 25001.83, 25035.96, 25026.08, 
    25036.19, 25029.75, 24878.71, 24885.78, 24881.96, 24889.15, 24884.08, 
    24906.84, 24913.75, 24946.62, 24932.99, 24954.75, 24935.18, 24938.62, 
    24955.47, 24936.23, 24978.55, 24949.75, 25003.72, 24974.47, 25005.58, 
    24999.85, 25009.35, 25017.94, 25028.85, 25049.32, 25044.54, 25061.92, 
    24896.39, 24905.72, 24904.89, 24914.72, 24922.02, 24938.03, 24964.23, 
    24954.3, 24972.49, 24976.14, 24948.54, 24965.51, 24912, 24920.46, 
    24915.41, 24897.12, 24956.59, 24925.68, 24983.19, 24966.17, 25016.71, 
    24991.25, 25041.92, 25064.44, 25086.12, 25111.87, 24910.84, 24904.46, 
    24915.89, 24931.85, 24946.9, 24967.2, 24969.27, 24973.07, 24982.99, 
    24991.4, 24974.28, 24993.52, 24922.44, 24959.31, 24902.06, 24919, 
    24930.9, 24925.66, 24953.17, 24959.76, 24986.64, 24972.7, 25058.83, 
    25019.76, 25131.71, 25099.51, 24902.25, 24910.82, 24941.08, 24926.57, 
    24968.55, 24979, 24987.57, 24998.64, 24999.85, 25006.47, 24995.63, 
    25006.04, 24967.25, 24984.39, 24937.57, 24948.85, 24943.65, 24937.97, 
    24955.59, 24974.55, 24974.95, 24981.06, 24998.48, 24968.72, 25064, 
    25004.05, 24920.2, 24936.99, 24939.41, 24932.86, 24977.95, 24961.51, 
    25006.31, 24994.02, 25014.25, 25004.14, 25002.66, 24989.86, 24981.97, 
    24962.27, 24946.3, 24933.81, 24936.7, 24950.47, 24975.71, 24999.96, 
    24994.59, 25012.69, 24965.5, 24985.01, 24977.42, 24997.33, 24954.04, 
    24990.82, 24944.75, 24948.74, 24961.19, 24986.35, 24991.98, 24998.04, 
    24994.3, 24976.35, 24973.44, 24960.88, 24957.41, 24947.87, 24940.04, 
    24947.19, 24954.76, 24976.36, 24996.08, 25018.06, 25023.52, 25050.02, 
    25028.39, 25064.35, 25033.7, 25087.38, 24992.98, 25032.81, 24961.76, 
    24969.21, 24982.75, 25014.52, 24997.24, 25017.48, 24973.33, 24950.95, 
    24945.2, 24934.56, 24945.45, 24944.56, 24955.07, 24951.68, 24977.08, 
    24963.45, 25002.62, 25017.32, 25060.08, 25087.27, 25115.48, 25128.06, 
    25131.91, 25133.53 ;

 HCSOI =
  24856.9, 24877.73, 24873.65, 24890.69, 24881.21, 24892.41, 24861.09, 
    24878.57, 24867.38, 24858.76, 24924.51, 24891.46, 24959.89, 24938.02, 
    24993.41, 24956.46, 25001, 24992.32, 25018.67, 25011.05, 25045.57, 
    25022.21, 25063.97, 25039.94, 25043.66, 25021.45, 24898.04, 24920.35, 
    24896.73, 24899.88, 24898.46, 24881.4, 24872.9, 24855.33, 24858.49, 
    24871.42, 24901.3, 24891.06, 24917.04, 24916.45, 24946.03, 24932.58, 
    24983.31, 24968.79, 25011.37, 25000.48, 25010.85, 25007.7, 25010.89, 
    24994.98, 25001.77, 24987.88, 24935.09, 24950.44, 24905.31, 24878.99, 
    24861.85, 24849.86, 24851.55, 24854.77, 24871.49, 24887.46, 24899.78, 
    24908.12, 24916.36, 24941.7, 24955.36, 24986.28, 24980.65, 24990.2, 
    24999.4, 25015.06, 25012.47, 25019.43, 24989.94, 25009.44, 24977.46, 
    24986.11, 24918.62, 24893.81, 24883.44, 24874.44, 24852.85, 24867.71, 
    24861.82, 24875.88, 24884.9, 24880.43, 24908.35, 24897.4, 24956.18, 
    24930.47, 24998.33, 24981.8, 25002.33, 24991.8, 25009.91, 24993.6, 
    25022.04, 25028.34, 25024.03, 25040.71, 24992.7, 25010.85, 24880.3, 
    24881.03, 24884.43, 24869.57, 24868.66, 24855.24, 24867.18, 24872.3, 
    24885.43, 24893.26, 24900.77, 24917.44, 24936.32, 24963.32, 24982.87, 
    24996.17, 24987.99, 24995.21, 24987.14, 24983.39, 25025.98, 25001.83, 
    25038.29, 25036.24, 25019.6, 25036.47, 24881.54, 24877.36, 24862.95, 
    24874.21, 24853.79, 24865.17, 24871.77, 24897.63, 24903.4, 24908.78, 
    24919.44, 24933.27, 24957.99, 24979.76, 24999.94, 24998.45, 24998.97, 
    25003.54, 24992.27, 25005.4, 25007.62, 25001.83, 25035.96, 25026.08, 
    25036.19, 25029.75, 24878.71, 24885.78, 24881.96, 24889.15, 24884.08, 
    24906.84, 24913.75, 24946.62, 24932.99, 24954.75, 24935.18, 24938.62, 
    24955.47, 24936.23, 24978.55, 24949.75, 25003.72, 24974.47, 25005.58, 
    24999.85, 25009.35, 25017.94, 25028.85, 25049.32, 25044.54, 25061.92, 
    24896.39, 24905.72, 24904.89, 24914.72, 24922.02, 24938.03, 24964.23, 
    24954.3, 24972.49, 24976.14, 24948.54, 24965.51, 24912, 24920.46, 
    24915.41, 24897.12, 24956.59, 24925.68, 24983.19, 24966.17, 25016.71, 
    24991.25, 25041.92, 25064.44, 25086.12, 25111.87, 24910.84, 24904.46, 
    24915.89, 24931.85, 24946.9, 24967.2, 24969.27, 24973.07, 24982.99, 
    24991.4, 24974.28, 24993.52, 24922.44, 24959.31, 24902.06, 24919, 
    24930.9, 24925.66, 24953.17, 24959.76, 24986.64, 24972.7, 25058.83, 
    25019.76, 25131.71, 25099.51, 24902.25, 24910.82, 24941.08, 24926.57, 
    24968.55, 24979, 24987.57, 24998.64, 24999.85, 25006.47, 24995.63, 
    25006.04, 24967.25, 24984.39, 24937.57, 24948.85, 24943.65, 24937.97, 
    24955.59, 24974.55, 24974.95, 24981.06, 24998.48, 24968.72, 25064, 
    25004.05, 24920.2, 24936.99, 24939.41, 24932.86, 24977.95, 24961.51, 
    25006.31, 24994.02, 25014.25, 25004.14, 25002.66, 24989.86, 24981.97, 
    24962.27, 24946.3, 24933.81, 24936.7, 24950.47, 24975.71, 24999.96, 
    24994.59, 25012.69, 24965.5, 24985.01, 24977.42, 24997.33, 24954.04, 
    24990.82, 24944.75, 24948.74, 24961.19, 24986.35, 24991.98, 24998.04, 
    24994.3, 24976.35, 24973.44, 24960.88, 24957.41, 24947.87, 24940.04, 
    24947.19, 24954.76, 24976.36, 24996.08, 25018.06, 25023.52, 25050.02, 
    25028.39, 25064.35, 25033.7, 25087.38, 24992.98, 25032.81, 24961.76, 
    24969.21, 24982.75, 25014.52, 24997.24, 25017.48, 24973.33, 24950.95, 
    24945.2, 24934.56, 24945.45, 24944.56, 24955.07, 24951.68, 24977.08, 
    24963.45, 25002.62, 25017.32, 25060.08, 25087.27, 25115.48, 25128.06, 
    25131.91, 25133.53 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 HR_vr =
  2.694543e-07, 2.70184e-07, 2.700423e-07, 2.706303e-07, 2.703043e-07, 
    2.706891e-07, 2.696024e-07, 2.702129e-07, 2.698233e-07, 2.695202e-07, 
    2.717696e-07, 2.706565e-07, 2.729249e-07, 2.722163e-07, 2.739952e-07, 
    2.728145e-07, 2.74233e-07, 2.739614e-07, 2.747792e-07, 2.74545e-07, 
    2.755894e-07, 2.748872e-07, 2.761305e-07, 2.754219e-07, 2.755327e-07, 
    2.74864e-07, 2.708809e-07, 2.716311e-07, 2.708364e-07, 2.709434e-07, 
    2.708954e-07, 2.703109e-07, 2.70016e-07, 2.693987e-07, 2.695108e-07, 
    2.699643e-07, 2.709916e-07, 2.706432e-07, 2.715213e-07, 2.715015e-07, 
    2.724776e-07, 2.720377e-07, 2.736763e-07, 2.73211e-07, 2.745548e-07, 
    2.742171e-07, 2.745389e-07, 2.744414e-07, 2.745402e-07, 2.740448e-07, 
    2.742571e-07, 2.738211e-07, 2.7212e-07, 2.726204e-07, 2.711269e-07, 
    2.70227e-07, 2.696292e-07, 2.692045e-07, 2.692645e-07, 2.693789e-07, 
    2.69967e-07, 2.705196e-07, 2.709403e-07, 2.712216e-07, 2.714986e-07, 
    2.723359e-07, 2.727792e-07, 2.737702e-07, 2.735917e-07, 2.738943e-07, 
    2.741835e-07, 2.746685e-07, 2.745887e-07, 2.748023e-07, 2.738865e-07, 
    2.744952e-07, 2.734899e-07, 2.73765e-07, 2.715731e-07, 2.707372e-07, 
    2.703809e-07, 2.700695e-07, 2.693107e-07, 2.698348e-07, 2.696282e-07, 
    2.701197e-07, 2.704317e-07, 2.702774e-07, 2.712293e-07, 2.708593e-07, 
    2.728055e-07, 2.719679e-07, 2.741498e-07, 2.736284e-07, 2.742747e-07, 
    2.73945e-07, 2.745098e-07, 2.740015e-07, 2.748818e-07, 2.750732e-07, 
    2.749424e-07, 2.754451e-07, 2.739733e-07, 2.745388e-07, 2.702731e-07, 
    2.702982e-07, 2.704155e-07, 2.698998e-07, 2.698683e-07, 2.693956e-07, 
    2.698163e-07, 2.699953e-07, 2.704498e-07, 2.707184e-07, 2.709737e-07, 
    2.715346e-07, 2.721604e-07, 2.730347e-07, 2.736622e-07, 2.740824e-07, 
    2.738248e-07, 2.740522e-07, 2.73798e-07, 2.736788e-07, 2.750014e-07, 
    2.74259e-07, 2.753728e-07, 2.753112e-07, 2.748073e-07, 2.753182e-07, 
    2.703159e-07, 2.701711e-07, 2.696679e-07, 2.700617e-07, 2.693441e-07, 
    2.697458e-07, 2.699766e-07, 2.708669e-07, 2.710626e-07, 2.712437e-07, 
    2.716014e-07, 2.720602e-07, 2.728641e-07, 2.73563e-07, 2.742004e-07, 
    2.741537e-07, 2.741701e-07, 2.743124e-07, 2.739599e-07, 2.743702e-07, 
    2.74439e-07, 2.74259e-07, 2.75303e-07, 2.750049e-07, 2.753099e-07, 
    2.751159e-07, 2.702182e-07, 2.704619e-07, 2.703302e-07, 2.705777e-07, 
    2.704033e-07, 2.711784e-07, 2.714106e-07, 2.724963e-07, 2.720511e-07, 
    2.727597e-07, 2.721232e-07, 2.72236e-07, 2.727824e-07, 2.721576e-07, 
    2.735243e-07, 2.725978e-07, 2.743179e-07, 2.733935e-07, 2.743757e-07, 
    2.741976e-07, 2.744926e-07, 2.747566e-07, 2.750887e-07, 2.757008e-07, 
    2.755591e-07, 2.760708e-07, 2.70825e-07, 2.711407e-07, 2.71113e-07, 
    2.714434e-07, 2.716875e-07, 2.722165e-07, 2.73064e-07, 2.727455e-07, 
    2.733303e-07, 2.734476e-07, 2.725592e-07, 2.731046e-07, 2.71352e-07, 
    2.716353e-07, 2.714667e-07, 2.708498e-07, 2.728187e-07, 2.718089e-07, 
    2.736725e-07, 2.731264e-07, 2.747189e-07, 2.739273e-07, 2.754811e-07, 
    2.761438e-07, 2.767675e-07, 2.774948e-07, 2.713131e-07, 2.710986e-07, 
    2.714827e-07, 2.720134e-07, 2.725058e-07, 2.731597e-07, 2.732266e-07, 
    2.73349e-07, 2.736661e-07, 2.739324e-07, 2.733876e-07, 2.739992e-07, 
    2.717007e-07, 2.729064e-07, 2.710174e-07, 2.715866e-07, 2.719821e-07, 
    2.718088e-07, 2.727091e-07, 2.729211e-07, 2.737817e-07, 2.73337e-07, 
    2.759802e-07, 2.748121e-07, 2.780485e-07, 2.771457e-07, 2.710237e-07, 
    2.713124e-07, 2.723161e-07, 2.718388e-07, 2.732034e-07, 2.735388e-07, 
    2.738115e-07, 2.741596e-07, 2.741973e-07, 2.744035e-07, 2.740655e-07, 
    2.743902e-07, 2.731611e-07, 2.737107e-07, 2.722016e-07, 2.725692e-07, 
    2.724002e-07, 2.722146e-07, 2.72787e-07, 2.733961e-07, 2.734093e-07, 
    2.736045e-07, 2.741536e-07, 2.732089e-07, 2.761303e-07, 2.743273e-07, 
    2.716271e-07, 2.721823e-07, 2.722619e-07, 2.720468e-07, 2.735052e-07, 
    2.729771e-07, 2.743985e-07, 2.740147e-07, 2.746435e-07, 2.743311e-07, 
    2.742851e-07, 2.738837e-07, 2.736336e-07, 2.730013e-07, 2.724865e-07, 
    2.72078e-07, 2.721731e-07, 2.726216e-07, 2.734334e-07, 2.742006e-07, 
    2.740326e-07, 2.745957e-07, 2.731045e-07, 2.737301e-07, 2.734883e-07, 
    2.741186e-07, 2.72737e-07, 2.73913e-07, 2.72436e-07, 2.725656e-07, 
    2.729666e-07, 2.737723e-07, 2.739508e-07, 2.741409e-07, 2.740237e-07, 
    2.73454e-07, 2.733608e-07, 2.72957e-07, 2.728453e-07, 2.725374e-07, 
    2.722823e-07, 2.725154e-07, 2.727599e-07, 2.734544e-07, 2.740794e-07, 
    2.747603e-07, 2.749269e-07, 2.757207e-07, 2.750743e-07, 2.761403e-07, 
    2.752336e-07, 2.768026e-07, 2.739814e-07, 2.752074e-07, 2.729849e-07, 
    2.732248e-07, 2.736581e-07, 2.746515e-07, 2.741157e-07, 2.747424e-07, 
    2.733571e-07, 2.72637e-07, 2.724508e-07, 2.721029e-07, 2.724587e-07, 
    2.724298e-07, 2.727702e-07, 2.726609e-07, 2.734774e-07, 2.730389e-07, 
    2.742839e-07, 2.747375e-07, 2.760171e-07, 2.768001e-07, 2.775965e-07, 
    2.779476e-07, 2.780545e-07, 2.780991e-07,
  2.336853e-07, 2.345734e-07, 2.344009e-07, 2.351167e-07, 2.347197e-07, 
    2.351883e-07, 2.338655e-07, 2.346086e-07, 2.341343e-07, 2.337654e-07, 
    2.365042e-07, 2.351486e-07, 2.37911e-07, 2.370478e-07, 2.392149e-07, 
    2.377766e-07, 2.395046e-07, 2.391736e-07, 2.401701e-07, 2.398847e-07, 
    2.411577e-07, 2.403017e-07, 2.418172e-07, 2.409535e-07, 2.410886e-07, 
    2.402735e-07, 2.354218e-07, 2.363355e-07, 2.353676e-07, 2.354979e-07, 
    2.354395e-07, 2.347279e-07, 2.34369e-07, 2.336175e-07, 2.33754e-07, 
    2.34306e-07, 2.355565e-07, 2.351323e-07, 2.362014e-07, 2.361773e-07, 
    2.373661e-07, 2.368302e-07, 2.388263e-07, 2.382594e-07, 2.398966e-07, 
    2.394851e-07, 2.398773e-07, 2.397584e-07, 2.398788e-07, 2.392753e-07, 
    2.395339e-07, 2.390027e-07, 2.369306e-07, 2.3754e-07, 2.357213e-07, 
    2.346259e-07, 2.338981e-07, 2.333811e-07, 2.334542e-07, 2.335935e-07, 
    2.343092e-07, 2.349818e-07, 2.35494e-07, 2.358365e-07, 2.361738e-07, 
    2.371937e-07, 2.377335e-07, 2.389407e-07, 2.387231e-07, 2.390919e-07, 
    2.394442e-07, 2.400352e-07, 2.39938e-07, 2.401983e-07, 2.390823e-07, 
    2.39824e-07, 2.385991e-07, 2.389343e-07, 2.362649e-07, 2.352468e-07, 
    2.348132e-07, 2.34434e-07, 2.335104e-07, 2.341483e-07, 2.338969e-07, 
    2.344951e-07, 2.348749e-07, 2.346871e-07, 2.358458e-07, 2.353955e-07, 
    2.377655e-07, 2.367454e-07, 2.394031e-07, 2.387678e-07, 2.395553e-07, 
    2.391536e-07, 2.398418e-07, 2.392225e-07, 2.402952e-07, 2.405285e-07, 
    2.40369e-07, 2.409816e-07, 2.391881e-07, 2.398772e-07, 2.346818e-07, 
    2.347124e-07, 2.348552e-07, 2.342275e-07, 2.341891e-07, 2.336137e-07, 
    2.341258e-07, 2.343437e-07, 2.348969e-07, 2.352239e-07, 2.355347e-07, 
    2.362177e-07, 2.369798e-07, 2.380446e-07, 2.38809e-07, 2.39321e-07, 
    2.390071e-07, 2.392842e-07, 2.389745e-07, 2.388292e-07, 2.40441e-07, 
    2.395363e-07, 2.408935e-07, 2.408185e-07, 2.402044e-07, 2.40827e-07, 
    2.347339e-07, 2.345576e-07, 2.339451e-07, 2.344245e-07, 2.33551e-07, 
    2.3404e-07, 2.34321e-07, 2.354048e-07, 2.356429e-07, 2.358634e-07, 
    2.36299e-07, 2.368577e-07, 2.378369e-07, 2.386882e-07, 2.394647e-07, 
    2.394079e-07, 2.394279e-07, 2.396012e-07, 2.391717e-07, 2.396717e-07, 
    2.397555e-07, 2.395362e-07, 2.408085e-07, 2.404452e-07, 2.408169e-07, 
    2.405804e-07, 2.34615e-07, 2.349116e-07, 2.347513e-07, 2.350527e-07, 
    2.348403e-07, 2.35784e-07, 2.360667e-07, 2.373889e-07, 2.368466e-07, 
    2.377097e-07, 2.369344e-07, 2.370718e-07, 2.377376e-07, 2.369763e-07, 
    2.386411e-07, 2.375126e-07, 2.396079e-07, 2.384818e-07, 2.396784e-07, 
    2.394613e-07, 2.398208e-07, 2.401426e-07, 2.405473e-07, 2.412934e-07, 
    2.411207e-07, 2.417445e-07, 2.353537e-07, 2.357381e-07, 2.357043e-07, 
    2.361065e-07, 2.364038e-07, 2.370481e-07, 2.380803e-07, 2.376923e-07, 
    2.384047e-07, 2.385476e-07, 2.374654e-07, 2.381299e-07, 2.359953e-07, 
    2.363404e-07, 2.36135e-07, 2.353839e-07, 2.377816e-07, 2.365518e-07, 
    2.388216e-07, 2.381563e-07, 2.400967e-07, 2.391321e-07, 2.410256e-07, 
    2.418336e-07, 2.425939e-07, 2.43481e-07, 2.359479e-07, 2.356868e-07, 
    2.361544e-07, 2.368007e-07, 2.374004e-07, 2.381969e-07, 2.382784e-07, 
    2.384275e-07, 2.388137e-07, 2.391383e-07, 2.384745e-07, 2.392196e-07, 
    2.364202e-07, 2.378883e-07, 2.355879e-07, 2.362811e-07, 2.367627e-07, 
    2.365516e-07, 2.37648e-07, 2.379062e-07, 2.389547e-07, 2.384129e-07, 
    2.416342e-07, 2.402103e-07, 2.441562e-07, 2.430552e-07, 2.355955e-07, 
    2.359471e-07, 2.371694e-07, 2.36588e-07, 2.382501e-07, 2.386587e-07, 
    2.389909e-07, 2.394151e-07, 2.39461e-07, 2.397123e-07, 2.393004e-07, 
    2.39696e-07, 2.381986e-07, 2.388681e-07, 2.370299e-07, 2.374776e-07, 
    2.372717e-07, 2.370458e-07, 2.377429e-07, 2.384849e-07, 2.38501e-07, 
    2.387387e-07, 2.394081e-07, 2.382568e-07, 2.418174e-07, 2.396198e-07, 
    2.363303e-07, 2.370065e-07, 2.371033e-07, 2.368414e-07, 2.386178e-07, 
    2.379745e-07, 2.397061e-07, 2.392385e-07, 2.400047e-07, 2.39624e-07, 
    2.39568e-07, 2.390788e-07, 2.387742e-07, 2.380039e-07, 2.373769e-07, 
    2.368794e-07, 2.369951e-07, 2.375415e-07, 2.385304e-07, 2.39465e-07, 
    2.392604e-07, 2.399465e-07, 2.381297e-07, 2.388918e-07, 2.385973e-07, 
    2.393652e-07, 2.37682e-07, 2.391149e-07, 2.373153e-07, 2.374733e-07, 
    2.379617e-07, 2.389434e-07, 2.391607e-07, 2.393923e-07, 2.392494e-07, 
    2.385555e-07, 2.384418e-07, 2.379499e-07, 2.378139e-07, 2.374389e-07, 
    2.371282e-07, 2.37412e-07, 2.3771e-07, 2.385559e-07, 2.393174e-07, 
    2.401471e-07, 2.403501e-07, 2.413179e-07, 2.405299e-07, 2.418296e-07, 
    2.407244e-07, 2.426369e-07, 2.391982e-07, 2.406922e-07, 2.37984e-07, 
    2.382762e-07, 2.388042e-07, 2.400146e-07, 2.393616e-07, 2.401254e-07, 
    2.384374e-07, 2.375602e-07, 2.373334e-07, 2.369096e-07, 2.373431e-07, 
    2.373078e-07, 2.377224e-07, 2.375892e-07, 2.385839e-07, 2.380498e-07, 
    2.395665e-07, 2.401194e-07, 2.416791e-07, 2.426337e-07, 2.436048e-07, 
    2.440331e-07, 2.441634e-07, 2.442178e-07,
  2.190408e-07, 2.200111e-07, 2.198226e-07, 2.206048e-07, 2.20171e-07, 
    2.206831e-07, 2.192376e-07, 2.200496e-07, 2.195313e-07, 2.191283e-07, 
    2.221216e-07, 2.206397e-07, 2.236599e-07, 2.227158e-07, 2.250865e-07, 
    2.23513e-07, 2.254036e-07, 2.250412e-07, 2.261318e-07, 2.258195e-07, 
    2.272133e-07, 2.26276e-07, 2.279356e-07, 2.269896e-07, 2.271376e-07, 
    2.26245e-07, 2.209381e-07, 2.219371e-07, 2.208789e-07, 2.210214e-07, 
    2.209575e-07, 2.201799e-07, 2.197878e-07, 2.189667e-07, 2.191158e-07, 
    2.197189e-07, 2.210855e-07, 2.206218e-07, 2.217903e-07, 2.21764e-07, 
    2.230639e-07, 2.224779e-07, 2.246612e-07, 2.24041e-07, 2.258325e-07, 
    2.253822e-07, 2.258114e-07, 2.256812e-07, 2.258131e-07, 2.251525e-07, 
    2.254355e-07, 2.248542e-07, 2.225876e-07, 2.23254e-07, 2.212656e-07, 
    2.200685e-07, 2.192732e-07, 2.187086e-07, 2.187884e-07, 2.189406e-07, 
    2.197225e-07, 2.204573e-07, 2.210171e-07, 2.213914e-07, 2.217602e-07, 
    2.228755e-07, 2.234658e-07, 2.247865e-07, 2.245483e-07, 2.249518e-07, 
    2.253373e-07, 2.259843e-07, 2.258778e-07, 2.261627e-07, 2.249413e-07, 
    2.257531e-07, 2.244126e-07, 2.247794e-07, 2.2186e-07, 2.207469e-07, 
    2.202733e-07, 2.198588e-07, 2.188498e-07, 2.195466e-07, 2.19272e-07, 
    2.199254e-07, 2.203405e-07, 2.201352e-07, 2.214017e-07, 2.209094e-07, 
    2.235008e-07, 2.223851e-07, 2.252924e-07, 2.245972e-07, 2.25459e-07, 
    2.250193e-07, 2.257725e-07, 2.250947e-07, 2.262688e-07, 2.265243e-07, 
    2.263497e-07, 2.270204e-07, 2.250571e-07, 2.258113e-07, 2.201295e-07, 
    2.201629e-07, 2.203189e-07, 2.196332e-07, 2.195912e-07, 2.189626e-07, 
    2.19522e-07, 2.197601e-07, 2.203646e-07, 2.207219e-07, 2.210616e-07, 
    2.218082e-07, 2.226415e-07, 2.238061e-07, 2.246423e-07, 2.252025e-07, 
    2.248591e-07, 2.251623e-07, 2.248233e-07, 2.246644e-07, 2.264285e-07, 
    2.254382e-07, 2.269239e-07, 2.268418e-07, 2.261695e-07, 2.26851e-07, 
    2.201865e-07, 2.199938e-07, 2.193247e-07, 2.198484e-07, 2.188942e-07, 
    2.194283e-07, 2.197353e-07, 2.209196e-07, 2.211798e-07, 2.214209e-07, 
    2.218971e-07, 2.225079e-07, 2.235788e-07, 2.245101e-07, 2.253598e-07, 
    2.252976e-07, 2.253195e-07, 2.255092e-07, 2.250391e-07, 2.255863e-07, 
    2.256781e-07, 2.254381e-07, 2.268308e-07, 2.26433e-07, 2.2684e-07, 
    2.265811e-07, 2.200564e-07, 2.203806e-07, 2.202054e-07, 2.205348e-07, 
    2.203027e-07, 2.213341e-07, 2.216432e-07, 2.230889e-07, 2.224958e-07, 
    2.234397e-07, 2.225918e-07, 2.22742e-07, 2.234703e-07, 2.226376e-07, 
    2.244587e-07, 2.232242e-07, 2.255165e-07, 2.242844e-07, 2.255937e-07, 
    2.253561e-07, 2.257495e-07, 2.261017e-07, 2.265448e-07, 2.273619e-07, 
    2.271727e-07, 2.278558e-07, 2.208637e-07, 2.212839e-07, 2.21247e-07, 
    2.216866e-07, 2.220117e-07, 2.227161e-07, 2.238451e-07, 2.234207e-07, 
    2.241999e-07, 2.243562e-07, 2.231724e-07, 2.238993e-07, 2.215651e-07, 
    2.219424e-07, 2.217178e-07, 2.208968e-07, 2.235184e-07, 2.221735e-07, 
    2.246561e-07, 2.239282e-07, 2.260515e-07, 2.249959e-07, 2.270686e-07, 
    2.279536e-07, 2.287863e-07, 2.297585e-07, 2.215132e-07, 2.212278e-07, 
    2.217389e-07, 2.224457e-07, 2.231014e-07, 2.239726e-07, 2.240618e-07, 
    2.242249e-07, 2.246474e-07, 2.250026e-07, 2.242764e-07, 2.250916e-07, 
    2.220297e-07, 2.236351e-07, 2.211198e-07, 2.218775e-07, 2.224041e-07, 
    2.221732e-07, 2.233722e-07, 2.236546e-07, 2.248017e-07, 2.242089e-07, 
    2.277351e-07, 2.26176e-07, 2.304985e-07, 2.292918e-07, 2.21128e-07, 
    2.215123e-07, 2.228488e-07, 2.222131e-07, 2.240308e-07, 2.244778e-07, 
    2.248413e-07, 2.253055e-07, 2.253557e-07, 2.256307e-07, 2.2518e-07, 
    2.25613e-07, 2.239745e-07, 2.247069e-07, 2.226962e-07, 2.231858e-07, 
    2.229606e-07, 2.227135e-07, 2.23476e-07, 2.242878e-07, 2.243053e-07, 
    2.245654e-07, 2.252982e-07, 2.240381e-07, 2.27936e-07, 2.255298e-07, 
    2.219312e-07, 2.226707e-07, 2.227765e-07, 2.2249e-07, 2.24433e-07, 
    2.237293e-07, 2.25624e-07, 2.251122e-07, 2.259508e-07, 2.255341e-07, 
    2.254728e-07, 2.249375e-07, 2.246041e-07, 2.237615e-07, 2.230756e-07, 
    2.225316e-07, 2.226581e-07, 2.232557e-07, 2.243375e-07, 2.253602e-07, 
    2.251362e-07, 2.258871e-07, 2.238991e-07, 2.247329e-07, 2.244107e-07, 
    2.252508e-07, 2.234094e-07, 2.249773e-07, 2.230083e-07, 2.23181e-07, 
    2.237153e-07, 2.247894e-07, 2.250271e-07, 2.252806e-07, 2.251242e-07, 
    2.243649e-07, 2.242406e-07, 2.237024e-07, 2.235537e-07, 2.231434e-07, 
    2.228037e-07, 2.231141e-07, 2.2344e-07, 2.243653e-07, 2.251987e-07, 
    2.261067e-07, 2.263289e-07, 2.273888e-07, 2.265259e-07, 2.279494e-07, 
    2.26739e-07, 2.288337e-07, 2.250683e-07, 2.267036e-07, 2.237397e-07, 
    2.240593e-07, 2.246371e-07, 2.259618e-07, 2.252469e-07, 2.26083e-07, 
    2.242357e-07, 2.232763e-07, 2.230281e-07, 2.225647e-07, 2.230387e-07, 
    2.230001e-07, 2.234536e-07, 2.233079e-07, 2.24396e-07, 2.238116e-07, 
    2.254713e-07, 2.260764e-07, 2.277842e-07, 2.2883e-07, 2.298941e-07, 
    2.303635e-07, 2.305064e-07, 2.305661e-07,
  2.100066e-07, 2.11004e-07, 2.108101e-07, 2.116145e-07, 2.111684e-07, 
    2.11695e-07, 2.102088e-07, 2.110436e-07, 2.105107e-07, 2.100964e-07, 
    2.131753e-07, 2.116504e-07, 2.147591e-07, 2.137868e-07, 2.162291e-07, 
    2.146078e-07, 2.16556e-07, 2.161824e-07, 2.173068e-07, 2.169847e-07, 
    2.184227e-07, 2.174555e-07, 2.191681e-07, 2.181918e-07, 2.183445e-07, 
    2.174236e-07, 2.119574e-07, 2.129855e-07, 2.118964e-07, 2.120431e-07, 
    2.119773e-07, 2.111776e-07, 2.107745e-07, 2.099304e-07, 2.100836e-07, 
    2.107036e-07, 2.12109e-07, 2.11632e-07, 2.128342e-07, 2.12807e-07, 
    2.141452e-07, 2.135419e-07, 2.157906e-07, 2.151516e-07, 2.169982e-07, 
    2.165338e-07, 2.169764e-07, 2.168422e-07, 2.169781e-07, 2.162971e-07, 
    2.165889e-07, 2.159896e-07, 2.136548e-07, 2.143411e-07, 2.122942e-07, 
    2.110632e-07, 2.102454e-07, 2.096651e-07, 2.097472e-07, 2.099036e-07, 
    2.107072e-07, 2.114628e-07, 2.120386e-07, 2.124237e-07, 2.128031e-07, 
    2.139514e-07, 2.145592e-07, 2.159198e-07, 2.156744e-07, 2.160903e-07, 
    2.164876e-07, 2.171546e-07, 2.170449e-07, 2.173387e-07, 2.160793e-07, 
    2.169163e-07, 2.155345e-07, 2.159125e-07, 2.129061e-07, 2.117607e-07, 
    2.112736e-07, 2.108474e-07, 2.098102e-07, 2.105265e-07, 2.102441e-07, 
    2.109159e-07, 2.113427e-07, 2.111316e-07, 2.124342e-07, 2.119278e-07, 
    2.145952e-07, 2.134464e-07, 2.164413e-07, 2.157248e-07, 2.16613e-07, 
    2.161598e-07, 2.169363e-07, 2.162375e-07, 2.174481e-07, 2.177117e-07, 
    2.175316e-07, 2.182235e-07, 2.161987e-07, 2.169763e-07, 2.111257e-07, 
    2.111601e-07, 2.113205e-07, 2.106154e-07, 2.105723e-07, 2.099262e-07, 
    2.105011e-07, 2.107459e-07, 2.113674e-07, 2.11735e-07, 2.120844e-07, 
    2.128525e-07, 2.137103e-07, 2.149096e-07, 2.157712e-07, 2.163486e-07, 
    2.159946e-07, 2.163072e-07, 2.159577e-07, 2.157939e-07, 2.176129e-07, 
    2.165916e-07, 2.18124e-07, 2.180392e-07, 2.173457e-07, 2.180487e-07, 
    2.111843e-07, 2.109862e-07, 2.102983e-07, 2.108366e-07, 2.098558e-07, 
    2.104048e-07, 2.107205e-07, 2.119384e-07, 2.12206e-07, 2.12454e-07, 
    2.12944e-07, 2.135727e-07, 2.146756e-07, 2.15635e-07, 2.165107e-07, 
    2.164466e-07, 2.164692e-07, 2.166648e-07, 2.161802e-07, 2.167443e-07, 
    2.16839e-07, 2.165915e-07, 2.180278e-07, 2.176175e-07, 2.180374e-07, 
    2.177702e-07, 2.110506e-07, 2.113839e-07, 2.112038e-07, 2.115425e-07, 
    2.113039e-07, 2.123648e-07, 2.126829e-07, 2.14171e-07, 2.135604e-07, 
    2.145323e-07, 2.136591e-07, 2.138138e-07, 2.145639e-07, 2.137063e-07, 
    2.155821e-07, 2.143104e-07, 2.166724e-07, 2.154026e-07, 2.167519e-07, 
    2.16507e-07, 2.169126e-07, 2.172758e-07, 2.177328e-07, 2.185759e-07, 
    2.183807e-07, 2.190857e-07, 2.118808e-07, 2.123131e-07, 2.122751e-07, 
    2.127274e-07, 2.13062e-07, 2.137871e-07, 2.149498e-07, 2.145126e-07, 
    2.153153e-07, 2.154764e-07, 2.14257e-07, 2.150057e-07, 2.126024e-07, 
    2.129907e-07, 2.127595e-07, 2.119149e-07, 2.146133e-07, 2.132286e-07, 
    2.157854e-07, 2.150354e-07, 2.17224e-07, 2.161357e-07, 2.182732e-07, 
    2.191867e-07, 2.200465e-07, 2.210509e-07, 2.12549e-07, 2.122553e-07, 
    2.127813e-07, 2.135088e-07, 2.141839e-07, 2.150812e-07, 2.15173e-07, 
    2.153411e-07, 2.157765e-07, 2.161425e-07, 2.153942e-07, 2.162343e-07, 
    2.130807e-07, 2.147335e-07, 2.121443e-07, 2.12924e-07, 2.134659e-07, 
    2.132282e-07, 2.144626e-07, 2.147536e-07, 2.159355e-07, 2.153246e-07, 
    2.189613e-07, 2.173525e-07, 2.218157e-07, 2.205688e-07, 2.121527e-07, 
    2.12548e-07, 2.139238e-07, 2.132693e-07, 2.151411e-07, 2.156017e-07, 
    2.159762e-07, 2.164549e-07, 2.165065e-07, 2.167901e-07, 2.163254e-07, 
    2.167718e-07, 2.150831e-07, 2.158378e-07, 2.137666e-07, 2.142708e-07, 
    2.140388e-07, 2.137844e-07, 2.145696e-07, 2.15406e-07, 2.154239e-07, 
    2.15692e-07, 2.164475e-07, 2.151487e-07, 2.191688e-07, 2.166863e-07, 
    2.129791e-07, 2.137405e-07, 2.138493e-07, 2.135544e-07, 2.155556e-07, 
    2.148305e-07, 2.167832e-07, 2.162555e-07, 2.171201e-07, 2.166905e-07, 
    2.166273e-07, 2.160755e-07, 2.157319e-07, 2.148638e-07, 2.141573e-07, 
    2.135971e-07, 2.137274e-07, 2.143428e-07, 2.154571e-07, 2.165112e-07, 
    2.162803e-07, 2.170544e-07, 2.150054e-07, 2.158646e-07, 2.155325e-07, 
    2.163985e-07, 2.14501e-07, 2.161167e-07, 2.140879e-07, 2.142658e-07, 
    2.148161e-07, 2.159229e-07, 2.161678e-07, 2.164292e-07, 2.162679e-07, 
    2.154854e-07, 2.153572e-07, 2.148028e-07, 2.146496e-07, 2.142271e-07, 
    2.138773e-07, 2.141969e-07, 2.145325e-07, 2.154858e-07, 2.163447e-07, 
    2.17281e-07, 2.175101e-07, 2.186038e-07, 2.177135e-07, 2.191826e-07, 
    2.179335e-07, 2.200957e-07, 2.162104e-07, 2.178968e-07, 2.148412e-07, 
    2.151704e-07, 2.157659e-07, 2.171316e-07, 2.163944e-07, 2.172565e-07, 
    2.153522e-07, 2.14364e-07, 2.141083e-07, 2.136312e-07, 2.141192e-07, 
    2.140795e-07, 2.145465e-07, 2.143964e-07, 2.155174e-07, 2.149153e-07, 
    2.166257e-07, 2.172497e-07, 2.190118e-07, 2.200918e-07, 2.211909e-07, 
    2.216761e-07, 2.218238e-07, 2.218855e-07,
  2.030027e-07, 2.039495e-07, 2.037654e-07, 2.045295e-07, 2.041056e-07, 
    2.04606e-07, 2.031946e-07, 2.039871e-07, 2.034812e-07, 2.030879e-07, 
    2.060135e-07, 2.045636e-07, 2.075213e-07, 2.065953e-07, 2.089227e-07, 
    2.073772e-07, 2.092346e-07, 2.088781e-07, 2.099513e-07, 2.096438e-07, 
    2.110176e-07, 2.100933e-07, 2.117303e-07, 2.107968e-07, 2.109428e-07, 
    2.100628e-07, 2.048552e-07, 2.058329e-07, 2.047973e-07, 2.049367e-07, 
    2.048741e-07, 2.041143e-07, 2.037316e-07, 2.029304e-07, 2.030758e-07, 
    2.036643e-07, 2.049994e-07, 2.04546e-07, 2.056888e-07, 2.05663e-07, 
    2.069365e-07, 2.063622e-07, 2.085045e-07, 2.078952e-07, 2.096566e-07, 
    2.092134e-07, 2.096358e-07, 2.095077e-07, 2.096375e-07, 2.089875e-07, 
    2.092659e-07, 2.086942e-07, 2.064697e-07, 2.071231e-07, 2.051754e-07, 
    2.040058e-07, 2.032294e-07, 2.026787e-07, 2.027566e-07, 2.02905e-07, 
    2.036677e-07, 2.043853e-07, 2.049324e-07, 2.052985e-07, 2.056593e-07, 
    2.067521e-07, 2.073309e-07, 2.086277e-07, 2.083936e-07, 2.087903e-07, 
    2.091693e-07, 2.09806e-07, 2.097012e-07, 2.099818e-07, 2.087798e-07, 
    2.095785e-07, 2.082602e-07, 2.086206e-07, 2.057575e-07, 2.046683e-07, 
    2.042057e-07, 2.038008e-07, 2.028164e-07, 2.034961e-07, 2.032281e-07, 
    2.038658e-07, 2.042711e-07, 2.040706e-07, 2.053085e-07, 2.048271e-07, 
    2.073652e-07, 2.062714e-07, 2.091251e-07, 2.084416e-07, 2.09289e-07, 
    2.088565e-07, 2.095976e-07, 2.089306e-07, 2.100862e-07, 2.10338e-07, 
    2.10166e-07, 2.10827e-07, 2.088937e-07, 2.096358e-07, 2.04065e-07, 
    2.040977e-07, 2.042501e-07, 2.035806e-07, 2.035396e-07, 2.029264e-07, 
    2.03472e-07, 2.037044e-07, 2.042946e-07, 2.046439e-07, 2.049759e-07, 
    2.057063e-07, 2.065225e-07, 2.076647e-07, 2.084859e-07, 2.090367e-07, 
    2.086989e-07, 2.089971e-07, 2.086638e-07, 2.085076e-07, 2.102437e-07, 
    2.092685e-07, 2.107319e-07, 2.106509e-07, 2.099885e-07, 2.1066e-07, 
    2.041207e-07, 2.039325e-07, 2.032795e-07, 2.037905e-07, 2.028596e-07, 
    2.033806e-07, 2.036803e-07, 2.048372e-07, 2.050915e-07, 2.053274e-07, 
    2.057933e-07, 2.063915e-07, 2.074417e-07, 2.083561e-07, 2.091914e-07, 
    2.091301e-07, 2.091517e-07, 2.093384e-07, 2.08876e-07, 2.094143e-07, 
    2.095047e-07, 2.092684e-07, 2.106401e-07, 2.10248e-07, 2.106492e-07, 
    2.103939e-07, 2.039937e-07, 2.043103e-07, 2.041392e-07, 2.04461e-07, 
    2.042343e-07, 2.052426e-07, 2.05545e-07, 2.069612e-07, 2.063798e-07, 
    2.073052e-07, 2.064737e-07, 2.06621e-07, 2.073354e-07, 2.065186e-07, 
    2.083057e-07, 2.070939e-07, 2.093456e-07, 2.081346e-07, 2.094216e-07, 
    2.091878e-07, 2.095749e-07, 2.099217e-07, 2.103582e-07, 2.11164e-07, 
    2.109773e-07, 2.116515e-07, 2.047824e-07, 2.051934e-07, 2.051572e-07, 
    2.055873e-07, 2.059056e-07, 2.065955e-07, 2.07703e-07, 2.072864e-07, 
    2.080512e-07, 2.082049e-07, 2.070429e-07, 2.077562e-07, 2.054685e-07, 
    2.058378e-07, 2.056179e-07, 2.048149e-07, 2.073824e-07, 2.060641e-07, 
    2.084995e-07, 2.077845e-07, 2.098723e-07, 2.088336e-07, 2.108746e-07, 
    2.117482e-07, 2.125709e-07, 2.135331e-07, 2.054177e-07, 2.051384e-07, 
    2.056385e-07, 2.063308e-07, 2.069733e-07, 2.078281e-07, 2.079156e-07, 
    2.080758e-07, 2.084909e-07, 2.0884e-07, 2.081265e-07, 2.089276e-07, 
    2.059235e-07, 2.074969e-07, 2.050328e-07, 2.057744e-07, 2.062899e-07, 
    2.060637e-07, 2.072388e-07, 2.075159e-07, 2.086427e-07, 2.080601e-07, 
    2.115325e-07, 2.09995e-07, 2.142662e-07, 2.130711e-07, 2.050408e-07, 
    2.054167e-07, 2.067258e-07, 2.061028e-07, 2.078852e-07, 2.083244e-07, 
    2.086814e-07, 2.091381e-07, 2.091874e-07, 2.09458e-07, 2.090146e-07, 
    2.094405e-07, 2.0783e-07, 2.085494e-07, 2.06576e-07, 2.070561e-07, 
    2.068352e-07, 2.06593e-07, 2.073407e-07, 2.081378e-07, 2.081548e-07, 
    2.084105e-07, 2.091313e-07, 2.078925e-07, 2.117312e-07, 2.093591e-07, 
    2.058267e-07, 2.065513e-07, 2.066548e-07, 2.06374e-07, 2.082803e-07, 
    2.075893e-07, 2.094514e-07, 2.089479e-07, 2.09773e-07, 2.093629e-07, 
    2.093026e-07, 2.087761e-07, 2.084484e-07, 2.07621e-07, 2.069481e-07, 
    2.064147e-07, 2.065387e-07, 2.071247e-07, 2.081865e-07, 2.091919e-07, 
    2.089716e-07, 2.097103e-07, 2.077559e-07, 2.085751e-07, 2.082584e-07, 
    2.090842e-07, 2.072754e-07, 2.088156e-07, 2.068819e-07, 2.070514e-07, 
    2.075756e-07, 2.086307e-07, 2.088642e-07, 2.091136e-07, 2.089597e-07, 
    2.082135e-07, 2.080913e-07, 2.075628e-07, 2.07417e-07, 2.070145e-07, 
    2.066814e-07, 2.069857e-07, 2.073054e-07, 2.082138e-07, 2.09033e-07, 
    2.099267e-07, 2.101455e-07, 2.111908e-07, 2.103398e-07, 2.117444e-07, 
    2.105502e-07, 2.126181e-07, 2.089049e-07, 2.10515e-07, 2.075994e-07, 
    2.079132e-07, 2.08481e-07, 2.097841e-07, 2.090804e-07, 2.099034e-07, 
    2.080865e-07, 2.071449e-07, 2.069014e-07, 2.064472e-07, 2.069117e-07, 
    2.068739e-07, 2.073186e-07, 2.071757e-07, 2.08244e-07, 2.0767e-07, 
    2.093011e-07, 2.098969e-07, 2.115808e-07, 2.126143e-07, 2.136671e-07, 
    2.141323e-07, 2.142739e-07, 2.143331e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.652399e-13, 9.678468e-13, 9.673404e-13, 9.69441e-13, 9.682762e-13, 
    9.696512e-13, 9.65769e-13, 9.679499e-13, 9.665581e-13, 9.654752e-13, 
    9.735113e-13, 9.695348e-13, 9.776379e-13, 9.751066e-13, 9.814612e-13, 
    9.772438e-13, 9.823108e-13, 9.813404e-13, 9.842616e-13, 9.834251e-13, 
    9.871558e-13, 9.846476e-13, 9.890884e-13, 9.865574e-13, 9.869532e-13, 
    9.845646e-13, 9.703362e-13, 9.730164e-13, 9.701772e-13, 9.705597e-13, 
    9.703883e-13, 9.683001e-13, 9.672466e-13, 9.650411e-13, 9.654418e-13, 
    9.670618e-13, 9.707316e-13, 9.69487e-13, 9.726239e-13, 9.725531e-13, 
    9.760401e-13, 9.744686e-13, 9.803222e-13, 9.786601e-13, 9.834602e-13, 
    9.822538e-13, 9.834034e-13, 9.830549e-13, 9.834079e-13, 9.816385e-13, 
    9.823967e-13, 9.808393e-13, 9.747628e-13, 9.765501e-13, 9.712151e-13, 
    9.680003e-13, 9.658645e-13, 9.643473e-13, 9.645619e-13, 9.649706e-13, 
    9.670714e-13, 9.690454e-13, 9.705484e-13, 9.715532e-13, 9.725429e-13, 
    9.755342e-13, 9.771176e-13, 9.806576e-13, 9.800199e-13, 9.811007e-13, 
    9.821338e-13, 9.838663e-13, 9.835813e-13, 9.843441e-13, 9.810728e-13, 
    9.832472e-13, 9.796564e-13, 9.80639e-13, 9.728094e-13, 9.69823e-13, 
    9.685502e-13, 9.674376e-13, 9.647268e-13, 9.66599e-13, 9.658611e-13, 
    9.676169e-13, 9.687315e-13, 9.681804e-13, 9.715807e-13, 9.702592e-13, 
    9.772114e-13, 9.742194e-13, 9.820133e-13, 9.801509e-13, 9.824597e-13, 
    9.812819e-13, 9.832993e-13, 9.814838e-13, 9.846282e-13, 9.85312e-13, 
    9.848446e-13, 9.866401e-13, 9.813831e-13, 9.83403e-13, 9.681649e-13, 
    9.682548e-13, 9.686737e-13, 9.668314e-13, 9.667188e-13, 9.650299e-13, 
    9.66533e-13, 9.671725e-13, 9.687963e-13, 9.697559e-13, 9.706678e-13, 
    9.726715e-13, 9.74907e-13, 9.7803e-13, 9.802715e-13, 9.817727e-13, 
    9.808526e-13, 9.816649e-13, 9.807566e-13, 9.803309e-13, 9.850556e-13, 
    9.824036e-13, 9.86382e-13, 9.861621e-13, 9.843621e-13, 9.861868e-13, 
    9.683179e-13, 9.678006e-13, 9.660028e-13, 9.674099e-13, 9.64846e-13, 
    9.662811e-13, 9.671057e-13, 9.702864e-13, 9.709851e-13, 9.716322e-13, 
    9.729102e-13, 9.74549e-13, 9.774209e-13, 9.799172e-13, 9.82194e-13, 
    9.820273e-13, 9.820859e-13, 9.82594e-13, 9.813349e-13, 9.828006e-13, 
    9.830463e-13, 9.824036e-13, 9.861326e-13, 9.850679e-13, 9.861574e-13, 
    9.854643e-13, 9.679688e-13, 9.688393e-13, 9.683689e-13, 9.692532e-13, 
    9.6863e-13, 9.71399e-13, 9.722285e-13, 9.761069e-13, 9.745166e-13, 
    9.770478e-13, 9.747741e-13, 9.75177e-13, 9.771292e-13, 9.748971e-13, 
    9.797791e-13, 9.764694e-13, 9.826137e-13, 9.793118e-13, 9.828205e-13, 
    9.821842e-13, 9.832379e-13, 9.841808e-13, 9.853672e-13, 9.875536e-13, 
    9.870476e-13, 9.888752e-13, 9.701366e-13, 9.712643e-13, 9.711655e-13, 
    9.723455e-13, 9.732176e-13, 9.751076e-13, 9.781349e-13, 9.769971e-13, 
    9.790861e-13, 9.79505e-13, 9.763315e-13, 9.782801e-13, 9.720191e-13, 
    9.730312e-13, 9.724291e-13, 9.702253e-13, 9.772586e-13, 9.736515e-13, 
    9.803085e-13, 9.783578e-13, 9.840464e-13, 9.812186e-13, 9.867688e-13, 
    9.891361e-13, 9.913638e-13, 9.939616e-13, 9.7188e-13, 9.71114e-13, 
    9.724859e-13, 9.743818e-13, 9.761409e-13, 9.784767e-13, 9.787158e-13, 
    9.79153e-13, 9.802855e-13, 9.81237e-13, 9.792907e-13, 9.814755e-13, 
    9.73265e-13, 9.775718e-13, 9.708239e-13, 9.728572e-13, 9.742703e-13, 
    9.73651e-13, 9.768671e-13, 9.776243e-13, 9.806985e-13, 9.791101e-13, 
    9.885516e-13, 9.843794e-13, 9.959391e-13, 9.927146e-13, 9.708461e-13, 
    9.718776e-13, 9.754633e-13, 9.73758e-13, 9.786328e-13, 9.798309e-13, 
    9.808048e-13, 9.820484e-13, 9.821831e-13, 9.829196e-13, 9.817124e-13, 
    9.828721e-13, 9.784816e-13, 9.804448e-13, 9.750543e-13, 9.763672e-13, 
    9.757635e-13, 9.751008e-13, 9.771456e-13, 9.793212e-13, 9.793685e-13, 
    9.800655e-13, 9.820272e-13, 9.786526e-13, 9.89088e-13, 9.826478e-13, 
    9.730018e-13, 9.749854e-13, 9.752695e-13, 9.745013e-13, 9.797108e-13, 
    9.778245e-13, 9.829017e-13, 9.815308e-13, 9.837768e-13, 9.826609e-13, 
    9.824966e-13, 9.810628e-13, 9.801694e-13, 9.779108e-13, 9.760718e-13, 
    9.746128e-13, 9.749522e-13, 9.765546e-13, 9.794544e-13, 9.821949e-13, 
    9.815947e-13, 9.836062e-13, 9.782796e-13, 9.805143e-13, 9.796506e-13, 
    9.819021e-13, 9.769667e-13, 9.811677e-13, 9.758914e-13, 9.763546e-13, 
    9.77787e-13, 9.806652e-13, 9.813027e-13, 9.819817e-13, 9.815629e-13, 
    9.795281e-13, 9.791949e-13, 9.777524e-13, 9.773535e-13, 9.762538e-13, 
    9.753425e-13, 9.76175e-13, 9.770486e-13, 9.795293e-13, 9.817621e-13, 
    9.841942e-13, 9.847893e-13, 9.876248e-13, 9.853158e-13, 9.891237e-13, 
    9.85885e-13, 9.914891e-13, 9.814121e-13, 9.857913e-13, 9.778525e-13, 
    9.787092e-13, 9.802573e-13, 9.838056e-13, 9.818915e-13, 9.841302e-13, 
    9.791819e-13, 9.766094e-13, 9.759444e-13, 9.747013e-13, 9.759728e-13, 
    9.758695e-13, 9.770854e-13, 9.766947e-13, 9.796117e-13, 9.780453e-13, 
    9.824923e-13, 9.841127e-13, 9.886835e-13, 9.914802e-13, 9.943246e-13, 
    9.955787e-13, 9.959604e-13, 9.961199e-13 ;

 LITR1C =
  3.066846e-05, 3.066834e-05, 3.066836e-05, 3.066827e-05, 3.066832e-05, 
    3.066826e-05, 3.066843e-05, 3.066833e-05, 3.06684e-05, 3.066845e-05, 
    3.066808e-05, 3.066826e-05, 3.06679e-05, 3.066801e-05, 3.066772e-05, 
    3.066791e-05, 3.066768e-05, 3.066773e-05, 3.066759e-05, 3.066763e-05, 
    3.066746e-05, 3.066758e-05, 3.066738e-05, 3.066749e-05, 3.066747e-05, 
    3.066758e-05, 3.066823e-05, 3.06681e-05, 3.066823e-05, 3.066822e-05, 
    3.066822e-05, 3.066832e-05, 3.066837e-05, 3.066846e-05, 3.066845e-05, 
    3.066837e-05, 3.066821e-05, 3.066826e-05, 3.066812e-05, 3.066812e-05, 
    3.066797e-05, 3.066804e-05, 3.066777e-05, 3.066785e-05, 3.066763e-05, 
    3.066768e-05, 3.066763e-05, 3.066765e-05, 3.066763e-05, 3.066771e-05, 
    3.066768e-05, 3.066775e-05, 3.066802e-05, 3.066794e-05, 3.066819e-05, 
    3.066833e-05, 3.066843e-05, 3.06685e-05, 3.066849e-05, 3.066847e-05, 
    3.066837e-05, 3.066829e-05, 3.066822e-05, 3.066817e-05, 3.066812e-05, 
    3.066799e-05, 3.066792e-05, 3.066776e-05, 3.066779e-05, 3.066774e-05, 
    3.066769e-05, 3.066761e-05, 3.066763e-05, 3.066759e-05, 3.066774e-05, 
    3.066764e-05, 3.06678e-05, 3.066776e-05, 3.066811e-05, 3.066825e-05, 
    3.066831e-05, 3.066836e-05, 3.066848e-05, 3.066839e-05, 3.066843e-05, 
    3.066835e-05, 3.06683e-05, 3.066832e-05, 3.066817e-05, 3.066823e-05, 
    3.066791e-05, 3.066805e-05, 3.06677e-05, 3.066778e-05, 3.066768e-05, 
    3.066773e-05, 3.066764e-05, 3.066772e-05, 3.066758e-05, 3.066755e-05, 
    3.066757e-05, 3.066749e-05, 3.066772e-05, 3.066763e-05, 3.066833e-05, 
    3.066832e-05, 3.06683e-05, 3.066838e-05, 3.066839e-05, 3.066847e-05, 
    3.06684e-05, 3.066837e-05, 3.06683e-05, 3.066825e-05, 3.066821e-05, 
    3.066812e-05, 3.066802e-05, 3.066788e-05, 3.066778e-05, 3.066771e-05, 
    3.066775e-05, 3.066771e-05, 3.066775e-05, 3.066777e-05, 3.066756e-05, 
    3.066768e-05, 3.06675e-05, 3.066751e-05, 3.066759e-05, 3.066751e-05, 
    3.066832e-05, 3.066834e-05, 3.066842e-05, 3.066836e-05, 3.066847e-05, 
    3.066841e-05, 3.066837e-05, 3.066823e-05, 3.066819e-05, 3.066816e-05, 
    3.066811e-05, 3.066803e-05, 3.06679e-05, 3.066779e-05, 3.066769e-05, 
    3.06677e-05, 3.066769e-05, 3.066767e-05, 3.066773e-05, 3.066766e-05, 
    3.066765e-05, 3.066768e-05, 3.066751e-05, 3.066756e-05, 3.066751e-05, 
    3.066754e-05, 3.066833e-05, 3.066829e-05, 3.066831e-05, 3.066827e-05, 
    3.06683e-05, 3.066818e-05, 3.066814e-05, 3.066796e-05, 3.066804e-05, 
    3.066792e-05, 3.066802e-05, 3.0668e-05, 3.066792e-05, 3.066802e-05, 
    3.06678e-05, 3.066795e-05, 3.066767e-05, 3.066782e-05, 3.066766e-05, 
    3.066769e-05, 3.066764e-05, 3.06676e-05, 3.066755e-05, 3.066744e-05, 
    3.066747e-05, 3.066739e-05, 3.066823e-05, 3.066818e-05, 3.066819e-05, 
    3.066814e-05, 3.06681e-05, 3.066801e-05, 3.066787e-05, 3.066792e-05, 
    3.066783e-05, 3.066781e-05, 3.066795e-05, 3.066787e-05, 3.066815e-05, 
    3.06681e-05, 3.066813e-05, 3.066823e-05, 3.066791e-05, 3.066807e-05, 
    3.066777e-05, 3.066786e-05, 3.06676e-05, 3.066773e-05, 3.066748e-05, 
    3.066738e-05, 3.066727e-05, 3.066716e-05, 3.066815e-05, 3.066819e-05, 
    3.066813e-05, 3.066804e-05, 3.066796e-05, 3.066786e-05, 3.066784e-05, 
    3.066783e-05, 3.066778e-05, 3.066773e-05, 3.066782e-05, 3.066772e-05, 
    3.066809e-05, 3.06679e-05, 3.06682e-05, 3.066811e-05, 3.066805e-05, 
    3.066807e-05, 3.066793e-05, 3.06679e-05, 3.066776e-05, 3.066783e-05, 
    3.06674e-05, 3.066759e-05, 3.066707e-05, 3.066721e-05, 3.06682e-05, 
    3.066815e-05, 3.066799e-05, 3.066807e-05, 3.066785e-05, 3.066779e-05, 
    3.066775e-05, 3.06677e-05, 3.066769e-05, 3.066766e-05, 3.066771e-05, 
    3.066766e-05, 3.066786e-05, 3.066777e-05, 3.066801e-05, 3.066795e-05, 
    3.066798e-05, 3.066801e-05, 3.066792e-05, 3.066782e-05, 3.066782e-05, 
    3.066779e-05, 3.06677e-05, 3.066785e-05, 3.066738e-05, 3.066767e-05, 
    3.06681e-05, 3.066802e-05, 3.0668e-05, 3.066804e-05, 3.06678e-05, 
    3.066788e-05, 3.066766e-05, 3.066772e-05, 3.066762e-05, 3.066767e-05, 
    3.066767e-05, 3.066774e-05, 3.066778e-05, 3.066788e-05, 3.066796e-05, 
    3.066803e-05, 3.066802e-05, 3.066794e-05, 3.066781e-05, 3.066769e-05, 
    3.066771e-05, 3.066762e-05, 3.066787e-05, 3.066776e-05, 3.06678e-05, 
    3.06677e-05, 3.066792e-05, 3.066774e-05, 3.066797e-05, 3.066795e-05, 
    3.066789e-05, 3.066776e-05, 3.066773e-05, 3.06677e-05, 3.066772e-05, 
    3.066781e-05, 3.066782e-05, 3.066789e-05, 3.066791e-05, 3.066796e-05, 
    3.0668e-05, 3.066796e-05, 3.066792e-05, 3.066781e-05, 3.066771e-05, 
    3.06676e-05, 3.066757e-05, 3.066744e-05, 3.066755e-05, 3.066738e-05, 
    3.066752e-05, 3.066727e-05, 3.066772e-05, 3.066752e-05, 3.066788e-05, 
    3.066784e-05, 3.066778e-05, 3.066762e-05, 3.06677e-05, 3.06676e-05, 
    3.066783e-05, 3.066794e-05, 3.066797e-05, 3.066803e-05, 3.066797e-05, 
    3.066798e-05, 3.066792e-05, 3.066794e-05, 3.06678e-05, 3.066788e-05, 
    3.066767e-05, 3.06676e-05, 3.066739e-05, 3.066727e-05, 3.066714e-05, 
    3.066708e-05, 3.066707e-05, 3.066706e-05 ;

 LITR1C_TO_SOIL1C =
  6.428924e-13, 6.446283e-13, 6.442911e-13, 6.456899e-13, 6.449143e-13, 
    6.458299e-13, 6.432447e-13, 6.44697e-13, 6.437701e-13, 6.43049e-13, 
    6.484004e-13, 6.457524e-13, 6.511484e-13, 6.494627e-13, 6.536944e-13, 
    6.508859e-13, 6.542601e-13, 6.536139e-13, 6.555592e-13, 6.550022e-13, 
    6.574864e-13, 6.558162e-13, 6.587734e-13, 6.57088e-13, 6.573516e-13, 
    6.55761e-13, 6.462861e-13, 6.480708e-13, 6.461802e-13, 6.464348e-13, 
    6.463207e-13, 6.449302e-13, 6.442286e-13, 6.427599e-13, 6.430268e-13, 
    6.441056e-13, 6.465494e-13, 6.457206e-13, 6.478095e-13, 6.477623e-13, 
    6.500844e-13, 6.490378e-13, 6.529358e-13, 6.518291e-13, 6.550255e-13, 
    6.542222e-13, 6.549877e-13, 6.547557e-13, 6.549907e-13, 6.538124e-13, 
    6.543173e-13, 6.532803e-13, 6.492338e-13, 6.50424e-13, 6.468713e-13, 
    6.447306e-13, 6.433083e-13, 6.422979e-13, 6.424408e-13, 6.42713e-13, 
    6.441119e-13, 6.454265e-13, 6.464274e-13, 6.470965e-13, 6.477556e-13, 
    6.497475e-13, 6.508019e-13, 6.531593e-13, 6.527345e-13, 6.534543e-13, 
    6.541423e-13, 6.552959e-13, 6.551062e-13, 6.556141e-13, 6.534356e-13, 
    6.548837e-13, 6.524924e-13, 6.531468e-13, 6.47933e-13, 6.459443e-13, 
    6.450968e-13, 6.443559e-13, 6.425506e-13, 6.437974e-13, 6.43306e-13, 
    6.444752e-13, 6.452175e-13, 6.448505e-13, 6.471148e-13, 6.462348e-13, 
    6.508643e-13, 6.48872e-13, 6.54062e-13, 6.528218e-13, 6.543592e-13, 
    6.53575e-13, 6.549183e-13, 6.537094e-13, 6.558033e-13, 6.562586e-13, 
    6.559474e-13, 6.571431e-13, 6.536423e-13, 6.549875e-13, 6.448401e-13, 
    6.449e-13, 6.45179e-13, 6.439522e-13, 6.438771e-13, 6.427526e-13, 
    6.437534e-13, 6.441793e-13, 6.452606e-13, 6.458996e-13, 6.465068e-13, 
    6.478412e-13, 6.493298e-13, 6.514095e-13, 6.529022e-13, 6.539018e-13, 
    6.532891e-13, 6.538301e-13, 6.532252e-13, 6.529417e-13, 6.560879e-13, 
    6.543219e-13, 6.569712e-13, 6.568247e-13, 6.556262e-13, 6.568412e-13, 
    6.44942e-13, 6.445975e-13, 6.434004e-13, 6.443373e-13, 6.4263e-13, 
    6.435857e-13, 6.441348e-13, 6.462529e-13, 6.467182e-13, 6.471491e-13, 
    6.480001e-13, 6.490914e-13, 6.510039e-13, 6.526662e-13, 6.541823e-13, 
    6.540714e-13, 6.541104e-13, 6.544487e-13, 6.536103e-13, 6.545864e-13, 
    6.5475e-13, 6.543219e-13, 6.568051e-13, 6.560962e-13, 6.568216e-13, 
    6.563601e-13, 6.447095e-13, 6.452892e-13, 6.44976e-13, 6.455649e-13, 
    6.451499e-13, 6.469937e-13, 6.475461e-13, 6.501289e-13, 6.490698e-13, 
    6.507554e-13, 6.492413e-13, 6.495096e-13, 6.508096e-13, 6.493233e-13, 
    6.525742e-13, 6.503703e-13, 6.544619e-13, 6.52263e-13, 6.545995e-13, 
    6.541758e-13, 6.548775e-13, 6.555054e-13, 6.562954e-13, 6.577514e-13, 
    6.574144e-13, 6.586315e-13, 6.461531e-13, 6.469041e-13, 6.468383e-13, 
    6.47624e-13, 6.482049e-13, 6.494634e-13, 6.514794e-13, 6.507217e-13, 
    6.521127e-13, 6.523917e-13, 6.502784e-13, 6.51576e-13, 6.474067e-13, 
    6.480808e-13, 6.476797e-13, 6.462122e-13, 6.508958e-13, 6.484937e-13, 
    6.529268e-13, 6.516277e-13, 6.554159e-13, 6.535328e-13, 6.572288e-13, 
    6.588052e-13, 6.602886e-13, 6.620186e-13, 6.473141e-13, 6.46804e-13, 
    6.477176e-13, 6.489801e-13, 6.501515e-13, 6.517069e-13, 6.518662e-13, 
    6.521573e-13, 6.529114e-13, 6.53545e-13, 6.52249e-13, 6.537039e-13, 
    6.482364e-13, 6.511043e-13, 6.466108e-13, 6.479648e-13, 6.489058e-13, 
    6.484934e-13, 6.506351e-13, 6.511394e-13, 6.531865e-13, 6.521287e-13, 
    6.584159e-13, 6.556376e-13, 6.633354e-13, 6.611882e-13, 6.466257e-13, 
    6.473126e-13, 6.497003e-13, 6.485647e-13, 6.518109e-13, 6.526087e-13, 
    6.532573e-13, 6.540854e-13, 6.541751e-13, 6.546655e-13, 6.538617e-13, 
    6.546339e-13, 6.517102e-13, 6.530175e-13, 6.494279e-13, 6.503022e-13, 
    6.499002e-13, 6.494588e-13, 6.508205e-13, 6.522693e-13, 6.523008e-13, 
    6.52765e-13, 6.540713e-13, 6.51824e-13, 6.587732e-13, 6.544845e-13, 
    6.480611e-13, 6.49382e-13, 6.495712e-13, 6.490596e-13, 6.525288e-13, 
    6.512726e-13, 6.546536e-13, 6.537407e-13, 6.552363e-13, 6.544933e-13, 
    6.543839e-13, 6.53429e-13, 6.528341e-13, 6.513301e-13, 6.501055e-13, 
    6.491339e-13, 6.493599e-13, 6.50427e-13, 6.52358e-13, 6.541829e-13, 
    6.537833e-13, 6.551227e-13, 6.515757e-13, 6.530638e-13, 6.524886e-13, 
    6.539879e-13, 6.507014e-13, 6.53499e-13, 6.499853e-13, 6.502938e-13, 
    6.512477e-13, 6.531643e-13, 6.535888e-13, 6.54041e-13, 6.537621e-13, 
    6.524071e-13, 6.521852e-13, 6.512246e-13, 6.50959e-13, 6.502267e-13, 
    6.496199e-13, 6.501742e-13, 6.50756e-13, 6.524079e-13, 6.538947e-13, 
    6.555143e-13, 6.559105e-13, 6.577988e-13, 6.562612e-13, 6.587969e-13, 
    6.566403e-13, 6.603721e-13, 6.536617e-13, 6.565778e-13, 6.512912e-13, 
    6.518618e-13, 6.528927e-13, 6.552555e-13, 6.539809e-13, 6.554717e-13, 
    6.521766e-13, 6.504635e-13, 6.500206e-13, 6.491929e-13, 6.500395e-13, 
    6.499707e-13, 6.507804e-13, 6.505203e-13, 6.524627e-13, 6.514197e-13, 
    6.54381e-13, 6.554601e-13, 6.585038e-13, 6.603661e-13, 6.622603e-13, 
    6.630954e-13, 6.633495e-13, 6.634557e-13 ;

 LITR1C_vr =
  0.001751201, 0.001751194, 0.001751195, 0.00175119, 0.001751193, 
    0.001751189, 0.001751199, 0.001751194, 0.001751197, 0.0017512, 
    0.001751179, 0.001751189, 0.001751169, 0.001751175, 0.001751159, 
    0.001751169, 0.001751156, 0.001751159, 0.001751151, 0.001751153, 
    0.001751144, 0.00175115, 0.001751139, 0.001751145, 0.001751144, 
    0.001751151, 0.001751187, 0.00175118, 0.001751188, 0.001751187, 
    0.001751187, 0.001751193, 0.001751195, 0.001751201, 0.0017512, 
    0.001751196, 0.001751186, 0.00175119, 0.001751181, 0.001751182, 
    0.001751173, 0.001751177, 0.001751162, 0.001751166, 0.001751153, 
    0.001751157, 0.001751154, 0.001751154, 0.001751154, 0.001751158, 
    0.001751156, 0.00175116, 0.001751176, 0.001751171, 0.001751185, 
    0.001751193, 0.001751199, 0.001751203, 0.001751202, 0.001751201, 
    0.001751196, 0.001751191, 0.001751187, 0.001751184, 0.001751182, 
    0.001751174, 0.00175117, 0.001751161, 0.001751162, 0.00175116, 
    0.001751157, 0.001751152, 0.001751153, 0.001751151, 0.00175116, 
    0.001751154, 0.001751163, 0.001751161, 0.001751181, 0.001751189, 
    0.001751192, 0.001751195, 0.001751202, 0.001751197, 0.001751199, 
    0.001751194, 0.001751191, 0.001751193, 0.001751184, 0.001751188, 
    0.00175117, 0.001751177, 0.001751157, 0.001751162, 0.001751156, 
    0.001751159, 0.001751154, 0.001751159, 0.00175115, 0.001751149, 
    0.00175115, 0.001751145, 0.001751159, 0.001751154, 0.001751193, 
    0.001751193, 0.001751192, 0.001751196, 0.001751197, 0.001751201, 
    0.001751197, 0.001751196, 0.001751191, 0.001751189, 0.001751186, 
    0.001751181, 0.001751175, 0.001751167, 0.001751162, 0.001751158, 
    0.00175116, 0.001751158, 0.00175116, 0.001751162, 0.001751149, 
    0.001751156, 0.001751146, 0.001751146, 0.001751151, 0.001751146, 
    0.001751193, 0.001751194, 0.001751199, 0.001751195, 0.001751202, 
    0.001751198, 0.001751196, 0.001751187, 0.001751186, 0.001751184, 
    0.001751181, 0.001751176, 0.001751169, 0.001751163, 0.001751157, 
    0.001751157, 0.001751157, 0.001751156, 0.001751159, 0.001751155, 
    0.001751155, 0.001751156, 0.001751147, 0.001751149, 0.001751147, 
    0.001751148, 0.001751193, 0.001751191, 0.001751192, 0.00175119, 
    0.001751192, 0.001751185, 0.001751182, 0.001751172, 0.001751177, 
    0.00175117, 0.001751176, 0.001751175, 0.00175117, 0.001751176, 
    0.001751163, 0.001751172, 0.001751156, 0.001751164, 0.001751155, 
    0.001751157, 0.001751154, 0.001751152, 0.001751148, 0.001751143, 
    0.001751144, 0.001751139, 0.001751188, 0.001751185, 0.001751185, 
    0.001751182, 0.00175118, 0.001751175, 0.001751167, 0.00175117, 
    0.001751165, 0.001751164, 0.001751172, 0.001751167, 0.001751183, 
    0.00175118, 0.001751182, 0.001751188, 0.001751169, 0.001751179, 
    0.001751162, 0.001751167, 0.001751152, 0.001751159, 0.001751145, 
    0.001751139, 0.001751133, 0.001751126, 0.001751183, 0.001751185, 
    0.001751182, 0.001751177, 0.001751172, 0.001751166, 0.001751166, 
    0.001751165, 0.001751162, 0.001751159, 0.001751164, 0.001751159, 
    0.00175118, 0.001751169, 0.001751186, 0.001751181, 0.001751177, 
    0.001751179, 0.00175117, 0.001751169, 0.001751161, 0.001751165, 
    0.00175114, 0.001751151, 0.001751121, 0.00175113, 0.001751186, 
    0.001751183, 0.001751174, 0.001751179, 0.001751166, 0.001751163, 
    0.00175116, 0.001751157, 0.001751157, 0.001751155, 0.001751158, 
    0.001751155, 0.001751166, 0.001751161, 0.001751175, 0.001751172, 
    0.001751173, 0.001751175, 0.00175117, 0.001751164, 0.001751164, 
    0.001751162, 0.001751157, 0.001751166, 0.001751139, 0.001751155, 
    0.001751181, 0.001751175, 0.001751175, 0.001751177, 0.001751163, 
    0.001751168, 0.001751155, 0.001751158, 0.001751153, 0.001751155, 
    0.001751156, 0.00175116, 0.001751162, 0.001751168, 0.001751172, 
    0.001751176, 0.001751175, 0.001751171, 0.001751164, 0.001751157, 
    0.001751158, 0.001751153, 0.001751167, 0.001751161, 0.001751163, 
    0.001751157, 0.00175117, 0.001751159, 0.001751173, 0.001751172, 
    0.001751168, 0.001751161, 0.001751159, 0.001751157, 0.001751158, 
    0.001751164, 0.001751164, 0.001751168, 0.001751169, 0.001751172, 
    0.001751174, 0.001751172, 0.00175117, 0.001751164, 0.001751158, 
    0.001751152, 0.00175115, 0.001751143, 0.001751149, 0.001751139, 
    0.001751147, 0.001751133, 0.001751159, 0.001751147, 0.001751168, 
    0.001751166, 0.001751162, 0.001751153, 0.001751157, 0.001751152, 
    0.001751164, 0.001751171, 0.001751173, 0.001751176, 0.001751173, 
    0.001751173, 0.00175117, 0.001751171, 0.001751163, 0.001751167, 
    0.001751156, 0.001751152, 0.00175114, 0.001751133, 0.001751125, 
    0.001751122, 0.001751121, 0.001751121,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.733029e-07, 9.732992e-07, 9.732998e-07, 9.732968e-07, 9.732985e-07, 
    9.732966e-07, 9.733021e-07, 9.732989e-07, 9.73301e-07, 9.733026e-07, 
    9.73291e-07, 9.732967e-07, 9.732851e-07, 9.732887e-07, 9.732796e-07, 
    9.732856e-07, 9.732784e-07, 9.732797e-07, 9.732755e-07, 9.732768e-07, 
    9.732714e-07, 9.73275e-07, 9.732686e-07, 9.732722e-07, 9.732717e-07, 
    9.732751e-07, 9.732955e-07, 9.732917e-07, 9.732958e-07, 9.732952e-07, 
    9.732955e-07, 9.732985e-07, 9.733e-07, 9.733031e-07, 9.733026e-07, 
    9.733003e-07, 9.73295e-07, 9.732968e-07, 9.732922e-07, 9.732923e-07, 
    9.732873e-07, 9.732896e-07, 9.732812e-07, 9.732836e-07, 9.732767e-07, 
    9.732785e-07, 9.732768e-07, 9.732772e-07, 9.732768e-07, 9.732793e-07, 
    9.732782e-07, 9.732804e-07, 9.732892e-07, 9.732867e-07, 9.732943e-07, 
    9.732989e-07, 9.73302e-07, 9.733042e-07, 9.733038e-07, 9.733033e-07, 
    9.733002e-07, 9.732973e-07, 9.732952e-07, 9.732938e-07, 9.732923e-07, 
    9.732881e-07, 9.732858e-07, 9.732807e-07, 9.732817e-07, 9.732801e-07, 
    9.732786e-07, 9.732761e-07, 9.732765e-07, 9.732754e-07, 9.732802e-07, 
    9.73277e-07, 9.732821e-07, 9.732807e-07, 9.73292e-07, 9.732963e-07, 
    9.732981e-07, 9.732997e-07, 9.733036e-07, 9.733009e-07, 9.73302e-07, 
    9.732995e-07, 9.732978e-07, 9.732986e-07, 9.732937e-07, 9.732956e-07, 
    9.732856e-07, 9.7329e-07, 9.732788e-07, 9.732814e-07, 9.732781e-07, 
    9.732798e-07, 9.732769e-07, 9.732795e-07, 9.732751e-07, 9.73274e-07, 
    9.732747e-07, 9.732721e-07, 9.732797e-07, 9.732768e-07, 9.732987e-07, 
    9.732985e-07, 9.732979e-07, 9.733005e-07, 9.733008e-07, 9.733031e-07, 
    9.73301e-07, 9.733001e-07, 9.732978e-07, 9.732964e-07, 9.732951e-07, 
    9.732922e-07, 9.732889e-07, 9.732845e-07, 9.732813e-07, 9.732792e-07, 
    9.732804e-07, 9.732793e-07, 9.732806e-07, 9.732812e-07, 9.732744e-07, 
    9.732782e-07, 9.732724e-07, 9.732728e-07, 9.732754e-07, 9.732728e-07, 
    9.732985e-07, 9.732992e-07, 9.733018e-07, 9.732997e-07, 9.733035e-07, 
    9.733013e-07, 9.733002e-07, 9.732956e-07, 9.732946e-07, 9.732937e-07, 
    9.732919e-07, 9.732895e-07, 9.732854e-07, 9.732818e-07, 9.732785e-07, 
    9.732787e-07, 9.732787e-07, 9.732779e-07, 9.732797e-07, 9.732777e-07, 
    9.732773e-07, 9.732782e-07, 9.732729e-07, 9.732744e-07, 9.732728e-07, 
    9.732738e-07, 9.732989e-07, 9.732977e-07, 9.732984e-07, 9.732971e-07, 
    9.73298e-07, 9.73294e-07, 9.732928e-07, 9.732872e-07, 9.732895e-07, 
    9.732859e-07, 9.732892e-07, 9.732886e-07, 9.732858e-07, 9.73289e-07, 
    9.73282e-07, 9.732868e-07, 9.732779e-07, 9.732827e-07, 9.732776e-07, 
    9.732785e-07, 9.73277e-07, 9.732756e-07, 9.732739e-07, 9.732709e-07, 
    9.732715e-07, 9.732689e-07, 9.732959e-07, 9.732942e-07, 9.732944e-07, 
    9.732927e-07, 9.732914e-07, 9.732887e-07, 9.732844e-07, 9.73286e-07, 
    9.73283e-07, 9.732823e-07, 9.732869e-07, 9.732842e-07, 9.732931e-07, 
    9.732917e-07, 9.732926e-07, 9.732958e-07, 9.732856e-07, 9.732908e-07, 
    9.732812e-07, 9.73284e-07, 9.732759e-07, 9.7328e-07, 9.73272e-07, 
    9.732686e-07, 9.732653e-07, 9.732616e-07, 9.732934e-07, 9.732944e-07, 
    9.732925e-07, 9.732897e-07, 9.732872e-07, 9.732838e-07, 9.732835e-07, 
    9.732829e-07, 9.732812e-07, 9.732798e-07, 9.732827e-07, 9.732795e-07, 
    9.732913e-07, 9.732852e-07, 9.732948e-07, 9.732919e-07, 9.732898e-07, 
    9.732908e-07, 9.732862e-07, 9.732851e-07, 9.732806e-07, 9.732829e-07, 
    9.732694e-07, 9.732754e-07, 9.732588e-07, 9.732634e-07, 9.732948e-07, 
    9.732934e-07, 9.732881e-07, 9.732906e-07, 9.732836e-07, 9.732819e-07, 
    9.732805e-07, 9.732787e-07, 9.732785e-07, 9.732775e-07, 9.732792e-07, 
    9.732776e-07, 9.732838e-07, 9.73281e-07, 9.732888e-07, 9.732869e-07, 
    9.732878e-07, 9.732887e-07, 9.732858e-07, 9.732827e-07, 9.732826e-07, 
    9.732815e-07, 9.732787e-07, 9.732836e-07, 9.732686e-07, 9.732779e-07, 
    9.732917e-07, 9.732888e-07, 9.732885e-07, 9.732896e-07, 9.732821e-07, 
    9.732848e-07, 9.732775e-07, 9.732795e-07, 9.732762e-07, 9.732778e-07, 
    9.732781e-07, 9.732802e-07, 9.732814e-07, 9.732846e-07, 9.732873e-07, 
    9.732894e-07, 9.732889e-07, 9.732867e-07, 9.732825e-07, 9.732785e-07, 
    9.732794e-07, 9.732764e-07, 9.732842e-07, 9.73281e-07, 9.732821e-07, 
    9.732789e-07, 9.73286e-07, 9.7328e-07, 9.732876e-07, 9.732869e-07, 
    9.732848e-07, 9.732807e-07, 9.732798e-07, 9.732788e-07, 9.732794e-07, 
    9.732823e-07, 9.732828e-07, 9.732848e-07, 9.732855e-07, 9.73287e-07, 
    9.732884e-07, 9.732871e-07, 9.732859e-07, 9.732823e-07, 9.732792e-07, 
    9.732756e-07, 9.732748e-07, 9.732707e-07, 9.73274e-07, 9.732686e-07, 
    9.732732e-07, 9.732652e-07, 9.732796e-07, 9.732734e-07, 9.732847e-07, 
    9.732835e-07, 9.732813e-07, 9.732762e-07, 9.732789e-07, 9.732757e-07, 
    9.732828e-07, 9.732865e-07, 9.732875e-07, 9.732893e-07, 9.732875e-07, 
    9.732876e-07, 9.732859e-07, 9.732864e-07, 9.732822e-07, 9.732845e-07, 
    9.732781e-07, 9.732757e-07, 9.732692e-07, 9.732652e-07, 9.732611e-07, 
    9.732593e-07, 9.732587e-07, 9.732585e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  8.82326e-25, -6.372354e-26, 1.274471e-25, 1.176435e-25, -3.480286e-25, 
    1.960724e-26, -4.999847e-25, 8.431115e-25, -1.519561e-25, -1.56858e-25, 
    2.941087e-25, -1.911706e-25, 4.803775e-25, 1.960724e-26, -7.842898e-25, 
    -3.970467e-25, -1.078398e-25, -3.921449e-26, -9.803622e-27, 
    -4.117521e-25, -3.823413e-25, 4.999847e-25, -2.548942e-25, 1.862688e-25, 
    9.803622e-26, 3.039123e-25, -4.41163e-26, -2.352869e-25, 2.843051e-25, 
    2.254833e-25, -3.578322e-25, -5.588064e-25, 2.450906e-25, 3.333231e-25, 
    9.166386e-25, -1.372507e-25, -3.333231e-25, -6.862535e-26, 5.244938e-25, 
    -2.646978e-25, -4.901811e-26, -3.431268e-26, 9.803622e-27, 4.705739e-25, 
    -4.607703e-25, 3.774394e-25, 6.764499e-25, 2.941087e-26, 9.460495e-25, 
    8.333079e-26, 2.646978e-25, 3.431268e-25, 6.274318e-25, -3.921449e-26, 
    1.02938e-25, -3.725376e-25, -4.607703e-25, -6.862535e-26, -2.941087e-25, 
    2.058761e-25, 3.774394e-25, 1.078398e-25, -1.666616e-25, -2.941087e-25, 
    -4.901811e-26, 9.117368e-25, -1.009773e-24, 4.901811e-27, -5.98021e-25, 
    4.41163e-25, 1.176435e-25, 6.960572e-25, 9.803622e-26, 1.421525e-25, 
    -5.490028e-25, 6.176282e-25, -3.823413e-25, -3.921449e-26, 4.803775e-25, 
    -2.401887e-25, -1.098006e-24, -2.058761e-25, -1.323489e-25, 
    -1.666616e-25, -4.019485e-25, 1.421525e-25, 4.901811e-25, -3.921449e-26, 
    6.122413e-41, -1.196042e-24, 1.235256e-24, 5.391992e-26, 5.146902e-25, 
    -3.480286e-25, 2.058761e-25, 7.058608e-25, 3.529304e-25, 1.176435e-25, 
    5.637083e-25, -2.745014e-25, 1.147024e-24, -9.803622e-26, 6.862535e-26, 
    -1.715634e-25, -4.901811e-26, 3.62734e-25, -3.235195e-25, 1.607794e-24, 
    9.803622e-27, -7.940934e-25, -7.401734e-25, -4.607703e-25, -1.078398e-25, 
    4.313593e-25, 2.548942e-25, -2.058761e-25, 1.323489e-25, 3.431268e-25, 
    4.999847e-25, 6.029227e-25, 3.088141e-25, 4.509666e-25, -2.156797e-25, 
    2.941087e-25, -8.82326e-26, -4.019485e-25, -4.999847e-25, -1.764652e-25, 
    2.254833e-25, 5.490028e-25, 4.019485e-25, 1.666616e-25, 5.490028e-25, 
    1.519561e-25, -5.784137e-25, 2.450906e-25, 4.019485e-25, 2.941087e-26, 
    -6.176282e-25, -1.274471e-25, 1.519561e-25, 6.176282e-25, -4.754757e-25, 
    2.107779e-25, -2.745014e-25, -3.137159e-25, -1.127417e-25, 6.127264e-25, 
    -2.156797e-25, -3.725376e-25, 3.62734e-25, 5.882173e-26, 1.911706e-25, 
    3.431268e-26, 1.470543e-25, 6.862535e-25, -2.941087e-25, 7.205662e-25, 
    -4.313593e-25, 3.921449e-25, -5.833155e-25, 1.960724e-25, -1.372507e-25, 
    8.82326e-26, 6.764499e-25, 5.19592e-25, -7.548789e-25, 5.048866e-25, 
    -3.823413e-25, 2.107779e-25, -7.842898e-25, -4.215557e-25, -9.019333e-25, 
    1.519561e-25, -5.342974e-25, 3.431268e-26, 4.117521e-25, -4.705739e-25, 
    3.431268e-26, -1.764652e-25, 1.862688e-25, 3.137159e-25, 2.352869e-25, 
    -6.519409e-25, -2.646978e-25, -1.274471e-25, 1.764652e-25, -3.137159e-25, 
    0, 4.607703e-25, 2.745014e-25, -5.293956e-25, 7.058608e-25, 3.921449e-26, 
    5.931191e-25, 6.911554e-25, -6.122413e-41, -3.529304e-25, 4.901811e-27, 
    -9.803622e-27, -4.117521e-25, -1.058791e-24, -1.56858e-25, 5.882173e-25, 
    -3.676358e-25, -4.901811e-25, -2.941087e-25, -3.725376e-25, 5.19592e-25, 
    1.960724e-26, -3.137159e-25, 1.862688e-25, -2.941087e-25, 7.744861e-25, 
    -6.078246e-25, 6.274318e-25, 3.872431e-25, 8.235043e-25, -3.529304e-25, 
    -3.039123e-25, -1.470543e-25, 6.372354e-26, 6.029227e-25, -3.921449e-26, 
    -2.499924e-25, 9.313441e-26, -3.725376e-25, -4.509666e-25, 3.235195e-25, 
    4.705739e-25, 3.039123e-25, -1.044086e-24, -3.529304e-25, 3.725376e-25, 
    3.235195e-25, 4.509666e-25, -4.705739e-25, 8.03897e-25, 7.107626e-25, 
    -6.862535e-26, 8.333079e-26, -2.941087e-25, 1.176435e-25, 1.862688e-25, 
    -2.745014e-25, 1.039184e-24, -5.391992e-26, -4.705739e-25, -3.872431e-25, 
    2.646978e-25, 9.950677e-25, 5.784137e-25, 2.941087e-25, -6.274318e-25, 
    1.862688e-25, 4.901811e-27, -4.509666e-25, 4.068503e-25, 1.078398e-25, 
    3.823413e-25, -2.548942e-25, -6.862535e-26, 6.323336e-25, 6.519409e-25, 
    -1.960724e-25, -3.039123e-25, 2.745014e-25, -5.882173e-26, 3.62734e-25, 
    -9.313441e-25, -3.137159e-25, -1.960724e-26, -1.911706e-25, 6.666463e-25, 
    -3.137159e-25, 7.058608e-25, 2.843051e-25, -1.274471e-25, -7.548789e-25, 
    3.921449e-25, -4.019485e-25, 4.705739e-25, -2.695996e-25, 1.573481e-24, 
    4.215557e-25, 5.588064e-25, -7.499771e-25, 5.146902e-25, 2.745014e-25, 
    8.333079e-26, 4.901811e-27, -3.137159e-25, 1.098006e-24, -1.81367e-25, 
    5.490028e-25, 4.901811e-25, -2.058761e-25, 9.411477e-25, 1.56858e-25, 
    -1.470543e-25, 1.372507e-25, -3.823413e-25, 1.764652e-25, 4.264576e-25, 
    -2.352869e-25, -5.784137e-25, 1.088202e-24, 6.372354e-26, 1.225453e-25, 
    -2.058761e-25, -4.901811e-25, 9.754604e-25, 3.235195e-25, -1.715634e-25, 
    3.62734e-25, 4.166539e-25, 3.676358e-25, 5.19592e-25, 3.039123e-25, 
    3.921449e-25, 1.960724e-25, -2.499924e-25, 6.372354e-25, -1.470543e-26, 
    -1.313685e-24, 5.882173e-26, -6.764499e-25, 5.588064e-25, 1.078398e-25, 
    -6.47039e-25, 4.754757e-25, -3.823413e-25, 2.548942e-25, -6.862535e-25, 
    -1.519561e-25, 1.666616e-25, 8.235043e-25, -2.303851e-25,
  9.436869e-32, 9.436832e-32, 9.436839e-32, 9.436809e-32, 9.436825e-32, 
    9.436806e-32, 9.436862e-32, 9.43683e-32, 9.43685e-32, 9.436866e-32, 
    9.43675e-32, 9.436807e-32, 9.43669e-32, 9.436727e-32, 9.436635e-32, 
    9.436696e-32, 9.436623e-32, 9.436637e-32, 9.436595e-32, 9.436607e-32, 
    9.436553e-32, 9.436589e-32, 9.436525e-32, 9.436561e-32, 9.436556e-32, 
    9.43659e-32, 9.436796e-32, 9.436757e-32, 9.436798e-32, 9.436792e-32, 
    9.436795e-32, 9.436825e-32, 9.43684e-32, 9.436872e-32, 9.436866e-32, 
    9.436843e-32, 9.43679e-32, 9.436808e-32, 9.436763e-32, 9.436763e-32, 
    9.436713e-32, 9.436736e-32, 9.436652e-32, 9.436675e-32, 9.436606e-32, 
    9.436624e-32, 9.436607e-32, 9.436612e-32, 9.436607e-32, 9.436632e-32, 
    9.436622e-32, 9.436644e-32, 9.436732e-32, 9.436706e-32, 9.436783e-32, 
    9.436829e-32, 9.43686e-32, 9.436882e-32, 9.436879e-32, 9.436873e-32, 
    9.436843e-32, 9.436814e-32, 9.436792e-32, 9.436778e-32, 9.436764e-32, 
    9.436721e-32, 9.436698e-32, 9.436646e-32, 9.436656e-32, 9.43664e-32, 
    9.436625e-32, 9.4366e-32, 9.436604e-32, 9.436594e-32, 9.436641e-32, 
    9.436609e-32, 9.436661e-32, 9.436647e-32, 9.43676e-32, 9.436803e-32, 
    9.436822e-32, 9.436837e-32, 9.436876e-32, 9.436849e-32, 9.43686e-32, 
    9.436835e-32, 9.436819e-32, 9.436827e-32, 9.436778e-32, 9.436797e-32, 
    9.436696e-32, 9.436739e-32, 9.436627e-32, 9.436654e-32, 9.436621e-32, 
    9.436638e-32, 9.436608e-32, 9.436635e-32, 9.436589e-32, 9.436579e-32, 
    9.436586e-32, 9.43656e-32, 9.436636e-32, 9.436607e-32, 9.436827e-32, 
    9.436826e-32, 9.43682e-32, 9.436846e-32, 9.436848e-32, 9.436872e-32, 
    9.43685e-32, 9.436841e-32, 9.436818e-32, 9.436804e-32, 9.436791e-32, 
    9.436762e-32, 9.436729e-32, 9.436685e-32, 9.436652e-32, 9.436631e-32, 
    9.436644e-32, 9.436632e-32, 9.436645e-32, 9.436651e-32, 9.436583e-32, 
    9.436621e-32, 9.436564e-32, 9.436567e-32, 9.436593e-32, 9.436567e-32, 
    9.436825e-32, 9.436832e-32, 9.436858e-32, 9.436838e-32, 9.436875e-32, 
    9.436854e-32, 9.436842e-32, 9.436796e-32, 9.436786e-32, 9.436777e-32, 
    9.436759e-32, 9.436735e-32, 9.436693e-32, 9.436657e-32, 9.436625e-32, 
    9.436627e-32, 9.436626e-32, 9.436619e-32, 9.436637e-32, 9.436616e-32, 
    9.436612e-32, 9.436621e-32, 9.436568e-32, 9.436583e-32, 9.436567e-32, 
    9.436577e-32, 9.43683e-32, 9.436817e-32, 9.436824e-32, 9.436811e-32, 
    9.43682e-32, 9.43678e-32, 9.436768e-32, 9.436712e-32, 9.436735e-32, 
    9.436699e-32, 9.436732e-32, 9.436726e-32, 9.436698e-32, 9.43673e-32, 
    9.436659e-32, 9.436707e-32, 9.436618e-32, 9.436666e-32, 9.436615e-32, 
    9.436625e-32, 9.436609e-32, 9.436596e-32, 9.436579e-32, 9.436547e-32, 
    9.436554e-32, 9.436528e-32, 9.436799e-32, 9.436782e-32, 9.436783e-32, 
    9.436766e-32, 9.436754e-32, 9.436727e-32, 9.436683e-32, 9.436699e-32, 
    9.436669e-32, 9.436664e-32, 9.436709e-32, 9.436681e-32, 9.436771e-32, 
    9.436757e-32, 9.436765e-32, 9.436797e-32, 9.436696e-32, 9.436748e-32, 
    9.436652e-32, 9.43668e-32, 9.436598e-32, 9.436638e-32, 9.436558e-32, 
    9.436524e-32, 9.436492e-32, 9.436455e-32, 9.436773e-32, 9.436785e-32, 
    9.436765e-32, 9.436737e-32, 9.436712e-32, 9.436678e-32, 9.436675e-32, 
    9.436668e-32, 9.436652e-32, 9.436638e-32, 9.436666e-32, 9.436635e-32, 
    9.436753e-32, 9.436691e-32, 9.436789e-32, 9.436759e-32, 9.436739e-32, 
    9.436748e-32, 9.436701e-32, 9.436691e-32, 9.436646e-32, 9.436669e-32, 
    9.436532e-32, 9.436593e-32, 9.436426e-32, 9.436473e-32, 9.436788e-32, 
    9.436773e-32, 9.436722e-32, 9.436746e-32, 9.436676e-32, 9.436659e-32, 
    9.436645e-32, 9.436626e-32, 9.436625e-32, 9.436614e-32, 9.436631e-32, 
    9.436615e-32, 9.436678e-32, 9.436649e-32, 9.436728e-32, 9.436709e-32, 
    9.436717e-32, 9.436727e-32, 9.436698e-32, 9.436666e-32, 9.436665e-32, 
    9.436655e-32, 9.436627e-32, 9.436676e-32, 9.436525e-32, 9.436618e-32, 
    9.436757e-32, 9.436729e-32, 9.436725e-32, 9.436735e-32, 9.436661e-32, 
    9.436688e-32, 9.436614e-32, 9.436634e-32, 9.436602e-32, 9.436618e-32, 
    9.43662e-32, 9.436641e-32, 9.436654e-32, 9.436686e-32, 9.436713e-32, 
    9.436734e-32, 9.436729e-32, 9.436706e-32, 9.436664e-32, 9.436625e-32, 
    9.436633e-32, 9.436604e-32, 9.436681e-32, 9.436649e-32, 9.436661e-32, 
    9.436629e-32, 9.4367e-32, 9.436639e-32, 9.436715e-32, 9.436709e-32, 
    9.436688e-32, 9.436646e-32, 9.436637e-32, 9.436628e-32, 9.436634e-32, 
    9.436663e-32, 9.436668e-32, 9.436689e-32, 9.436694e-32, 9.43671e-32, 
    9.436723e-32, 9.436711e-32, 9.436699e-32, 9.436663e-32, 9.436631e-32, 
    9.436595e-32, 9.436587e-32, 9.436546e-32, 9.436579e-32, 9.436524e-32, 
    9.436571e-32, 9.43649e-32, 9.436636e-32, 9.436572e-32, 9.436687e-32, 
    9.436675e-32, 9.436652e-32, 9.436601e-32, 9.436629e-32, 9.436597e-32, 
    9.436668e-32, 9.436705e-32, 9.436715e-32, 9.436733e-32, 9.436714e-32, 
    9.436716e-32, 9.436698e-32, 9.436704e-32, 9.436662e-32, 9.436684e-32, 
    9.43662e-32, 9.436597e-32, 9.436531e-32, 9.43649e-32, 9.43645e-32, 
    9.436431e-32, 9.436425e-32, 9.436424e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.533999e-14, 4.546242e-14, 4.543864e-14, 4.553729e-14, 4.548259e-14, 
    4.554716e-14, 4.536483e-14, 4.546726e-14, 4.540189e-14, 4.535104e-14, 
    4.572844e-14, 4.554169e-14, 4.592225e-14, 4.580336e-14, 4.61018e-14, 
    4.590373e-14, 4.61417e-14, 4.609613e-14, 4.623332e-14, 4.619404e-14, 
    4.636924e-14, 4.625144e-14, 4.646e-14, 4.634114e-14, 4.635973e-14, 
    4.624755e-14, 4.557933e-14, 4.57052e-14, 4.557186e-14, 4.558982e-14, 
    4.558177e-14, 4.54837e-14, 4.543423e-14, 4.533065e-14, 4.534947e-14, 
    4.542555e-14, 4.55979e-14, 4.553945e-14, 4.568677e-14, 4.568344e-14, 
    4.584721e-14, 4.57734e-14, 4.604831e-14, 4.597025e-14, 4.619568e-14, 
    4.613902e-14, 4.619301e-14, 4.617665e-14, 4.619322e-14, 4.611013e-14, 
    4.614573e-14, 4.60726e-14, 4.578722e-14, 4.587116e-14, 4.562061e-14, 
    4.546963e-14, 4.536932e-14, 4.529807e-14, 4.530814e-14, 4.532734e-14, 
    4.5426e-14, 4.551871e-14, 4.55893e-14, 4.563649e-14, 4.568297e-14, 
    4.582345e-14, 4.589781e-14, 4.606406e-14, 4.603411e-14, 4.608487e-14, 
    4.613339e-14, 4.621475e-14, 4.620137e-14, 4.623719e-14, 4.608356e-14, 
    4.618568e-14, 4.601704e-14, 4.606318e-14, 4.569548e-14, 4.555522e-14, 
    4.549545e-14, 4.54432e-14, 4.531589e-14, 4.540382e-14, 4.536916e-14, 
    4.545162e-14, 4.550397e-14, 4.547809e-14, 4.563778e-14, 4.557572e-14, 
    4.590221e-14, 4.57617e-14, 4.612773e-14, 4.604026e-14, 4.614869e-14, 
    4.609338e-14, 4.618812e-14, 4.610286e-14, 4.625053e-14, 4.628265e-14, 
    4.62607e-14, 4.634502e-14, 4.609813e-14, 4.6193e-14, 4.547735e-14, 
    4.548158e-14, 4.550125e-14, 4.541473e-14, 4.540944e-14, 4.533013e-14, 
    4.540072e-14, 4.543075e-14, 4.550701e-14, 4.555207e-14, 4.55949e-14, 
    4.5689e-14, 4.579399e-14, 4.594066e-14, 4.604593e-14, 4.611643e-14, 
    4.607322e-14, 4.611137e-14, 4.606871e-14, 4.604872e-14, 4.62706e-14, 
    4.614606e-14, 4.63329e-14, 4.632257e-14, 4.623804e-14, 4.632373e-14, 
    4.548454e-14, 4.546025e-14, 4.537582e-14, 4.544189e-14, 4.532149e-14, 
    4.538889e-14, 4.542761e-14, 4.557699e-14, 4.560981e-14, 4.56402e-14, 
    4.570021e-14, 4.577718e-14, 4.591205e-14, 4.602929e-14, 4.613621e-14, 
    4.612839e-14, 4.613114e-14, 4.6155e-14, 4.609587e-14, 4.616471e-14, 
    4.617625e-14, 4.614606e-14, 4.632119e-14, 4.627119e-14, 4.632235e-14, 
    4.62898e-14, 4.546815e-14, 4.550903e-14, 4.548694e-14, 4.552846e-14, 
    4.54992e-14, 4.562924e-14, 4.56682e-14, 4.585034e-14, 4.577566e-14, 
    4.589453e-14, 4.578775e-14, 4.580667e-14, 4.589835e-14, 4.579353e-14, 
    4.60228e-14, 4.586737e-14, 4.615593e-14, 4.600086e-14, 4.616564e-14, 
    4.613575e-14, 4.618524e-14, 4.622953e-14, 4.628524e-14, 4.638792e-14, 
    4.636416e-14, 4.644999e-14, 4.556996e-14, 4.562292e-14, 4.561828e-14, 
    4.567369e-14, 4.571465e-14, 4.580341e-14, 4.594558e-14, 4.589215e-14, 
    4.599025e-14, 4.600993e-14, 4.586089e-14, 4.59524e-14, 4.565837e-14, 
    4.57059e-14, 4.567762e-14, 4.557412e-14, 4.590444e-14, 4.573503e-14, 
    4.604767e-14, 4.595605e-14, 4.622321e-14, 4.609041e-14, 4.635107e-14, 
    4.646224e-14, 4.656686e-14, 4.668886e-14, 4.565183e-14, 4.561586e-14, 
    4.568029e-14, 4.576933e-14, 4.585194e-14, 4.596164e-14, 4.597287e-14, 
    4.59934e-14, 4.604658e-14, 4.609127e-14, 4.599987e-14, 4.610247e-14, 
    4.571688e-14, 4.591914e-14, 4.560223e-14, 4.569773e-14, 4.576409e-14, 
    4.573501e-14, 4.588605e-14, 4.592161e-14, 4.606598e-14, 4.599139e-14, 
    4.643479e-14, 4.623885e-14, 4.678173e-14, 4.66303e-14, 4.560328e-14, 
    4.565172e-14, 4.582012e-14, 4.574003e-14, 4.596897e-14, 4.602524e-14, 
    4.607098e-14, 4.612938e-14, 4.61357e-14, 4.617029e-14, 4.61136e-14, 
    4.616806e-14, 4.596187e-14, 4.605407e-14, 4.580091e-14, 4.586257e-14, 
    4.583422e-14, 4.580309e-14, 4.589912e-14, 4.60013e-14, 4.600352e-14, 
    4.603625e-14, 4.612838e-14, 4.59699e-14, 4.645998e-14, 4.615753e-14, 
    4.570452e-14, 4.579767e-14, 4.581101e-14, 4.577493e-14, 4.601959e-14, 
    4.593101e-14, 4.616945e-14, 4.610507e-14, 4.621055e-14, 4.615814e-14, 
    4.615043e-14, 4.608309e-14, 4.604113e-14, 4.593506e-14, 4.584869e-14, 
    4.578017e-14, 4.579611e-14, 4.587137e-14, 4.600755e-14, 4.613625e-14, 
    4.610807e-14, 4.620254e-14, 4.595238e-14, 4.605733e-14, 4.601677e-14, 
    4.612251e-14, 4.589072e-14, 4.608802e-14, 4.584022e-14, 4.586198e-14, 
    4.592925e-14, 4.606442e-14, 4.609436e-14, 4.612625e-14, 4.610658e-14, 
    4.601102e-14, 4.599537e-14, 4.592762e-14, 4.590889e-14, 4.585724e-14, 
    4.581445e-14, 4.585354e-14, 4.589457e-14, 4.601107e-14, 4.611593e-14, 
    4.623015e-14, 4.62581e-14, 4.639127e-14, 4.628283e-14, 4.646166e-14, 
    4.630956e-14, 4.657275e-14, 4.60995e-14, 4.630516e-14, 4.593232e-14, 
    4.597256e-14, 4.604526e-14, 4.62119e-14, 4.612201e-14, 4.622715e-14, 
    4.599476e-14, 4.587395e-14, 4.584271e-14, 4.578433e-14, 4.584404e-14, 
    4.583919e-14, 4.589629e-14, 4.587795e-14, 4.601494e-14, 4.594138e-14, 
    4.615023e-14, 4.622633e-14, 4.644098e-14, 4.657233e-14, 4.670591e-14, 
    4.676481e-14, 4.678273e-14, 4.679022e-14 ;

 LITR1N_vr =
  5.55766e-05, 5.557639e-05, 5.557643e-05, 5.557626e-05, 5.557635e-05, 
    5.557624e-05, 5.557655e-05, 5.557638e-05, 5.557649e-05, 5.557658e-05, 
    5.557592e-05, 5.557625e-05, 5.557558e-05, 5.557579e-05, 5.557527e-05, 
    5.557562e-05, 5.55752e-05, 5.557528e-05, 5.557504e-05, 5.557511e-05, 
    5.55748e-05, 5.557501e-05, 5.557464e-05, 5.557485e-05, 5.557482e-05, 
    5.557502e-05, 5.557618e-05, 5.557596e-05, 5.557619e-05, 5.557616e-05, 
    5.557618e-05, 5.557635e-05, 5.557643e-05, 5.557662e-05, 5.557658e-05, 
    5.557645e-05, 5.557615e-05, 5.557625e-05, 5.557599e-05, 5.5576e-05, 
    5.557571e-05, 5.557584e-05, 5.557536e-05, 5.55755e-05, 5.557511e-05, 
    5.55752e-05, 5.557511e-05, 5.557514e-05, 5.557511e-05, 5.557526e-05, 
    5.557519e-05, 5.557532e-05, 5.557582e-05, 5.557567e-05, 5.557611e-05, 
    5.557637e-05, 5.557655e-05, 5.557667e-05, 5.557666e-05, 5.557662e-05, 
    5.557645e-05, 5.557629e-05, 5.557617e-05, 5.557608e-05, 5.5576e-05, 
    5.557575e-05, 5.557563e-05, 5.557534e-05, 5.557539e-05, 5.55753e-05, 
    5.557521e-05, 5.557507e-05, 5.55751e-05, 5.557503e-05, 5.55753e-05, 
    5.557512e-05, 5.557542e-05, 5.557534e-05, 5.557598e-05, 5.557622e-05, 
    5.557633e-05, 5.557642e-05, 5.557664e-05, 5.557649e-05, 5.557655e-05, 
    5.557641e-05, 5.557631e-05, 5.557636e-05, 5.557608e-05, 5.557619e-05, 
    5.557562e-05, 5.557586e-05, 5.557522e-05, 5.557538e-05, 5.557519e-05, 
    5.557528e-05, 5.557512e-05, 5.557527e-05, 5.557501e-05, 5.557495e-05, 
    5.557499e-05, 5.557484e-05, 5.557527e-05, 5.557511e-05, 5.557636e-05, 
    5.557635e-05, 5.557632e-05, 5.557647e-05, 5.557648e-05, 5.557662e-05, 
    5.557649e-05, 5.557644e-05, 5.557631e-05, 5.557623e-05, 5.557615e-05, 
    5.557599e-05, 5.557581e-05, 5.557555e-05, 5.557536e-05, 5.557524e-05, 
    5.557532e-05, 5.557525e-05, 5.557532e-05, 5.557536e-05, 5.557498e-05, 
    5.557519e-05, 5.557487e-05, 5.557488e-05, 5.557503e-05, 5.557488e-05, 
    5.557635e-05, 5.557639e-05, 5.557654e-05, 5.557642e-05, 5.557663e-05, 
    5.557651e-05, 5.557645e-05, 5.557619e-05, 5.557613e-05, 5.557607e-05, 
    5.557597e-05, 5.557583e-05, 5.55756e-05, 5.557539e-05, 5.557521e-05, 
    5.557522e-05, 5.557522e-05, 5.557518e-05, 5.557528e-05, 5.557516e-05, 
    5.557514e-05, 5.557519e-05, 5.557488e-05, 5.557497e-05, 5.557488e-05, 
    5.557494e-05, 5.557638e-05, 5.55763e-05, 5.557634e-05, 5.557627e-05, 
    5.557632e-05, 5.557609e-05, 5.557603e-05, 5.557571e-05, 5.557584e-05, 
    5.557563e-05, 5.557582e-05, 5.557578e-05, 5.557562e-05, 5.557581e-05, 
    5.557541e-05, 5.557568e-05, 5.557518e-05, 5.557545e-05, 5.557516e-05, 
    5.557521e-05, 5.557512e-05, 5.557504e-05, 5.557495e-05, 5.557477e-05, 
    5.557481e-05, 5.557466e-05, 5.55762e-05, 5.557611e-05, 5.557611e-05, 
    5.557602e-05, 5.557594e-05, 5.557579e-05, 5.557554e-05, 5.557563e-05, 
    5.557546e-05, 5.557543e-05, 5.557569e-05, 5.557553e-05, 5.557605e-05, 
    5.557596e-05, 5.557601e-05, 5.557619e-05, 5.557561e-05, 5.557591e-05, 
    5.557536e-05, 5.557553e-05, 5.557506e-05, 5.557529e-05, 5.557483e-05, 
    5.557464e-05, 5.557446e-05, 5.557424e-05, 5.557606e-05, 5.557612e-05, 
    5.557601e-05, 5.557585e-05, 5.557571e-05, 5.557551e-05, 5.55755e-05, 
    5.557546e-05, 5.557536e-05, 5.557529e-05, 5.557545e-05, 5.557527e-05, 
    5.557594e-05, 5.557559e-05, 5.557614e-05, 5.557598e-05, 5.557586e-05, 
    5.557591e-05, 5.557565e-05, 5.557558e-05, 5.557533e-05, 5.557546e-05, 
    5.557469e-05, 5.557503e-05, 5.557408e-05, 5.557435e-05, 5.557614e-05, 
    5.557606e-05, 5.557576e-05, 5.55759e-05, 5.55755e-05, 5.55754e-05, 
    5.557532e-05, 5.557522e-05, 5.557521e-05, 5.557515e-05, 5.557525e-05, 
    5.557515e-05, 5.557551e-05, 5.557535e-05, 5.557579e-05, 5.557569e-05, 
    5.557574e-05, 5.557579e-05, 5.557562e-05, 5.557545e-05, 5.557544e-05, 
    5.557538e-05, 5.557522e-05, 5.55755e-05, 5.557464e-05, 5.557517e-05, 
    5.557596e-05, 5.55758e-05, 5.557578e-05, 5.557584e-05, 5.557541e-05, 
    5.557557e-05, 5.557515e-05, 5.557526e-05, 5.557508e-05, 5.557517e-05, 
    5.557518e-05, 5.55753e-05, 5.557538e-05, 5.557556e-05, 5.557571e-05, 
    5.557583e-05, 5.55758e-05, 5.557567e-05, 5.557543e-05, 5.557521e-05, 
    5.557526e-05, 5.557509e-05, 5.557553e-05, 5.557535e-05, 5.557542e-05, 
    5.557523e-05, 5.557564e-05, 5.557529e-05, 5.557573e-05, 5.557569e-05, 
    5.557557e-05, 5.557534e-05, 5.557528e-05, 5.557523e-05, 5.557526e-05, 
    5.557543e-05, 5.557546e-05, 5.557557e-05, 5.557561e-05, 5.55757e-05, 
    5.557577e-05, 5.55757e-05, 5.557563e-05, 5.557543e-05, 5.557524e-05, 
    5.557504e-05, 5.5575e-05, 5.557476e-05, 5.557495e-05, 5.557464e-05, 
    5.557491e-05, 5.557444e-05, 5.557527e-05, 5.557491e-05, 5.557557e-05, 
    5.55755e-05, 5.557537e-05, 5.557508e-05, 5.557523e-05, 5.557505e-05, 
    5.557546e-05, 5.557567e-05, 5.557572e-05, 5.557582e-05, 5.557572e-05, 
    5.557573e-05, 5.557563e-05, 5.557566e-05, 5.557542e-05, 5.557555e-05, 
    5.557518e-05, 5.557505e-05, 5.557468e-05, 5.557445e-05, 5.557422e-05, 
    5.557411e-05, 5.557408e-05, 5.557407e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.857573e-13, 7.87879e-13, 7.874669e-13, 7.891766e-13, 7.882286e-13, 
    7.893476e-13, 7.86188e-13, 7.87963e-13, 7.868302e-13, 7.859488e-13, 
    7.924893e-13, 7.892529e-13, 7.95848e-13, 7.937878e-13, 7.989598e-13, 
    7.955272e-13, 7.996513e-13, 7.988615e-13, 8.01239e-13, 8.005582e-13, 
    8.035945e-13, 8.015532e-13, 8.051675e-13, 8.031076e-13, 8.034297e-13, 
    8.014857e-13, 7.899053e-13, 7.920865e-13, 7.897758e-13, 7.90087e-13, 
    7.899475e-13, 7.88248e-13, 7.873906e-13, 7.855955e-13, 7.859216e-13, 
    7.872402e-13, 7.90227e-13, 7.89214e-13, 7.917672e-13, 7.917095e-13, 
    7.945476e-13, 7.932685e-13, 7.980327e-13, 7.9668e-13, 8.005867e-13, 
    7.996049e-13, 8.005405e-13, 8.002569e-13, 8.005441e-13, 7.991041e-13, 
    7.997212e-13, 7.984536e-13, 7.93508e-13, 7.949626e-13, 7.906206e-13, 
    7.88004e-13, 7.862657e-13, 7.850308e-13, 7.852054e-13, 7.855381e-13, 
    7.872479e-13, 7.888546e-13, 7.900779e-13, 7.908957e-13, 7.917012e-13, 
    7.941359e-13, 7.954245e-13, 7.983058e-13, 7.977866e-13, 7.986664e-13, 
    7.995072e-13, 8.009173e-13, 8.006853e-13, 8.013062e-13, 7.986436e-13, 
    8.004134e-13, 7.974908e-13, 7.982905e-13, 7.919181e-13, 7.894875e-13, 
    7.884516e-13, 7.875461e-13, 7.853396e-13, 7.868635e-13, 7.862629e-13, 
    7.87692e-13, 7.885992e-13, 7.881506e-13, 7.909181e-13, 7.898425e-13, 
    7.955009e-13, 7.930657e-13, 7.994091e-13, 7.978933e-13, 7.997724e-13, 
    7.988139e-13, 8.004558e-13, 7.989781e-13, 8.015373e-13, 8.020939e-13, 
    8.017135e-13, 8.031749e-13, 7.988962e-13, 8.005402e-13, 7.881379e-13, 
    7.882111e-13, 7.885521e-13, 7.870526e-13, 7.86961e-13, 7.855864e-13, 
    7.868097e-13, 7.873303e-13, 7.886519e-13, 7.894328e-13, 7.90175e-13, 
    7.918059e-13, 7.936253e-13, 7.961672e-13, 7.979916e-13, 7.992133e-13, 
    7.984644e-13, 7.991256e-13, 7.983864e-13, 7.980399e-13, 8.018852e-13, 
    7.997268e-13, 8.029647e-13, 8.027858e-13, 8.013208e-13, 8.02806e-13, 
    7.882625e-13, 7.878414e-13, 7.863782e-13, 7.875234e-13, 7.854367e-13, 
    7.866048e-13, 7.872759e-13, 7.898646e-13, 7.904334e-13, 7.9096e-13, 
    7.920001e-13, 7.933339e-13, 7.956714e-13, 7.977031e-13, 7.995562e-13, 
    7.994205e-13, 7.994683e-13, 7.998818e-13, 7.98857e-13, 8.0005e-13, 
    8.002499e-13, 7.997268e-13, 8.027618e-13, 8.018953e-13, 8.02782e-13, 
    8.022179e-13, 7.879784e-13, 7.886868e-13, 7.88304e-13, 7.890237e-13, 
    7.885166e-13, 7.907701e-13, 7.914453e-13, 7.94602e-13, 7.933076e-13, 
    7.953677e-13, 7.935171e-13, 7.938451e-13, 7.95434e-13, 7.936173e-13, 
    7.975907e-13, 7.94897e-13, 7.998979e-13, 7.972104e-13, 8.000661e-13, 
    7.995482e-13, 8.004058e-13, 8.011733e-13, 8.021388e-13, 8.039183e-13, 
    8.035065e-13, 8.04994e-13, 7.897427e-13, 7.906606e-13, 7.905802e-13, 
    7.915406e-13, 7.922504e-13, 7.937885e-13, 7.962525e-13, 7.953265e-13, 
    7.970266e-13, 7.973676e-13, 7.947848e-13, 7.963706e-13, 7.912749e-13, 
    7.920987e-13, 7.916085e-13, 7.898149e-13, 7.955394e-13, 7.926035e-13, 
    7.980216e-13, 7.964339e-13, 8.010639e-13, 7.987623e-13, 8.032796e-13, 
    8.052063e-13, 8.070194e-13, 8.091338e-13, 7.911617e-13, 7.905382e-13, 
    7.916548e-13, 7.931979e-13, 7.946296e-13, 7.965307e-13, 7.967253e-13, 
    7.970811e-13, 7.980028e-13, 7.987773e-13, 7.971932e-13, 7.989714e-13, 
    7.922889e-13, 7.957941e-13, 7.903021e-13, 7.91957e-13, 7.931071e-13, 
    7.926031e-13, 7.952207e-13, 7.95837e-13, 7.98339e-13, 7.970463e-13, 
    8.047306e-13, 8.013348e-13, 8.107433e-13, 8.081189e-13, 7.903202e-13, 
    7.911598e-13, 7.940781e-13, 7.926902e-13, 7.966578e-13, 7.976329e-13, 
    7.984256e-13, 7.994377e-13, 7.995473e-13, 8.001467e-13, 7.991643e-13, 
    8.001081e-13, 7.965348e-13, 7.981325e-13, 7.937452e-13, 7.948138e-13, 
    7.943225e-13, 7.93783e-13, 7.954473e-13, 7.97218e-13, 7.972565e-13, 
    7.978238e-13, 7.994204e-13, 7.966738e-13, 8.051672e-13, 7.999255e-13, 
    7.920747e-13, 7.936891e-13, 7.939204e-13, 7.932951e-13, 7.975352e-13, 
    7.959998e-13, 8.001322e-13, 7.990165e-13, 8.008444e-13, 7.999362e-13, 
    7.998026e-13, 7.986355e-13, 7.979084e-13, 7.960701e-13, 7.945733e-13, 
    7.933859e-13, 7.936621e-13, 7.949663e-13, 7.973265e-13, 7.995569e-13, 
    7.990684e-13, 8.007056e-13, 7.963703e-13, 7.981891e-13, 7.974862e-13, 
    7.993186e-13, 7.953017e-13, 7.98721e-13, 7.944265e-13, 7.948036e-13, 
    7.959694e-13, 7.983119e-13, 7.988308e-13, 7.993835e-13, 7.990426e-13, 
    7.973865e-13, 7.971153e-13, 7.959412e-13, 7.956166e-13, 7.947215e-13, 
    7.939798e-13, 7.946573e-13, 7.953684e-13, 7.973874e-13, 7.992047e-13, 
    8.011842e-13, 8.016685e-13, 8.039763e-13, 8.02097e-13, 8.051962e-13, 
    8.025603e-13, 8.071215e-13, 7.989198e-13, 8.02484e-13, 7.960226e-13, 
    7.967199e-13, 7.9798e-13, 8.008678e-13, 7.9931e-13, 8.011321e-13, 
    7.971047e-13, 7.95011e-13, 7.944696e-13, 7.93458e-13, 7.944928e-13, 
    7.944086e-13, 7.953983e-13, 7.950804e-13, 7.974544e-13, 7.961796e-13, 
    7.99799e-13, 8.011179e-13, 8.04838e-13, 8.071142e-13, 8.094292e-13, 
    8.1045e-13, 8.107606e-13, 8.108904e-13 ;

 LITR2C =
  1.939607e-05, 1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939605e-05, 
    1.939604e-05, 1.939607e-05, 1.939605e-05, 1.939606e-05, 1.939607e-05, 
    1.939601e-05, 1.939604e-05, 1.939598e-05, 1.939599e-05, 1.939595e-05, 
    1.939598e-05, 1.939594e-05, 1.939595e-05, 1.939593e-05, 1.939593e-05, 
    1.93959e-05, 1.939592e-05, 1.939589e-05, 1.939591e-05, 1.939591e-05, 
    1.939592e-05, 1.939603e-05, 1.939601e-05, 1.939603e-05, 1.939603e-05, 
    1.939603e-05, 1.939605e-05, 1.939605e-05, 1.939607e-05, 1.939607e-05, 
    1.939606e-05, 1.939603e-05, 1.939604e-05, 1.939601e-05, 1.939601e-05, 
    1.939599e-05, 1.9396e-05, 1.939596e-05, 1.939597e-05, 1.939593e-05, 
    1.939594e-05, 1.939593e-05, 1.939593e-05, 1.939593e-05, 1.939595e-05, 
    1.939594e-05, 1.939595e-05, 1.9396e-05, 1.939598e-05, 1.939603e-05, 
    1.939605e-05, 1.939607e-05, 1.939608e-05, 1.939608e-05, 1.939607e-05, 
    1.939606e-05, 1.939604e-05, 1.939603e-05, 1.939602e-05, 1.939601e-05, 
    1.939599e-05, 1.939598e-05, 1.939595e-05, 1.939596e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939593e-05, 1.939593e-05, 1.939595e-05, 
    1.939593e-05, 1.939596e-05, 1.939595e-05, 1.939601e-05, 1.939603e-05, 
    1.939605e-05, 1.939605e-05, 1.939608e-05, 1.939606e-05, 1.939607e-05, 
    1.939605e-05, 1.939604e-05, 1.939605e-05, 1.939602e-05, 1.939603e-05, 
    1.939598e-05, 1.9396e-05, 1.939594e-05, 1.939596e-05, 1.939594e-05, 
    1.939595e-05, 1.939593e-05, 1.939595e-05, 1.939592e-05, 1.939592e-05, 
    1.939592e-05, 1.939591e-05, 1.939595e-05, 1.939593e-05, 1.939605e-05, 
    1.939605e-05, 1.939604e-05, 1.939606e-05, 1.939606e-05, 1.939607e-05, 
    1.939606e-05, 1.939605e-05, 1.939604e-05, 1.939604e-05, 1.939603e-05, 
    1.939601e-05, 1.9396e-05, 1.939597e-05, 1.939596e-05, 1.939595e-05, 
    1.939595e-05, 1.939595e-05, 1.939595e-05, 1.939596e-05, 1.939592e-05, 
    1.939594e-05, 1.939591e-05, 1.939591e-05, 1.939593e-05, 1.939591e-05, 
    1.939605e-05, 1.939605e-05, 1.939606e-05, 1.939605e-05, 1.939607e-05, 
    1.939606e-05, 1.939606e-05, 1.939603e-05, 1.939603e-05, 1.939602e-05, 
    1.939601e-05, 1.9396e-05, 1.939598e-05, 1.939596e-05, 1.939594e-05, 
    1.939594e-05, 1.939594e-05, 1.939594e-05, 1.939595e-05, 1.939594e-05, 
    1.939593e-05, 1.939594e-05, 1.939591e-05, 1.939592e-05, 1.939591e-05, 
    1.939592e-05, 1.939605e-05, 1.939604e-05, 1.939605e-05, 1.939604e-05, 
    1.939604e-05, 1.939602e-05, 1.939602e-05, 1.939599e-05, 1.9396e-05, 
    1.939598e-05, 1.9396e-05, 1.939599e-05, 1.939598e-05, 1.9396e-05, 
    1.939596e-05, 1.939599e-05, 1.939594e-05, 1.939596e-05, 1.939594e-05, 
    1.939594e-05, 1.939593e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 
    1.939591e-05, 1.939589e-05, 1.939603e-05, 1.939602e-05, 1.939603e-05, 
    1.939602e-05, 1.939601e-05, 1.939599e-05, 1.939597e-05, 1.939598e-05, 
    1.939597e-05, 1.939596e-05, 1.939599e-05, 1.939597e-05, 1.939602e-05, 
    1.939601e-05, 1.939602e-05, 1.939603e-05, 1.939598e-05, 1.939601e-05, 
    1.939596e-05, 1.939597e-05, 1.939593e-05, 1.939595e-05, 1.939591e-05, 
    1.939589e-05, 1.939587e-05, 1.939585e-05, 1.939602e-05, 1.939603e-05, 
    1.939601e-05, 1.9396e-05, 1.939599e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939596e-05, 1.939595e-05, 1.939596e-05, 1.939595e-05, 
    1.939601e-05, 1.939598e-05, 1.939603e-05, 1.939601e-05, 1.9396e-05, 
    1.939601e-05, 1.939598e-05, 1.939598e-05, 1.939595e-05, 1.939597e-05, 
    1.939589e-05, 1.939593e-05, 1.939584e-05, 1.939586e-05, 1.939603e-05, 
    1.939602e-05, 1.939599e-05, 1.939601e-05, 1.939597e-05, 1.939596e-05, 
    1.939595e-05, 1.939594e-05, 1.939594e-05, 1.939594e-05, 1.939595e-05, 
    1.939594e-05, 1.939597e-05, 1.939595e-05, 1.9396e-05, 1.939599e-05, 
    1.939599e-05, 1.939599e-05, 1.939598e-05, 1.939596e-05, 1.939596e-05, 
    1.939596e-05, 1.939594e-05, 1.939597e-05, 1.939589e-05, 1.939594e-05, 
    1.939601e-05, 1.9396e-05, 1.939599e-05, 1.9396e-05, 1.939596e-05, 
    1.939597e-05, 1.939594e-05, 1.939595e-05, 1.939593e-05, 1.939594e-05, 
    1.939594e-05, 1.939595e-05, 1.939596e-05, 1.939597e-05, 1.939599e-05, 
    1.9396e-05, 1.9396e-05, 1.939598e-05, 1.939596e-05, 1.939594e-05, 
    1.939595e-05, 1.939593e-05, 1.939597e-05, 1.939595e-05, 1.939596e-05, 
    1.939594e-05, 1.939598e-05, 1.939595e-05, 1.939599e-05, 1.939599e-05, 
    1.939597e-05, 1.939595e-05, 1.939595e-05, 1.939594e-05, 1.939595e-05, 
    1.939596e-05, 1.939596e-05, 1.939597e-05, 1.939598e-05, 1.939599e-05, 
    1.939599e-05, 1.939599e-05, 1.939598e-05, 1.939596e-05, 1.939595e-05, 
    1.939593e-05, 1.939592e-05, 1.93959e-05, 1.939592e-05, 1.939589e-05, 
    1.939591e-05, 1.939587e-05, 1.939595e-05, 1.939591e-05, 1.939597e-05, 
    1.939597e-05, 1.939596e-05, 1.939593e-05, 1.939594e-05, 1.939593e-05, 
    1.939596e-05, 1.939598e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 
    1.939599e-05, 1.939598e-05, 1.939598e-05, 1.939596e-05, 1.939597e-05, 
    1.939594e-05, 1.939593e-05, 1.939589e-05, 1.939587e-05, 1.939585e-05, 
    1.939584e-05, 1.939584e-05, 1.939584e-05 ;

 LITR2C_TO_SOIL1C =
  1.196551e-13, 1.199785e-13, 1.199157e-13, 1.201763e-13, 1.200318e-13, 
    1.202024e-13, 1.197207e-13, 1.199913e-13, 1.198186e-13, 1.196843e-13, 
    1.206813e-13, 1.201879e-13, 1.211933e-13, 1.208792e-13, 1.216676e-13, 
    1.211444e-13, 1.21773e-13, 1.216526e-13, 1.220151e-13, 1.219113e-13, 
    1.223742e-13, 1.22063e-13, 1.226139e-13, 1.222999e-13, 1.22349e-13, 
    1.220527e-13, 1.202874e-13, 1.206199e-13, 1.202676e-13, 1.203151e-13, 
    1.202938e-13, 1.200347e-13, 1.19904e-13, 1.196304e-13, 1.196801e-13, 
    1.198811e-13, 1.203364e-13, 1.20182e-13, 1.205712e-13, 1.205624e-13, 
    1.20995e-13, 1.208e-13, 1.215263e-13, 1.213201e-13, 1.219156e-13, 
    1.21766e-13, 1.219086e-13, 1.218654e-13, 1.219092e-13, 1.216896e-13, 
    1.217837e-13, 1.215905e-13, 1.208366e-13, 1.210583e-13, 1.203964e-13, 
    1.199976e-13, 1.197326e-13, 1.195443e-13, 1.19571e-13, 1.196217e-13, 
    1.198823e-13, 1.201272e-13, 1.203137e-13, 1.204384e-13, 1.205611e-13, 
    1.209323e-13, 1.211287e-13, 1.215679e-13, 1.214888e-13, 1.216229e-13, 
    1.217511e-13, 1.21966e-13, 1.219307e-13, 1.220253e-13, 1.216194e-13, 
    1.218892e-13, 1.214437e-13, 1.215656e-13, 1.205942e-13, 1.202237e-13, 
    1.200658e-13, 1.199277e-13, 1.195914e-13, 1.198237e-13, 1.197321e-13, 
    1.1995e-13, 1.200883e-13, 1.200199e-13, 1.204418e-13, 1.202778e-13, 
    1.211403e-13, 1.207691e-13, 1.217361e-13, 1.21505e-13, 1.217915e-13, 
    1.216454e-13, 1.218957e-13, 1.216704e-13, 1.220606e-13, 1.221454e-13, 
    1.220874e-13, 1.223102e-13, 1.216579e-13, 1.219086e-13, 1.20018e-13, 
    1.200291e-13, 1.200811e-13, 1.198525e-13, 1.198386e-13, 1.19629e-13, 
    1.198155e-13, 1.198948e-13, 1.200963e-13, 1.202153e-13, 1.203285e-13, 
    1.205771e-13, 1.208544e-13, 1.212419e-13, 1.2152e-13, 1.217063e-13, 
    1.215921e-13, 1.216929e-13, 1.215802e-13, 1.215274e-13, 1.221136e-13, 
    1.217846e-13, 1.222782e-13, 1.222509e-13, 1.220276e-13, 1.222539e-13, 
    1.20037e-13, 1.199728e-13, 1.197497e-13, 1.199243e-13, 1.196062e-13, 
    1.197843e-13, 1.198866e-13, 1.202812e-13, 1.203679e-13, 1.204482e-13, 
    1.206067e-13, 1.2081e-13, 1.211663e-13, 1.214761e-13, 1.217585e-13, 
    1.217379e-13, 1.217451e-13, 1.218082e-13, 1.21652e-13, 1.218338e-13, 
    1.218643e-13, 1.217846e-13, 1.222472e-13, 1.221151e-13, 1.222503e-13, 
    1.221643e-13, 1.199936e-13, 1.201016e-13, 1.200433e-13, 1.20153e-13, 
    1.200757e-13, 1.204192e-13, 1.205221e-13, 1.210033e-13, 1.20806e-13, 
    1.211201e-13, 1.20838e-13, 1.208879e-13, 1.211302e-13, 1.208532e-13, 
    1.214589e-13, 1.210483e-13, 1.218106e-13, 1.214009e-13, 1.218363e-13, 
    1.217573e-13, 1.218881e-13, 1.220051e-13, 1.221522e-13, 1.224235e-13, 
    1.223607e-13, 1.225875e-13, 1.202626e-13, 1.204025e-13, 1.203902e-13, 
    1.205367e-13, 1.206449e-13, 1.208793e-13, 1.212549e-13, 1.211138e-13, 
    1.213729e-13, 1.214249e-13, 1.210312e-13, 1.212729e-13, 1.204962e-13, 
    1.206217e-13, 1.20547e-13, 1.202736e-13, 1.211462e-13, 1.206987e-13, 
    1.215246e-13, 1.212826e-13, 1.219884e-13, 1.216375e-13, 1.223262e-13, 
    1.226199e-13, 1.228963e-13, 1.232186e-13, 1.204789e-13, 1.203839e-13, 
    1.205541e-13, 1.207893e-13, 1.210075e-13, 1.212973e-13, 1.21327e-13, 
    1.213812e-13, 1.215218e-13, 1.216398e-13, 1.213983e-13, 1.216694e-13, 
    1.206507e-13, 1.211851e-13, 1.203479e-13, 1.206001e-13, 1.207755e-13, 
    1.206986e-13, 1.210976e-13, 1.211916e-13, 1.21573e-13, 1.213759e-13, 
    1.225473e-13, 1.220297e-13, 1.234639e-13, 1.230639e-13, 1.203506e-13, 
    1.204786e-13, 1.209235e-13, 1.207119e-13, 1.213167e-13, 1.214654e-13, 
    1.215862e-13, 1.217405e-13, 1.217572e-13, 1.218486e-13, 1.216988e-13, 
    1.218427e-13, 1.21298e-13, 1.215415e-13, 1.208727e-13, 1.210356e-13, 
    1.209607e-13, 1.208785e-13, 1.211322e-13, 1.214021e-13, 1.21408e-13, 
    1.214945e-13, 1.217379e-13, 1.213192e-13, 1.226139e-13, 1.218148e-13, 
    1.206181e-13, 1.208642e-13, 1.208994e-13, 1.208041e-13, 1.214505e-13, 
    1.212164e-13, 1.218464e-13, 1.216763e-13, 1.219549e-13, 1.218165e-13, 
    1.217961e-13, 1.216182e-13, 1.215074e-13, 1.212271e-13, 1.20999e-13, 
    1.208179e-13, 1.208601e-13, 1.210589e-13, 1.214186e-13, 1.217587e-13, 
    1.216842e-13, 1.219338e-13, 1.212729e-13, 1.215501e-13, 1.21443e-13, 
    1.217223e-13, 1.2111e-13, 1.216312e-13, 1.209766e-13, 1.210341e-13, 
    1.212118e-13, 1.215689e-13, 1.21648e-13, 1.217322e-13, 1.216802e-13, 
    1.214278e-13, 1.213864e-13, 1.212075e-13, 1.21158e-13, 1.210215e-13, 
    1.209085e-13, 1.210118e-13, 1.211202e-13, 1.214279e-13, 1.21705e-13, 
    1.220067e-13, 1.220805e-13, 1.224324e-13, 1.221459e-13, 1.226183e-13, 
    1.222165e-13, 1.229118e-13, 1.216615e-13, 1.222049e-13, 1.212199e-13, 
    1.213262e-13, 1.215183e-13, 1.219585e-13, 1.21721e-13, 1.219988e-13, 
    1.213848e-13, 1.210657e-13, 1.209832e-13, 1.208289e-13, 1.209867e-13, 
    1.209739e-13, 1.211247e-13, 1.210763e-13, 1.214382e-13, 1.212438e-13, 
    1.217956e-13, 1.219966e-13, 1.225637e-13, 1.229107e-13, 1.232636e-13, 
    1.234192e-13, 1.234666e-13, 1.234864e-13 ;

 LITR2C_vr =
  0.001107536, 0.001107535, 0.001107535, 0.001107534, 0.001107534, 
    0.001107534, 0.001107535, 0.001107535, 0.001107535, 0.001107536, 
    0.001107532, 0.001107534, 0.00110753, 0.001107531, 0.001107529, 
    0.00110753, 0.001107528, 0.001107529, 0.001107527, 0.001107528, 
    0.001107526, 0.001107527, 0.001107525, 0.001107526, 0.001107526, 
    0.001107527, 0.001107533, 0.001107532, 0.001107534, 0.001107533, 
    0.001107533, 0.001107534, 0.001107535, 0.001107536, 0.001107536, 
    0.001107535, 0.001107533, 0.001107534, 0.001107533, 0.001107533, 
    0.001107531, 0.001107532, 0.001107529, 0.00110753, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107528, 0.001107529, 
    0.001107528, 0.001107529, 0.001107532, 0.001107531, 0.001107533, 
    0.001107535, 0.001107535, 0.001107536, 0.001107536, 0.001107536, 
    0.001107535, 0.001107534, 0.001107533, 0.001107533, 0.001107533, 
    0.001107531, 0.001107531, 0.001107529, 0.001107529, 0.001107529, 
    0.001107528, 0.001107528, 0.001107528, 0.001107527, 0.001107529, 
    0.001107528, 0.001107529, 0.001107529, 0.001107532, 0.001107534, 
    0.001107534, 0.001107535, 0.001107536, 0.001107535, 0.001107535, 
    0.001107535, 0.001107534, 0.001107534, 0.001107533, 0.001107533, 
    0.00110753, 0.001107532, 0.001107528, 0.001107529, 0.001107528, 
    0.001107529, 0.001107528, 0.001107529, 0.001107527, 0.001107527, 
    0.001107527, 0.001107526, 0.001107529, 0.001107528, 0.001107534, 
    0.001107534, 0.001107534, 0.001107535, 0.001107535, 0.001107536, 
    0.001107535, 0.001107535, 0.001107534, 0.001107534, 0.001107533, 
    0.001107532, 0.001107531, 0.00110753, 0.001107529, 0.001107529, 
    0.001107529, 0.001107529, 0.001107529, 0.001107529, 0.001107527, 
    0.001107528, 0.001107526, 0.001107527, 0.001107527, 0.001107527, 
    0.001107534, 0.001107535, 0.001107535, 0.001107535, 0.001107536, 
    0.001107535, 0.001107535, 0.001107533, 0.001107533, 0.001107533, 
    0.001107532, 0.001107532, 0.00110753, 0.001107529, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107529, 0.001107528, 
    0.001107528, 0.001107528, 0.001107527, 0.001107527, 0.001107527, 
    0.001107527, 0.001107535, 0.001107534, 0.001107534, 0.001107534, 
    0.001107534, 0.001107533, 0.001107533, 0.001107531, 0.001107532, 
    0.001107531, 0.001107532, 0.001107531, 0.001107531, 0.001107531, 
    0.001107529, 0.001107531, 0.001107528, 0.00110753, 0.001107528, 
    0.001107528, 0.001107528, 0.001107528, 0.001107527, 0.001107526, 
    0.001107526, 0.001107525, 0.001107534, 0.001107533, 0.001107533, 
    0.001107533, 0.001107532, 0.001107531, 0.00110753, 0.001107531, 
    0.00110753, 0.00110753, 0.001107531, 0.00110753, 0.001107533, 
    0.001107532, 0.001107533, 0.001107533, 0.00110753, 0.001107532, 
    0.001107529, 0.00110753, 0.001107528, 0.001107529, 0.001107526, 
    0.001107525, 0.001107524, 0.001107523, 0.001107533, 0.001107533, 
    0.001107533, 0.001107532, 0.001107531, 0.00110753, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.00110753, 0.001107529, 
    0.001107532, 0.00110753, 0.001107533, 0.001107532, 0.001107532, 
    0.001107532, 0.001107531, 0.00110753, 0.001107529, 0.00110753, 
    0.001107526, 0.001107527, 0.001107522, 0.001107524, 0.001107533, 
    0.001107533, 0.001107531, 0.001107532, 0.00110753, 0.001107529, 
    0.001107529, 0.001107528, 0.001107528, 0.001107528, 0.001107529, 
    0.001107528, 0.00110753, 0.001107529, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.001107531, 0.00110753, 0.00110753, 
    0.001107529, 0.001107528, 0.00110753, 0.001107525, 0.001107528, 
    0.001107532, 0.001107531, 0.001107531, 0.001107532, 0.001107529, 
    0.00110753, 0.001107528, 0.001107529, 0.001107528, 0.001107528, 
    0.001107528, 0.001107529, 0.001107529, 0.00110753, 0.001107531, 
    0.001107532, 0.001107531, 0.001107531, 0.00110753, 0.001107528, 
    0.001107529, 0.001107528, 0.00110753, 0.001107529, 0.001107529, 
    0.001107528, 0.001107531, 0.001107529, 0.001107531, 0.001107531, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107529, 
    0.00110753, 0.00110753, 0.00110753, 0.00110753, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107527, 0.001107525, 0.001107527, 
    0.001107524, 0.001107529, 0.001107527, 0.00110753, 0.00110753, 
    0.001107529, 0.001107528, 0.001107528, 0.001107528, 0.00110753, 
    0.001107531, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.00110753, 0.001107528, 
    0.001107528, 0.001107526, 0.001107524, 0.001107523, 0.001107523, 
    0.001107522, 0.001107522,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684274e-07, 2.684271e-07, 2.684271e-07, 2.684269e-07, 2.68427e-07, 
    2.684269e-07, 2.684273e-07, 2.684271e-07, 2.684272e-07, 2.684273e-07, 
    2.684265e-07, 2.684269e-07, 2.68426e-07, 2.684263e-07, 2.684257e-07, 
    2.684261e-07, 2.684256e-07, 2.684257e-07, 2.684254e-07, 2.684255e-07, 
    2.684251e-07, 2.684253e-07, 2.684249e-07, 2.684251e-07, 2.684251e-07, 
    2.684253e-07, 2.684268e-07, 2.684265e-07, 2.684268e-07, 2.684268e-07, 
    2.684268e-07, 2.68427e-07, 2.684272e-07, 2.684274e-07, 2.684273e-07, 
    2.684272e-07, 2.684268e-07, 2.684269e-07, 2.684266e-07, 2.684266e-07, 
    2.684262e-07, 2.684264e-07, 2.684258e-07, 2.684259e-07, 2.684255e-07, 
    2.684256e-07, 2.684255e-07, 2.684255e-07, 2.684255e-07, 2.684256e-07, 
    2.684256e-07, 2.684257e-07, 2.684264e-07, 2.684262e-07, 2.684267e-07, 
    2.684271e-07, 2.684273e-07, 2.684274e-07, 2.684274e-07, 2.684274e-07, 
    2.684272e-07, 2.68427e-07, 2.684268e-07, 2.684267e-07, 2.684266e-07, 
    2.684263e-07, 2.684261e-07, 2.684257e-07, 2.684258e-07, 2.684257e-07, 
    2.684256e-07, 2.684254e-07, 2.684254e-07, 2.684253e-07, 2.684257e-07, 
    2.684255e-07, 2.684259e-07, 2.684257e-07, 2.684266e-07, 2.684269e-07, 
    2.68427e-07, 2.684271e-07, 2.684274e-07, 2.684272e-07, 2.684273e-07, 
    2.684271e-07, 2.68427e-07, 2.68427e-07, 2.684267e-07, 2.684268e-07, 
    2.684261e-07, 2.684264e-07, 2.684256e-07, 2.684258e-07, 2.684255e-07, 
    2.684257e-07, 2.684255e-07, 2.684257e-07, 2.684253e-07, 2.684253e-07, 
    2.684253e-07, 2.684251e-07, 2.684257e-07, 2.684255e-07, 2.68427e-07, 
    2.68427e-07, 2.68427e-07, 2.684272e-07, 2.684272e-07, 2.684274e-07, 
    2.684272e-07, 2.684272e-07, 2.68427e-07, 2.684269e-07, 2.684268e-07, 
    2.684266e-07, 2.684263e-07, 2.68426e-07, 2.684258e-07, 2.684256e-07, 
    2.684257e-07, 2.684256e-07, 2.684257e-07, 2.684258e-07, 2.684253e-07, 
    2.684256e-07, 2.684251e-07, 2.684252e-07, 2.684253e-07, 2.684252e-07, 
    2.68427e-07, 2.684271e-07, 2.684273e-07, 2.684271e-07, 2.684274e-07, 
    2.684272e-07, 2.684272e-07, 2.684268e-07, 2.684268e-07, 2.684267e-07, 
    2.684266e-07, 2.684264e-07, 2.684261e-07, 2.684258e-07, 2.684256e-07, 
    2.684256e-07, 2.684256e-07, 2.684255e-07, 2.684257e-07, 2.684255e-07, 
    2.684255e-07, 2.684256e-07, 2.684252e-07, 2.684253e-07, 2.684252e-07, 
    2.684252e-07, 2.684271e-07, 2.68427e-07, 2.68427e-07, 2.684269e-07, 
    2.68427e-07, 2.684267e-07, 2.684266e-07, 2.684262e-07, 2.684264e-07, 
    2.684261e-07, 2.684264e-07, 2.684263e-07, 2.684261e-07, 2.684263e-07, 
    2.684258e-07, 2.684262e-07, 2.684255e-07, 2.684259e-07, 2.684255e-07, 
    2.684256e-07, 2.684255e-07, 2.684254e-07, 2.684253e-07, 2.68425e-07, 
    2.684251e-07, 2.684249e-07, 2.684268e-07, 2.684267e-07, 2.684267e-07, 
    2.684266e-07, 2.684265e-07, 2.684263e-07, 2.68426e-07, 2.684261e-07, 
    2.684259e-07, 2.684259e-07, 2.684262e-07, 2.68426e-07, 2.684266e-07, 
    2.684265e-07, 2.684266e-07, 2.684268e-07, 2.684261e-07, 2.684265e-07, 
    2.684258e-07, 2.68426e-07, 2.684254e-07, 2.684257e-07, 2.684251e-07, 
    2.684249e-07, 2.684246e-07, 2.684243e-07, 2.684266e-07, 2.684267e-07, 
    2.684266e-07, 2.684264e-07, 2.684262e-07, 2.68426e-07, 2.684259e-07, 
    2.684259e-07, 2.684258e-07, 2.684257e-07, 2.684259e-07, 2.684257e-07, 
    2.684265e-07, 2.68426e-07, 2.684268e-07, 2.684266e-07, 2.684264e-07, 
    2.684265e-07, 2.684261e-07, 2.68426e-07, 2.684257e-07, 2.684259e-07, 
    2.684249e-07, 2.684253e-07, 2.684241e-07, 2.684245e-07, 2.684268e-07, 
    2.684266e-07, 2.684263e-07, 2.684264e-07, 2.684259e-07, 2.684258e-07, 
    2.684257e-07, 2.684256e-07, 2.684256e-07, 2.684255e-07, 2.684256e-07, 
    2.684255e-07, 2.68426e-07, 2.684258e-07, 2.684263e-07, 2.684262e-07, 
    2.684262e-07, 2.684263e-07, 2.684261e-07, 2.684259e-07, 2.684259e-07, 
    2.684258e-07, 2.684256e-07, 2.684259e-07, 2.684249e-07, 2.684255e-07, 
    2.684265e-07, 2.684263e-07, 2.684263e-07, 2.684264e-07, 2.684258e-07, 
    2.68426e-07, 2.684255e-07, 2.684257e-07, 2.684254e-07, 2.684255e-07, 
    2.684255e-07, 2.684257e-07, 2.684258e-07, 2.68426e-07, 2.684262e-07, 
    2.684264e-07, 2.684263e-07, 2.684262e-07, 2.684259e-07, 2.684256e-07, 
    2.684257e-07, 2.684254e-07, 2.68426e-07, 2.684258e-07, 2.684259e-07, 
    2.684256e-07, 2.684261e-07, 2.684257e-07, 2.684262e-07, 2.684262e-07, 
    2.68426e-07, 2.684257e-07, 2.684257e-07, 2.684256e-07, 2.684257e-07, 
    2.684259e-07, 2.684259e-07, 2.68426e-07, 2.684261e-07, 2.684262e-07, 
    2.684263e-07, 2.684262e-07, 2.684261e-07, 2.684259e-07, 2.684256e-07, 
    2.684254e-07, 2.684253e-07, 2.68425e-07, 2.684253e-07, 2.684249e-07, 
    2.684252e-07, 2.684246e-07, 2.684257e-07, 2.684252e-07, 2.68426e-07, 
    2.684259e-07, 2.684258e-07, 2.684254e-07, 2.684256e-07, 2.684254e-07, 
    2.684259e-07, 2.684262e-07, 2.684262e-07, 2.684264e-07, 2.684262e-07, 
    2.684262e-07, 2.684261e-07, 2.684262e-07, 2.684259e-07, 2.68426e-07, 
    2.684255e-07, 2.684254e-07, 2.684249e-07, 2.684246e-07, 2.684243e-07, 
    2.684242e-07, 2.684241e-07, 2.684241e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  5.146902e-26, 1.862688e-25, 1.495052e-25, -8.333079e-26, 1.54407e-25, 
    -8.578169e-26, -8.578169e-26, 4.65672e-26, -9.068351e-26, -4.142031e-25, 
    -6.372354e-26, 6.127264e-26, -3.676358e-26, 2.205815e-26, 1.004871e-25, 
    2.867559e-25, 1.151926e-25, -1.54407e-25, -1.81367e-25, -4.901811e-27, 
    -2.279342e-25, -1.838179e-25, -1.004871e-25, -2.695996e-26, 5.882173e-26, 
    -1.446034e-25, -9.803622e-26, -2.08327e-25, -2.32836e-25, 2.450905e-26, 
    -1.372507e-25, -2.009742e-25, 1.495052e-25, -2.941087e-26, -6.617445e-26, 
    2.475414e-25, -1.323489e-25, -1.666616e-25, 2.941087e-26, -4.043994e-25, 
    8.82326e-26, -3.725376e-25, -7.107626e-26, 1.470543e-26, 4.65672e-26, 
    -1.862688e-25, -7.352717e-27, -1.225453e-26, 5.391992e-26, -1.593089e-25, 
    5.882173e-26, -1.200944e-25, 2.107779e-25, 2.769523e-25, -1.838179e-25, 
    -1.960724e-26, -5.637083e-26, -3.431268e-26, 1.225453e-25, 9.313441e-26, 
    9.313441e-26, -3.676358e-26, -1.004871e-25, 1.764652e-25, 1.053889e-25, 
    1.127417e-25, -9.313441e-26, 1.323489e-25, -2.843051e-25, 1.176435e-25, 
    -5.882173e-26, -3.11265e-25, 1.691125e-25, 2.034252e-25, -1.274471e-25, 
    6.862535e-26, 0, -1.372507e-25, -1.960724e-25, -1.078398e-25, 
    -1.887197e-25, -3.137159e-25, -1.960724e-26, -9.558531e-26, 
    -1.372507e-25, 4.901811e-27, -5.637083e-26, 1.691125e-25, 1.56858e-25, 
    1.004871e-25, -1.421525e-25, 2.205815e-26, -7.107626e-26, 1.176435e-25, 
    -1.225453e-26, 7.352717e-26, -9.068351e-26, -1.372507e-25, -1.54407e-25, 
    5.637083e-26, 1.274471e-25, -1.397016e-25, 2.450906e-27, 2.745014e-25, 
    -7.107626e-26, -1.593089e-25, -1.053889e-25, 1.740143e-25, 7.352717e-27, 
    1.102908e-25, -2.205815e-26, -1.519561e-25, 5.391992e-26, 5.146902e-26, 
    1.470543e-26, -1.81367e-25, 2.034252e-25, 6.617445e-26, 1.176435e-25, 
    3.431268e-26, -5.146902e-26, -7.352717e-26, -1.200944e-25, 1.936215e-25, 
    9.803622e-27, 1.691125e-25, -9.068351e-26, -9.558531e-26, -1.960724e-26, 
    3.921449e-26, 5.391992e-26, -1.495052e-25, 1.446034e-25, 1.715634e-25, 
    6.127264e-26, 1.519561e-25, -1.446034e-25, -9.803622e-26, -1.960724e-25, 
    -2.941087e-26, 7.107626e-26, -8.333079e-26, -2.230324e-25, -2.450905e-26, 
    6.372354e-26, -1.372507e-25, 9.068351e-26, 4.41163e-26, -3.431268e-25, 
    3.921449e-26, 2.548942e-25, 7.597807e-26, 1.911706e-25, 3.676358e-26, 
    -1.666616e-25, -1.887197e-25, -2.695996e-26, 9.558531e-26, 9.803622e-26, 
    7.107626e-26, -7.842898e-26, -1.470543e-25, 6.127264e-26, -1.960724e-26, 
    -3.921449e-26, 2.230324e-25, -5.146902e-26, -7.107626e-26, -9.803622e-26, 
    -1.617598e-25, -4.901811e-26, 7.107626e-26, 9.068351e-26, -1.470543e-25, 
    3.676358e-26, 3.676358e-26, 1.470543e-25, -1.470543e-26, -2.132288e-25, 
    5.882173e-26, -1.617598e-25, -3.186177e-26, -1.397016e-25, 3.431268e-26, 
    6.127264e-26, -1.495052e-25, 8.087988e-26, -7.597807e-26, -4.65672e-26, 
    -6.862535e-26, 3.676358e-26, 1.985233e-25, -5.146902e-26, -2.450905e-26, 
    -5.146902e-26, -1.715634e-25, -7.597807e-26, -2.058761e-25, 7.352717e-26, 
    6.372354e-26, 2.205815e-26, -1.691125e-25, -1.617598e-25, 8.087988e-26, 
    1.397016e-25, -2.450906e-27, -2.941087e-26, 2.450906e-27, -6.617445e-26, 
    2.720505e-25, 2.671487e-25, -1.446034e-25, -7.352717e-27, 2.695996e-25, 
    -4.901811e-26, -1.274471e-25, -1.470543e-26, 2.941087e-26, -2.524433e-25, 
    6.127264e-26, -1.789161e-25, -2.279342e-25, 7.352717e-26, 2.745014e-25, 
    -8.578169e-26, -3.186177e-26, -5.146902e-26, 6.127264e-26, -2.205815e-26, 
    8.087988e-26, -2.205815e-26, 2.181306e-25, -4.65672e-26, -1.102908e-25, 
    -2.941087e-26, -1.02938e-25, -1.249962e-25, 3.186177e-26, -7.352717e-27, 
    -6.617445e-26, -1.078398e-25, -3.186177e-26, 1.323489e-25, -1.176435e-25, 
    1.54407e-25, 8.333079e-26, -2.475414e-25, 0, 8.578169e-26, -2.573451e-25, 
    1.715634e-26, 1.495052e-25, -6.862535e-26, -2.745014e-25, 1.102908e-25, 
    2.450905e-26, 6.127264e-26, -5.146902e-26, 1.176435e-25, 7.352717e-26, 
    1.004871e-25, 6.127264e-26, 1.225453e-26, 8.333079e-26, 8.333079e-26, 
    8.333079e-26, -4.65672e-26, -9.558531e-26, -4.65672e-26, 1.54407e-25, 
    -9.803622e-27, -4.901811e-27, -1.789161e-25, -1.470543e-25, 
    -4.901811e-27, -1.421525e-25, -3.186177e-26, -6.862535e-26, 3.676358e-26, 
    -1.911706e-25, 8.82326e-26, -2.720505e-25, 2.646978e-25, -1.642107e-25, 
    -4.41163e-26, -4.65672e-26, -1.887197e-25, -1.397016e-25, -1.004871e-25, 
    -2.401887e-25, 6.862535e-26, 7.107626e-26, -2.303851e-25, 1.960724e-26, 
    -8.333079e-26, -1.078398e-25, 3.431268e-26, 1.936215e-25, 7.597807e-26, 
    -1.151926e-25, -7.107626e-26, -6.127264e-26, 4.65672e-26, -1.54407e-25, 
    -1.200944e-25, -1.764652e-25, 1.81367e-25, 4.901811e-27, -2.548942e-25, 
    -1.715634e-26, -5.146902e-26, 1.764652e-25, 1.053889e-25, -7.352717e-26, 
    1.789161e-25, 1.249962e-25, -1.56858e-25, -5.637083e-26, 6.617445e-26, 
    1.495052e-25, 9.068351e-26, -1.715634e-26, 1.56858e-25, -2.205815e-26, 
    4.166539e-26, 2.450906e-27, -9.558531e-26, 2.941087e-26, -2.009742e-25, 
    -4.901811e-26, 9.803622e-26, 1.053889e-25, 3.186177e-26, 1.078398e-25, 
    -1.004871e-25, -9.803622e-26, -7.352717e-26, -1.102908e-25,
  2.67626e-32, 2.676257e-32, 2.676258e-32, 2.676255e-32, 2.676257e-32, 
    2.676255e-32, 2.676259e-32, 2.676257e-32, 2.676258e-32, 2.676259e-32, 
    2.676251e-32, 2.676255e-32, 2.676247e-32, 2.676249e-32, 2.676243e-32, 
    2.676247e-32, 2.676242e-32, 2.676243e-32, 2.67624e-32, 2.676241e-32, 
    2.676237e-32, 2.676239e-32, 2.676235e-32, 2.676237e-32, 2.676237e-32, 
    2.676239e-32, 2.676254e-32, 2.676252e-32, 2.676255e-32, 2.676254e-32, 
    2.676254e-32, 2.676257e-32, 2.676258e-32, 2.67626e-32, 2.676259e-32, 
    2.676258e-32, 2.676254e-32, 2.676255e-32, 2.676252e-32, 2.676252e-32, 
    2.676248e-32, 2.67625e-32, 2.676244e-32, 2.676246e-32, 2.676241e-32, 
    2.676242e-32, 2.676241e-32, 2.676241e-32, 2.676241e-32, 2.676242e-32, 
    2.676242e-32, 2.676243e-32, 2.67625e-32, 2.676248e-32, 2.676254e-32, 
    2.676257e-32, 2.676259e-32, 2.676261e-32, 2.676261e-32, 2.67626e-32, 
    2.676258e-32, 2.676256e-32, 2.676254e-32, 2.676253e-32, 2.676252e-32, 
    2.676249e-32, 2.676247e-32, 2.676244e-32, 2.676244e-32, 2.676243e-32, 
    2.676242e-32, 2.67624e-32, 2.67624e-32, 2.67624e-32, 2.676243e-32, 
    2.676241e-32, 2.676244e-32, 2.676244e-32, 2.676252e-32, 2.676255e-32, 
    2.676256e-32, 2.676257e-32, 2.67626e-32, 2.676258e-32, 2.676259e-32, 
    2.676257e-32, 2.676256e-32, 2.676257e-32, 2.676253e-32, 2.676254e-32, 
    2.676247e-32, 2.67625e-32, 2.676242e-32, 2.676244e-32, 2.676242e-32, 
    2.676243e-32, 2.676241e-32, 2.676243e-32, 2.676239e-32, 2.676239e-32, 
    2.676239e-32, 2.676237e-32, 2.676243e-32, 2.676241e-32, 2.676257e-32, 
    2.676257e-32, 2.676256e-32, 2.676258e-32, 2.676258e-32, 2.67626e-32, 
    2.676259e-32, 2.676258e-32, 2.676256e-32, 2.676255e-32, 2.676254e-32, 
    2.676252e-32, 2.67625e-32, 2.676246e-32, 2.676244e-32, 2.676242e-32, 
    2.676243e-32, 2.676242e-32, 2.676244e-32, 2.676244e-32, 2.676239e-32, 
    2.676242e-32, 2.676237e-32, 2.676238e-32, 2.67624e-32, 2.676238e-32, 
    2.676257e-32, 2.676257e-32, 2.676259e-32, 2.676257e-32, 2.67626e-32, 
    2.676259e-32, 2.676258e-32, 2.676254e-32, 2.676254e-32, 2.676253e-32, 
    2.676252e-32, 2.67625e-32, 2.676247e-32, 2.676244e-32, 2.676242e-32, 
    2.676242e-32, 2.676242e-32, 2.676242e-32, 2.676243e-32, 2.676241e-32, 
    2.676241e-32, 2.676242e-32, 2.676238e-32, 2.676239e-32, 2.676238e-32, 
    2.676239e-32, 2.676257e-32, 2.676256e-32, 2.676257e-32, 2.676256e-32, 
    2.676256e-32, 2.676253e-32, 2.676252e-32, 2.676248e-32, 2.67625e-32, 
    2.676247e-32, 2.67625e-32, 2.676249e-32, 2.676247e-32, 2.67625e-32, 
    2.676244e-32, 2.676248e-32, 2.676242e-32, 2.676245e-32, 2.676241e-32, 
    2.676242e-32, 2.676241e-32, 2.67624e-32, 2.676239e-32, 2.676236e-32, 
    2.676237e-32, 2.676235e-32, 2.676255e-32, 2.676254e-32, 2.676254e-32, 
    2.676252e-32, 2.676252e-32, 2.676249e-32, 2.676246e-32, 2.676247e-32, 
    2.676245e-32, 2.676245e-32, 2.676248e-32, 2.676246e-32, 2.676253e-32, 
    2.676252e-32, 2.676252e-32, 2.676254e-32, 2.676247e-32, 2.676251e-32, 
    2.676244e-32, 2.676246e-32, 2.67624e-32, 2.676243e-32, 2.676237e-32, 
    2.676234e-32, 2.676232e-32, 2.676229e-32, 2.676253e-32, 2.676254e-32, 
    2.676252e-32, 2.67625e-32, 2.676248e-32, 2.676246e-32, 2.676246e-32, 
    2.676245e-32, 2.676244e-32, 2.676243e-32, 2.676245e-32, 2.676243e-32, 
    2.676251e-32, 2.676247e-32, 2.676254e-32, 2.676252e-32, 2.67625e-32, 
    2.676251e-32, 2.676248e-32, 2.676247e-32, 2.676244e-32, 2.676245e-32, 
    2.676235e-32, 2.67624e-32, 2.676227e-32, 2.676231e-32, 2.676254e-32, 
    2.676253e-32, 2.676249e-32, 2.676251e-32, 2.676246e-32, 2.676244e-32, 
    2.676243e-32, 2.676242e-32, 2.676242e-32, 2.676241e-32, 2.676242e-32, 
    2.676241e-32, 2.676246e-32, 2.676244e-32, 2.676249e-32, 2.676248e-32, 
    2.676249e-32, 2.676249e-32, 2.676247e-32, 2.676245e-32, 2.676245e-32, 
    2.676244e-32, 2.676242e-32, 2.676246e-32, 2.676235e-32, 2.676242e-32, 
    2.676252e-32, 2.676249e-32, 2.676249e-32, 2.67625e-32, 2.676244e-32, 
    2.676247e-32, 2.676241e-32, 2.676243e-32, 2.67624e-32, 2.676242e-32, 
    2.676242e-32, 2.676243e-32, 2.676244e-32, 2.676247e-32, 2.676248e-32, 
    2.67625e-32, 2.676249e-32, 2.676248e-32, 2.676245e-32, 2.676242e-32, 
    2.676243e-32, 2.67624e-32, 2.676246e-32, 2.676244e-32, 2.676245e-32, 
    2.676242e-32, 2.676247e-32, 2.676243e-32, 2.676249e-32, 2.676248e-32, 
    2.676247e-32, 2.676244e-32, 2.676243e-32, 2.676242e-32, 2.676243e-32, 
    2.676245e-32, 2.676245e-32, 2.676247e-32, 2.676247e-32, 2.676248e-32, 
    2.676249e-32, 2.676248e-32, 2.676247e-32, 2.676245e-32, 2.676242e-32, 
    2.67624e-32, 2.676239e-32, 2.676236e-32, 2.676239e-32, 2.676235e-32, 
    2.676238e-32, 2.676232e-32, 2.676243e-32, 2.676238e-32, 2.676247e-32, 
    2.676246e-32, 2.676244e-32, 2.67624e-32, 2.676242e-32, 2.67624e-32, 
    2.676245e-32, 2.676248e-32, 2.676249e-32, 2.67625e-32, 2.676249e-32, 
    2.676249e-32, 2.676247e-32, 2.676248e-32, 2.676245e-32, 2.676246e-32, 
    2.676242e-32, 2.67624e-32, 2.676235e-32, 2.676232e-32, 2.676229e-32, 
    2.676228e-32, 2.676227e-32, 2.676227e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.311877e-15, 3.320829e-15, 3.31909e-15, 3.326303e-15, 3.322303e-15, 
    3.327025e-15, 3.313693e-15, 3.321183e-15, 3.316403e-15, 3.312684e-15, 
    3.340281e-15, 3.326625e-15, 3.354452e-15, 3.345759e-15, 3.367581e-15, 
    3.353098e-15, 3.370498e-15, 3.367166e-15, 3.377198e-15, 3.374326e-15, 
    3.387137e-15, 3.378523e-15, 3.393773e-15, 3.385082e-15, 3.386441e-15, 
    3.378238e-15, 3.329378e-15, 3.338581e-15, 3.328831e-15, 3.330145e-15, 
    3.329556e-15, 3.322385e-15, 3.318767e-15, 3.311194e-15, 3.31257e-15, 
    3.318133e-15, 3.330735e-15, 3.326461e-15, 3.337233e-15, 3.33699e-15, 
    3.348965e-15, 3.343568e-15, 3.363669e-15, 3.357962e-15, 3.374445e-15, 
    3.370303e-15, 3.37425e-15, 3.373054e-15, 3.374266e-15, 3.36819e-15, 
    3.370794e-15, 3.365445e-15, 3.344578e-15, 3.350716e-15, 3.332396e-15, 
    3.321356e-15, 3.314022e-15, 3.308811e-15, 3.309548e-15, 3.310952e-15, 
    3.318166e-15, 3.324945e-15, 3.330106e-15, 3.333557e-15, 3.336955e-15, 
    3.347228e-15, 3.352665e-15, 3.364822e-15, 3.362631e-15, 3.366343e-15, 
    3.369891e-15, 3.37584e-15, 3.374862e-15, 3.377481e-15, 3.366247e-15, 
    3.373714e-15, 3.361383e-15, 3.364757e-15, 3.33787e-15, 3.327615e-15, 
    3.323244e-15, 3.319424e-15, 3.310114e-15, 3.316544e-15, 3.31401e-15, 
    3.320039e-15, 3.323867e-15, 3.321974e-15, 3.333651e-15, 3.329113e-15, 
    3.352987e-15, 3.342712e-15, 3.369477e-15, 3.363081e-15, 3.37101e-15, 
    3.366965e-15, 3.373893e-15, 3.367659e-15, 3.378457e-15, 3.380805e-15, 
    3.3792e-15, 3.385366e-15, 3.367313e-15, 3.37425e-15, 3.321921e-15, 
    3.322229e-15, 3.323668e-15, 3.317342e-15, 3.316955e-15, 3.311156e-15, 
    3.316317e-15, 3.318513e-15, 3.324089e-15, 3.327384e-15, 3.330516e-15, 
    3.337397e-15, 3.345074e-15, 3.355798e-15, 3.363496e-15, 3.368651e-15, 
    3.365491e-15, 3.368281e-15, 3.365162e-15, 3.3637e-15, 3.379924e-15, 
    3.370817e-15, 3.384479e-15, 3.383724e-15, 3.377543e-15, 3.383809e-15, 
    3.322446e-15, 3.32067e-15, 3.314496e-15, 3.319328e-15, 3.310524e-15, 
    3.315452e-15, 3.318284e-15, 3.329206e-15, 3.331606e-15, 3.333828e-15, 
    3.338216e-15, 3.343844e-15, 3.353706e-15, 3.362279e-15, 3.370098e-15, 
    3.369525e-15, 3.369727e-15, 3.371471e-15, 3.367148e-15, 3.372181e-15, 
    3.373025e-15, 3.370817e-15, 3.383623e-15, 3.379967e-15, 3.383708e-15, 
    3.381328e-15, 3.321248e-15, 3.324237e-15, 3.322622e-15, 3.325658e-15, 
    3.323518e-15, 3.333027e-15, 3.335875e-15, 3.349194e-15, 3.343733e-15, 
    3.352425e-15, 3.344617e-15, 3.346001e-15, 3.352705e-15, 3.34504e-15, 
    3.361805e-15, 3.350439e-15, 3.371539e-15, 3.3602e-15, 3.372249e-15, 
    3.370064e-15, 3.373682e-15, 3.376921e-15, 3.380994e-15, 3.388503e-15, 
    3.386765e-15, 3.393042e-15, 3.328692e-15, 3.332564e-15, 3.332225e-15, 
    3.336277e-15, 3.339272e-15, 3.345762e-15, 3.356158e-15, 3.352251e-15, 
    3.359425e-15, 3.360863e-15, 3.349965e-15, 3.356657e-15, 3.335156e-15, 
    3.338632e-15, 3.336564e-15, 3.328996e-15, 3.353149e-15, 3.340762e-15, 
    3.363623e-15, 3.356923e-15, 3.376459e-15, 3.366748e-15, 3.385808e-15, 
    3.393937e-15, 3.401588e-15, 3.410509e-15, 3.334679e-15, 3.332048e-15, 
    3.336759e-15, 3.34327e-15, 3.349311e-15, 3.357332e-15, 3.358153e-15, 
    3.359654e-15, 3.363543e-15, 3.366811e-15, 3.360127e-15, 3.36763e-15, 
    3.339435e-15, 3.354224e-15, 3.331052e-15, 3.338034e-15, 3.342887e-15, 
    3.34076e-15, 3.351805e-15, 3.354405e-15, 3.364962e-15, 3.359507e-15, 
    3.39193e-15, 3.377602e-15, 3.4173e-15, 3.406227e-15, 3.331129e-15, 
    3.334671e-15, 3.346984e-15, 3.341128e-15, 3.357868e-15, 3.361983e-15, 
    3.365327e-15, 3.369598e-15, 3.37006e-15, 3.372589e-15, 3.368444e-15, 
    3.372426e-15, 3.357349e-15, 3.36409e-15, 3.345579e-15, 3.350088e-15, 
    3.348015e-15, 3.345739e-15, 3.352761e-15, 3.360232e-15, 3.360394e-15, 
    3.362788e-15, 3.369525e-15, 3.357936e-15, 3.393772e-15, 3.371656e-15, 
    3.338531e-15, 3.345343e-15, 3.346318e-15, 3.34368e-15, 3.36157e-15, 
    3.355092e-15, 3.372528e-15, 3.36782e-15, 3.375533e-15, 3.371701e-15, 
    3.371137e-15, 3.366213e-15, 3.363145e-15, 3.355389e-15, 3.349073e-15, 
    3.344063e-15, 3.345229e-15, 3.350731e-15, 3.36069e-15, 3.370101e-15, 
    3.36804e-15, 3.374947e-15, 3.356655e-15, 3.364329e-15, 3.361363e-15, 
    3.369095e-15, 3.352147e-15, 3.366573e-15, 3.348454e-15, 3.350045e-15, 
    3.354964e-15, 3.364848e-15, 3.367037e-15, 3.369369e-15, 3.36793e-15, 
    3.360943e-15, 3.359799e-15, 3.354845e-15, 3.353475e-15, 3.349699e-15, 
    3.346569e-15, 3.349428e-15, 3.352428e-15, 3.360947e-15, 3.368614e-15, 
    3.376966e-15, 3.37901e-15, 3.388747e-15, 3.380818e-15, 3.393895e-15, 
    3.382773e-15, 3.402018e-15, 3.367413e-15, 3.382451e-15, 3.355188e-15, 
    3.358131e-15, 3.363447e-15, 3.375632e-15, 3.369059e-15, 3.376747e-15, 
    3.359754e-15, 3.35092e-15, 3.348636e-15, 3.344367e-15, 3.348733e-15, 
    3.348378e-15, 3.352554e-15, 3.351213e-15, 3.361229e-15, 3.355851e-15, 
    3.371122e-15, 3.376687e-15, 3.392383e-15, 3.401987e-15, 3.411756e-15, 
    3.416062e-15, 3.417373e-15, 3.417921e-15 ;

 LITR2N_vr =
  1.532748e-05, 1.532746e-05, 1.532747e-05, 1.532745e-05, 1.532746e-05, 
    1.532745e-05, 1.532748e-05, 1.532746e-05, 1.532747e-05, 1.532748e-05, 
    1.532743e-05, 1.532745e-05, 1.53274e-05, 1.532742e-05, 1.532738e-05, 
    1.532741e-05, 1.532738e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532735e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 1.532735e-05, 
    1.532736e-05, 1.532745e-05, 1.532743e-05, 1.532745e-05, 1.532745e-05, 
    1.532745e-05, 1.532746e-05, 1.532747e-05, 1.532748e-05, 1.532748e-05, 
    1.532747e-05, 1.532745e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532741e-05, 1.532742e-05, 1.532739e-05, 1.53274e-05, 1.532737e-05, 
    1.532738e-05, 1.532737e-05, 1.532737e-05, 1.532737e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532742e-05, 1.532741e-05, 1.532744e-05, 
    1.532746e-05, 1.532748e-05, 1.532749e-05, 1.532748e-05, 1.532748e-05, 
    1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532738e-05, 
    1.532737e-05, 1.532739e-05, 1.532739e-05, 1.532743e-05, 1.532745e-05, 
    1.532746e-05, 1.532747e-05, 1.532748e-05, 1.532747e-05, 1.532748e-05, 
    1.532747e-05, 1.532746e-05, 1.532746e-05, 1.532744e-05, 1.532745e-05, 
    1.532741e-05, 1.532742e-05, 1.532738e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532738e-05, 1.532736e-05, 1.532736e-05, 
    1.532736e-05, 1.532735e-05, 1.532738e-05, 1.532737e-05, 1.532746e-05, 
    1.532746e-05, 1.532746e-05, 1.532747e-05, 1.532747e-05, 1.532748e-05, 
    1.532747e-05, 1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532745e-05, 
    1.532743e-05, 1.532742e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532739e-05, 1.532739e-05, 1.532736e-05, 
    1.532738e-05, 1.532735e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532746e-05, 1.532746e-05, 1.532747e-05, 1.532747e-05, 1.532748e-05, 
    1.532747e-05, 1.532747e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532743e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532738e-05, 1.532738e-05, 1.532737e-05, 
    1.532737e-05, 1.532738e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532736e-05, 1.532746e-05, 1.532746e-05, 1.532746e-05, 1.532746e-05, 
    1.532746e-05, 1.532744e-05, 1.532744e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532739e-05, 1.532741e-05, 1.532738e-05, 1.53274e-05, 1.532737e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532736e-05, 1.532734e-05, 
    1.532735e-05, 1.532734e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532743e-05, 1.532742e-05, 1.53274e-05, 1.532741e-05, 
    1.53274e-05, 1.532739e-05, 1.532741e-05, 1.53274e-05, 1.532744e-05, 
    1.532743e-05, 1.532744e-05, 1.532745e-05, 1.532741e-05, 1.532743e-05, 
    1.532739e-05, 1.53274e-05, 1.532737e-05, 1.532738e-05, 1.532735e-05, 
    1.532734e-05, 1.532732e-05, 1.532731e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532739e-05, 1.532738e-05, 1.53274e-05, 1.532738e-05, 
    1.532743e-05, 1.53274e-05, 1.532744e-05, 1.532743e-05, 1.532742e-05, 
    1.532743e-05, 1.532741e-05, 1.53274e-05, 1.532739e-05, 1.53274e-05, 
    1.532734e-05, 1.532736e-05, 1.53273e-05, 1.532731e-05, 1.532744e-05, 
    1.532744e-05, 1.532742e-05, 1.532743e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.532738e-05, 1.532737e-05, 1.532738e-05, 
    1.532737e-05, 1.53274e-05, 1.532739e-05, 1.532742e-05, 1.532741e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.53274e-05, 1.532734e-05, 1.532738e-05, 
    1.532743e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532739e-05, 
    1.53274e-05, 1.532737e-05, 1.532738e-05, 1.532737e-05, 1.532737e-05, 
    1.532738e-05, 1.532738e-05, 1.532739e-05, 1.53274e-05, 1.532741e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.53274e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532741e-05, 1.532738e-05, 1.532742e-05, 1.532741e-05, 
    1.53274e-05, 1.532739e-05, 1.532738e-05, 1.532738e-05, 1.532738e-05, 
    1.532739e-05, 1.53274e-05, 1.53274e-05, 1.532741e-05, 1.532741e-05, 
    1.532742e-05, 1.532741e-05, 1.532741e-05, 1.532739e-05, 1.532738e-05, 
    1.532736e-05, 1.532736e-05, 1.532734e-05, 1.532736e-05, 1.532734e-05, 
    1.532736e-05, 1.532732e-05, 1.532738e-05, 1.532736e-05, 1.53274e-05, 
    1.53274e-05, 1.532739e-05, 1.532737e-05, 1.532738e-05, 1.532737e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 
    1.532742e-05, 1.532741e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 
    1.532738e-05, 1.532737e-05, 1.532734e-05, 1.532732e-05, 1.53273e-05, 
    1.53273e-05, 1.53273e-05, 1.532729e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.196551e-13, 1.199785e-13, 1.199157e-13, 1.201763e-13, 1.200318e-13, 
    1.202024e-13, 1.197207e-13, 1.199913e-13, 1.198186e-13, 1.196843e-13, 
    1.206813e-13, 1.201879e-13, 1.211933e-13, 1.208792e-13, 1.216676e-13, 
    1.211444e-13, 1.21773e-13, 1.216526e-13, 1.220151e-13, 1.219113e-13, 
    1.223742e-13, 1.22063e-13, 1.226139e-13, 1.222999e-13, 1.22349e-13, 
    1.220527e-13, 1.202874e-13, 1.206199e-13, 1.202676e-13, 1.203151e-13, 
    1.202938e-13, 1.200347e-13, 1.19904e-13, 1.196304e-13, 1.196801e-13, 
    1.198811e-13, 1.203364e-13, 1.20182e-13, 1.205712e-13, 1.205624e-13, 
    1.20995e-13, 1.208e-13, 1.215263e-13, 1.213201e-13, 1.219156e-13, 
    1.21766e-13, 1.219086e-13, 1.218654e-13, 1.219092e-13, 1.216896e-13, 
    1.217837e-13, 1.215905e-13, 1.208366e-13, 1.210583e-13, 1.203964e-13, 
    1.199976e-13, 1.197326e-13, 1.195443e-13, 1.19571e-13, 1.196217e-13, 
    1.198823e-13, 1.201272e-13, 1.203137e-13, 1.204384e-13, 1.205611e-13, 
    1.209323e-13, 1.211287e-13, 1.215679e-13, 1.214888e-13, 1.216229e-13, 
    1.217511e-13, 1.21966e-13, 1.219307e-13, 1.220253e-13, 1.216194e-13, 
    1.218892e-13, 1.214437e-13, 1.215656e-13, 1.205942e-13, 1.202237e-13, 
    1.200658e-13, 1.199277e-13, 1.195914e-13, 1.198237e-13, 1.197321e-13, 
    1.1995e-13, 1.200883e-13, 1.200199e-13, 1.204418e-13, 1.202778e-13, 
    1.211403e-13, 1.207691e-13, 1.217361e-13, 1.21505e-13, 1.217915e-13, 
    1.216454e-13, 1.218957e-13, 1.216704e-13, 1.220606e-13, 1.221454e-13, 
    1.220874e-13, 1.223102e-13, 1.216579e-13, 1.219086e-13, 1.20018e-13, 
    1.200291e-13, 1.200811e-13, 1.198525e-13, 1.198386e-13, 1.19629e-13, 
    1.198155e-13, 1.198948e-13, 1.200963e-13, 1.202153e-13, 1.203285e-13, 
    1.205771e-13, 1.208544e-13, 1.212419e-13, 1.2152e-13, 1.217063e-13, 
    1.215921e-13, 1.216929e-13, 1.215802e-13, 1.215274e-13, 1.221136e-13, 
    1.217846e-13, 1.222782e-13, 1.222509e-13, 1.220276e-13, 1.222539e-13, 
    1.20037e-13, 1.199728e-13, 1.197497e-13, 1.199243e-13, 1.196062e-13, 
    1.197843e-13, 1.198866e-13, 1.202812e-13, 1.203679e-13, 1.204482e-13, 
    1.206067e-13, 1.2081e-13, 1.211663e-13, 1.214761e-13, 1.217585e-13, 
    1.217379e-13, 1.217451e-13, 1.218082e-13, 1.21652e-13, 1.218338e-13, 
    1.218643e-13, 1.217846e-13, 1.222472e-13, 1.221151e-13, 1.222503e-13, 
    1.221643e-13, 1.199936e-13, 1.201016e-13, 1.200433e-13, 1.20153e-13, 
    1.200757e-13, 1.204192e-13, 1.205221e-13, 1.210033e-13, 1.20806e-13, 
    1.211201e-13, 1.20838e-13, 1.208879e-13, 1.211302e-13, 1.208532e-13, 
    1.214589e-13, 1.210483e-13, 1.218106e-13, 1.214009e-13, 1.218363e-13, 
    1.217573e-13, 1.218881e-13, 1.220051e-13, 1.221522e-13, 1.224235e-13, 
    1.223607e-13, 1.225875e-13, 1.202626e-13, 1.204025e-13, 1.203902e-13, 
    1.205367e-13, 1.206449e-13, 1.208793e-13, 1.212549e-13, 1.211138e-13, 
    1.213729e-13, 1.214249e-13, 1.210312e-13, 1.212729e-13, 1.204962e-13, 
    1.206217e-13, 1.20547e-13, 1.202736e-13, 1.211462e-13, 1.206987e-13, 
    1.215246e-13, 1.212826e-13, 1.219884e-13, 1.216375e-13, 1.223262e-13, 
    1.226199e-13, 1.228963e-13, 1.232186e-13, 1.204789e-13, 1.203839e-13, 
    1.205541e-13, 1.207893e-13, 1.210075e-13, 1.212973e-13, 1.21327e-13, 
    1.213812e-13, 1.215218e-13, 1.216398e-13, 1.213983e-13, 1.216694e-13, 
    1.206507e-13, 1.211851e-13, 1.203479e-13, 1.206001e-13, 1.207755e-13, 
    1.206986e-13, 1.210976e-13, 1.211916e-13, 1.21573e-13, 1.213759e-13, 
    1.225473e-13, 1.220297e-13, 1.234639e-13, 1.230639e-13, 1.203506e-13, 
    1.204786e-13, 1.209235e-13, 1.207119e-13, 1.213167e-13, 1.214654e-13, 
    1.215862e-13, 1.217405e-13, 1.217572e-13, 1.218486e-13, 1.216988e-13, 
    1.218427e-13, 1.21298e-13, 1.215415e-13, 1.208727e-13, 1.210356e-13, 
    1.209607e-13, 1.208785e-13, 1.211322e-13, 1.214021e-13, 1.21408e-13, 
    1.214945e-13, 1.217379e-13, 1.213192e-13, 1.226139e-13, 1.218148e-13, 
    1.206181e-13, 1.208642e-13, 1.208994e-13, 1.208041e-13, 1.214505e-13, 
    1.212164e-13, 1.218464e-13, 1.216763e-13, 1.219549e-13, 1.218165e-13, 
    1.217961e-13, 1.216182e-13, 1.215074e-13, 1.212271e-13, 1.20999e-13, 
    1.208179e-13, 1.208601e-13, 1.210589e-13, 1.214186e-13, 1.217587e-13, 
    1.216842e-13, 1.219338e-13, 1.212729e-13, 1.215501e-13, 1.21443e-13, 
    1.217223e-13, 1.2111e-13, 1.216312e-13, 1.209766e-13, 1.210341e-13, 
    1.212118e-13, 1.215689e-13, 1.21648e-13, 1.217322e-13, 1.216802e-13, 
    1.214278e-13, 1.213864e-13, 1.212075e-13, 1.21158e-13, 1.210215e-13, 
    1.209085e-13, 1.210118e-13, 1.211202e-13, 1.214279e-13, 1.21705e-13, 
    1.220067e-13, 1.220805e-13, 1.224324e-13, 1.221459e-13, 1.226183e-13, 
    1.222165e-13, 1.229118e-13, 1.216615e-13, 1.222049e-13, 1.212199e-13, 
    1.213262e-13, 1.215183e-13, 1.219585e-13, 1.21721e-13, 1.219988e-13, 
    1.213848e-13, 1.210657e-13, 1.209832e-13, 1.208289e-13, 1.209867e-13, 
    1.209739e-13, 1.211247e-13, 1.210763e-13, 1.214382e-13, 1.212438e-13, 
    1.217956e-13, 1.219966e-13, 1.225637e-13, 1.229107e-13, 1.232636e-13, 
    1.234192e-13, 1.234666e-13, 1.234864e-13 ;

 LITR3C =
  9.698032e-06, 9.698022e-06, 9.698025e-06, 9.698017e-06, 9.698021e-06, 
    9.698016e-06, 9.69803e-06, 9.698022e-06, 9.698027e-06, 9.698031e-06, 
    9.698001e-06, 9.698016e-06, 9.697986e-06, 9.697995e-06, 9.697971e-06, 
    9.697987e-06, 9.697967e-06, 9.697971e-06, 9.69796e-06, 9.697964e-06, 
    9.697949e-06, 9.697958e-06, 9.697942e-06, 9.697952e-06, 9.69795e-06, 
    9.697959e-06, 9.698013e-06, 9.698003e-06, 9.698014e-06, 9.698012e-06, 
    9.698013e-06, 9.698021e-06, 9.698025e-06, 9.698033e-06, 9.698031e-06, 
    9.698026e-06, 9.698011e-06, 9.698017e-06, 9.698005e-06, 9.698005e-06, 
    9.697991e-06, 9.697997e-06, 9.697976e-06, 9.697981e-06, 9.697963e-06, 
    9.697967e-06, 9.697964e-06, 9.697965e-06, 9.697964e-06, 9.69797e-06, 
    9.697967e-06, 9.697973e-06, 9.697997e-06, 9.697989e-06, 9.698009e-06, 
    9.698022e-06, 9.69803e-06, 9.698036e-06, 9.698035e-06, 9.698033e-06, 
    9.698026e-06, 9.698017e-06, 9.698012e-06, 9.698008e-06, 9.698005e-06, 
    9.697993e-06, 9.697987e-06, 9.697974e-06, 9.697977e-06, 9.697972e-06, 
    9.697968e-06, 9.697962e-06, 9.697963e-06, 9.69796e-06, 9.697972e-06, 
    9.697964e-06, 9.697977e-06, 9.697974e-06, 9.698004e-06, 9.698015e-06, 
    9.69802e-06, 9.698024e-06, 9.698034e-06, 9.698027e-06, 9.69803e-06, 
    9.698023e-06, 9.698019e-06, 9.698021e-06, 9.698008e-06, 9.698013e-06, 
    9.697987e-06, 9.697998e-06, 9.697968e-06, 9.697976e-06, 9.697967e-06, 
    9.697972e-06, 9.697964e-06, 9.697971e-06, 9.697959e-06, 9.697957e-06, 
    9.697958e-06, 9.697951e-06, 9.697971e-06, 9.697964e-06, 9.698021e-06, 
    9.698021e-06, 9.698019e-06, 9.698027e-06, 9.698027e-06, 9.698033e-06, 
    9.698027e-06, 9.698025e-06, 9.698019e-06, 9.698016e-06, 9.698012e-06, 
    9.698004e-06, 9.697996e-06, 9.697984e-06, 9.697976e-06, 9.697969e-06, 
    9.697973e-06, 9.69797e-06, 9.697974e-06, 9.697975e-06, 9.697957e-06, 
    9.697967e-06, 9.697952e-06, 9.697953e-06, 9.69796e-06, 9.697953e-06, 
    9.698021e-06, 9.698023e-06, 9.698029e-06, 9.698024e-06, 9.698034e-06, 
    9.698028e-06, 9.698026e-06, 9.698013e-06, 9.69801e-06, 9.698008e-06, 
    9.698003e-06, 9.697997e-06, 9.697987e-06, 9.697977e-06, 9.697968e-06, 
    9.697968e-06, 9.697968e-06, 9.697967e-06, 9.697971e-06, 9.697966e-06, 
    9.697965e-06, 9.697967e-06, 9.697953e-06, 9.697957e-06, 9.697953e-06, 
    9.697956e-06, 9.698022e-06, 9.698018e-06, 9.69802e-06, 9.698017e-06, 
    9.698019e-06, 9.698009e-06, 9.698006e-06, 9.697991e-06, 9.697997e-06, 
    9.697987e-06, 9.697997e-06, 9.697995e-06, 9.697987e-06, 9.697996e-06, 
    9.697977e-06, 9.69799e-06, 9.697967e-06, 9.697979e-06, 9.697966e-06, 
    9.697968e-06, 9.697964e-06, 9.69796e-06, 9.697956e-06, 9.697947e-06, 
    9.697949e-06, 9.697943e-06, 9.698014e-06, 9.698009e-06, 9.69801e-06, 
    9.698006e-06, 9.698002e-06, 9.697995e-06, 9.697984e-06, 9.697987e-06, 
    9.69798e-06, 9.697978e-06, 9.69799e-06, 9.697983e-06, 9.698007e-06, 
    9.698003e-06, 9.698005e-06, 9.698014e-06, 9.697987e-06, 9.698e-06, 
    9.697976e-06, 9.697983e-06, 9.697961e-06, 9.697972e-06, 9.697951e-06, 
    9.697942e-06, 9.697934e-06, 9.697924e-06, 9.698007e-06, 9.69801e-06, 
    9.698005e-06, 9.697997e-06, 9.697991e-06, 9.697982e-06, 9.697981e-06, 
    9.697979e-06, 9.697976e-06, 9.697972e-06, 9.697979e-06, 9.697971e-06, 
    9.698002e-06, 9.697986e-06, 9.698011e-06, 9.698004e-06, 9.697998e-06, 
    9.698e-06, 9.697988e-06, 9.697986e-06, 9.697974e-06, 9.69798e-06, 
    9.697944e-06, 9.69796e-06, 9.697916e-06, 9.697928e-06, 9.698011e-06, 
    9.698007e-06, 9.697994e-06, 9.698e-06, 9.697982e-06, 9.697977e-06, 
    9.697973e-06, 9.697968e-06, 9.697968e-06, 9.697966e-06, 9.69797e-06, 
    9.697966e-06, 9.697982e-06, 9.697975e-06, 9.697995e-06, 9.69799e-06, 
    9.697992e-06, 9.697995e-06, 9.697987e-06, 9.697979e-06, 9.697978e-06, 
    9.697977e-06, 9.697968e-06, 9.697981e-06, 9.697942e-06, 9.697967e-06, 
    9.698003e-06, 9.697996e-06, 9.697995e-06, 9.697997e-06, 9.697977e-06, 
    9.697985e-06, 9.697966e-06, 9.69797e-06, 9.697962e-06, 9.697967e-06, 
    9.697967e-06, 9.697972e-06, 9.697976e-06, 9.697985e-06, 9.697991e-06, 
    9.697997e-06, 9.697996e-06, 9.697989e-06, 9.697978e-06, 9.697968e-06, 
    9.69797e-06, 9.697963e-06, 9.697983e-06, 9.697975e-06, 9.697977e-06, 
    9.697969e-06, 9.697987e-06, 9.697972e-06, 9.697992e-06, 9.69799e-06, 
    9.697985e-06, 9.697974e-06, 9.697971e-06, 9.697969e-06, 9.69797e-06, 
    9.697978e-06, 9.697979e-06, 9.697985e-06, 9.697987e-06, 9.69799e-06, 
    9.697994e-06, 9.697991e-06, 9.697987e-06, 9.697978e-06, 9.69797e-06, 
    9.69796e-06, 9.697958e-06, 9.697947e-06, 9.697957e-06, 9.697942e-06, 
    9.697954e-06, 9.697933e-06, 9.697971e-06, 9.697955e-06, 9.697985e-06, 
    9.697981e-06, 9.697976e-06, 9.697962e-06, 9.697969e-06, 9.697961e-06, 
    9.697979e-06, 9.697989e-06, 9.697992e-06, 9.697997e-06, 9.697992e-06, 
    9.697992e-06, 9.697987e-06, 9.697989e-06, 9.697977e-06, 9.697984e-06, 
    9.697967e-06, 9.697961e-06, 9.697944e-06, 9.697933e-06, 9.697922e-06, 
    9.697917e-06, 9.697916e-06, 9.697916e-06 ;

 LITR3C_TO_SOIL2C =
  5.982752e-14, 5.998923e-14, 5.995782e-14, 6.008813e-14, 6.001588e-14, 
    6.010117e-14, 5.986034e-14, 5.999564e-14, 5.990929e-14, 5.984211e-14, 
    6.034062e-14, 6.009395e-14, 6.059662e-14, 6.043959e-14, 6.08338e-14, 
    6.057217e-14, 6.08865e-14, 6.08263e-14, 6.100752e-14, 6.095563e-14, 
    6.118706e-14, 6.103146e-14, 6.130695e-14, 6.114994e-14, 6.117449e-14, 
    6.102632e-14, 6.014367e-14, 6.030992e-14, 6.01338e-14, 6.015752e-14, 
    6.014689e-14, 6.001735e-14, 5.9952e-14, 5.981518e-14, 5.984005e-14, 
    5.994054e-14, 6.016819e-14, 6.009098e-14, 6.028558e-14, 6.028119e-14, 
    6.04975e-14, 6.040001e-14, 6.076313e-14, 6.066003e-14, 6.09578e-14, 
    6.088297e-14, 6.095427e-14, 6.093266e-14, 6.095456e-14, 6.08448e-14, 
    6.089183e-14, 6.079522e-14, 6.041826e-14, 6.052914e-14, 6.019818e-14, 
    5.999876e-14, 5.986627e-14, 5.977215e-14, 5.978546e-14, 5.981082e-14, 
    5.994113e-14, 6.006359e-14, 6.015683e-14, 6.021916e-14, 6.028056e-14, 
    6.046612e-14, 6.056434e-14, 6.078394e-14, 6.074438e-14, 6.081144e-14, 
    6.087552e-14, 6.0983e-14, 6.096532e-14, 6.101264e-14, 6.080969e-14, 
    6.094459e-14, 6.072183e-14, 6.078279e-14, 6.029708e-14, 6.011182e-14, 
    6.003287e-14, 5.996385e-14, 5.979569e-14, 5.991183e-14, 5.986605e-14, 
    5.997497e-14, 6.004412e-14, 6.000993e-14, 6.022086e-14, 6.013889e-14, 
    6.057016e-14, 6.038455e-14, 6.086805e-14, 6.07525e-14, 6.089573e-14, 
    6.082267e-14, 6.094782e-14, 6.083519e-14, 6.103026e-14, 6.107267e-14, 
    6.104369e-14, 6.115507e-14, 6.082895e-14, 6.095426e-14, 6.000896e-14, 
    6.001454e-14, 6.004053e-14, 5.992625e-14, 5.991926e-14, 5.98145e-14, 
    5.990773e-14, 5.994741e-14, 6.004814e-14, 6.010766e-14, 6.016423e-14, 
    6.028853e-14, 6.042721e-14, 6.062095e-14, 6.076e-14, 6.085312e-14, 
    6.079603e-14, 6.084644e-14, 6.079009e-14, 6.076368e-14, 6.105677e-14, 
    6.089226e-14, 6.113905e-14, 6.112541e-14, 6.101376e-14, 6.112695e-14, 
    6.001846e-14, 5.998637e-14, 5.987484e-14, 5.996213e-14, 5.980309e-14, 
    5.989211e-14, 5.994326e-14, 6.014057e-14, 6.018392e-14, 6.022406e-14, 
    6.030334e-14, 6.0405e-14, 6.058316e-14, 6.073802e-14, 6.087925e-14, 
    6.086891e-14, 6.087255e-14, 6.090407e-14, 6.082596e-14, 6.091689e-14, 
    6.093213e-14, 6.089226e-14, 6.112358e-14, 6.105754e-14, 6.112512e-14, 
    6.108213e-14, 5.99968e-14, 6.00508e-14, 6.002162e-14, 6.007648e-14, 
    6.003782e-14, 6.020959e-14, 6.026105e-14, 6.050164e-14, 6.040299e-14, 
    6.056001e-14, 6.041896e-14, 6.044395e-14, 6.056506e-14, 6.04266e-14, 
    6.072945e-14, 6.052413e-14, 6.090529e-14, 6.070045e-14, 6.091812e-14, 
    6.087864e-14, 6.094401e-14, 6.100251e-14, 6.10761e-14, 6.121174e-14, 
    6.118035e-14, 6.129373e-14, 6.013128e-14, 6.020123e-14, 6.019511e-14, 
    6.026831e-14, 6.032241e-14, 6.043965e-14, 6.062745e-14, 6.055687e-14, 
    6.068645e-14, 6.071244e-14, 6.051558e-14, 6.063645e-14, 6.024806e-14, 
    6.031085e-14, 6.027349e-14, 6.013678e-14, 6.057309e-14, 6.034932e-14, 
    6.076229e-14, 6.064127e-14, 6.099416e-14, 6.081875e-14, 6.116306e-14, 
    6.13099e-14, 6.144811e-14, 6.160927e-14, 6.023943e-14, 6.019191e-14, 
    6.027702e-14, 6.039463e-14, 6.050375e-14, 6.064865e-14, 6.066348e-14, 
    6.06906e-14, 6.076086e-14, 6.081989e-14, 6.069915e-14, 6.083469e-14, 
    6.032535e-14, 6.059252e-14, 6.017391e-14, 6.030005e-14, 6.038771e-14, 
    6.03493e-14, 6.05488e-14, 6.059577e-14, 6.078648e-14, 6.068795e-14, 
    6.127365e-14, 6.101482e-14, 6.173194e-14, 6.153191e-14, 6.017529e-14, 
    6.023928e-14, 6.046172e-14, 6.035593e-14, 6.065833e-14, 6.073266e-14, 
    6.079308e-14, 6.087023e-14, 6.087858e-14, 6.092426e-14, 6.084938e-14, 
    6.092132e-14, 6.064896e-14, 6.077074e-14, 6.043635e-14, 6.051779e-14, 
    6.048034e-14, 6.043922e-14, 6.056607e-14, 6.070104e-14, 6.070397e-14, 
    6.074721e-14, 6.086891e-14, 6.065956e-14, 6.130693e-14, 6.09074e-14, 
    6.030902e-14, 6.043207e-14, 6.044969e-14, 6.040203e-14, 6.072521e-14, 
    6.060819e-14, 6.092316e-14, 6.083811e-14, 6.097744e-14, 6.090822e-14, 
    6.089803e-14, 6.080908e-14, 6.075365e-14, 6.061355e-14, 6.049946e-14, 
    6.040895e-14, 6.043001e-14, 6.052941e-14, 6.07093e-14, 6.087931e-14, 
    6.084208e-14, 6.096686e-14, 6.063643e-14, 6.077505e-14, 6.072147e-14, 
    6.086115e-14, 6.055498e-14, 6.081559e-14, 6.048827e-14, 6.051701e-14, 
    6.060586e-14, 6.078442e-14, 6.082397e-14, 6.086609e-14, 6.084011e-14, 
    6.071388e-14, 6.069321e-14, 6.060372e-14, 6.057898e-14, 6.051076e-14, 
    6.045423e-14, 6.050587e-14, 6.056006e-14, 6.071395e-14, 6.085246e-14, 
    6.100333e-14, 6.104025e-14, 6.121616e-14, 6.107291e-14, 6.130914e-14, 
    6.110823e-14, 6.145589e-14, 6.083075e-14, 6.110242e-14, 6.060992e-14, 
    6.066308e-14, 6.075911e-14, 6.097923e-14, 6.086049e-14, 6.099937e-14, 
    6.06924e-14, 6.053282e-14, 6.049156e-14, 6.041445e-14, 6.049332e-14, 
    6.048691e-14, 6.056234e-14, 6.053811e-14, 6.071906e-14, 6.062189e-14, 
    6.089776e-14, 6.099828e-14, 6.128183e-14, 6.145533e-14, 6.163179e-14, 
    6.170959e-14, 6.173327e-14, 6.174316e-14 ;

 LITR3C_vr =
  0.0005537677, 0.0005537671, 0.0005537672, 0.0005537667, 0.000553767, 
    0.0005537667, 0.0005537675, 0.0005537671, 0.0005537674, 0.0005537676, 
    0.0005537659, 0.0005537667, 0.000553765, 0.0005537655, 0.0005537642, 
    0.000553765, 0.000553764, 0.0005537642, 0.0005537635, 0.0005537638, 
    0.0005537629, 0.0005537635, 0.0005537625, 0.0005537631, 0.0005537629, 
    0.0005537635, 0.0005537666, 0.000553766, 0.0005537666, 0.0005537665, 
    0.0005537666, 0.000553767, 0.0005537673, 0.0005537677, 0.0005537676, 
    0.0005537673, 0.0005537665, 0.0005537667, 0.0005537661, 0.0005537661, 
    0.0005537653, 0.0005537657, 0.0005537644, 0.0005537648, 0.0005537637, 
    0.000553764, 0.0005537638, 0.0005537638, 0.0005537638, 0.0005537641, 
    0.0005537639, 0.0005537643, 0.0005537656, 0.0005537652, 0.0005537664, 
    0.0005537671, 0.0005537675, 0.0005537678, 0.0005537678, 0.0005537677, 
    0.0005537673, 0.0005537668, 0.0005537665, 0.0005537663, 0.0005537661, 
    0.0005537655, 0.0005537651, 0.0005537643, 0.0005537645, 0.0005537642, 
    0.000553764, 0.0005537636, 0.0005537637, 0.0005537635, 0.0005537642, 
    0.0005537638, 0.0005537646, 0.0005537643, 0.000553766, 0.0005537667, 
    0.000553767, 0.0005537672, 0.0005537678, 0.0005537674, 0.0005537675, 
    0.0005537671, 0.0005537669, 0.000553767, 0.0005537663, 0.0005537666, 
    0.0005537651, 0.0005537657, 0.0005537641, 0.0005537645, 0.0005537639, 
    0.0005537642, 0.0005537638, 0.0005537642, 0.0005537635, 0.0005537634, 
    0.0005537634, 0.0005537631, 0.0005537642, 0.0005537638, 0.000553767, 
    0.000553767, 0.0005537669, 0.0005537673, 0.0005537674, 0.0005537677, 
    0.0005537674, 0.0005537673, 0.0005537669, 0.0005537667, 0.0005537665, 
    0.000553766, 0.0005537656, 0.0005537649, 0.0005537644, 0.0005537641, 
    0.0005537643, 0.0005537641, 0.0005537643, 0.0005537644, 0.0005537634, 
    0.0005537639, 0.0005537631, 0.0005537631, 0.0005537635, 0.0005537631, 
    0.000553767, 0.0005537671, 0.0005537675, 0.0005537672, 0.0005537678, 
    0.0005537674, 0.0005537673, 0.0005537666, 0.0005537664, 0.0005537663, 
    0.000553766, 0.0005537657, 0.000553765, 0.0005537645, 0.000553764, 
    0.0005537641, 0.000553764, 0.0005537639, 0.0005537642, 0.0005537639, 
    0.0005537638, 0.0005537639, 0.0005537631, 0.0005537634, 0.0005537631, 
    0.0005537633, 0.0005537671, 0.0005537669, 0.000553767, 0.0005537668, 
    0.0005537669, 0.0005537663, 0.0005537661, 0.0005537653, 0.0005537657, 
    0.0005537651, 0.0005537656, 0.0005537655, 0.0005537651, 0.0005537656, 
    0.0005537645, 0.0005537652, 0.0005537639, 0.0005537646, 0.0005537639, 
    0.000553764, 0.0005537638, 0.0005537636, 0.0005537633, 0.0005537628, 
    0.0005537629, 0.0005537625, 0.0005537666, 0.0005537664, 0.0005537664, 
    0.0005537661, 0.0005537659, 0.0005537655, 0.0005537649, 0.0005537651, 
    0.0005537647, 0.0005537646, 0.0005537653, 0.0005537649, 0.0005537662, 
    0.000553766, 0.0005537661, 0.0005537666, 0.000553765, 0.0005537659, 
    0.0005537644, 0.0005537648, 0.0005537636, 0.0005537642, 0.000553763, 
    0.0005537625, 0.000553762, 0.0005537614, 0.0005537662, 0.0005537664, 
    0.0005537661, 0.0005537657, 0.0005537653, 0.0005537648, 0.0005537648, 
    0.0005537646, 0.0005537644, 0.0005537642, 0.0005537646, 0.0005537642, 
    0.0005537659, 0.000553765, 0.0005537664, 0.000553766, 0.0005537657, 
    0.0005537659, 0.0005537652, 0.000553765, 0.0005537643, 0.0005537647, 
    0.0005537626, 0.0005537635, 0.000553761, 0.0005537617, 0.0005537664, 
    0.0005537662, 0.0005537655, 0.0005537658, 0.0005537648, 0.0005537645, 
    0.0005537643, 0.0005537641, 0.000553764, 0.0005537638, 0.0005537641, 
    0.0005537639, 0.0005537648, 0.0005537644, 0.0005537656, 0.0005537653, 
    0.0005537654, 0.0005537655, 0.0005537651, 0.0005537646, 0.0005537646, 
    0.0005537645, 0.0005537641, 0.0005537648, 0.0005537625, 0.0005537639, 
    0.000553766, 0.0005537656, 0.0005537655, 0.0005537657, 0.0005537645, 
    0.0005537649, 0.0005537638, 0.0005537642, 0.0005537636, 0.0005537639, 
    0.0005537639, 0.0005537642, 0.0005537645, 0.0005537649, 0.0005537653, 
    0.0005537656, 0.0005537656, 0.0005537652, 0.0005537646, 0.000553764, 
    0.0005537641, 0.0005537637, 0.0005537649, 0.0005537643, 0.0005537646, 
    0.0005537641, 0.0005537652, 0.0005537642, 0.0005537654, 0.0005537653, 
    0.0005537649, 0.0005537643, 0.0005537642, 0.0005537641, 0.0005537641, 
    0.0005537646, 0.0005537646, 0.000553765, 0.000553765, 0.0005537653, 
    0.0005537655, 0.0005537653, 0.0005537651, 0.0005537646, 0.0005537641, 
    0.0005537636, 0.0005537634, 0.0005537628, 0.0005537633, 0.0005537625, 
    0.0005537632, 0.000553762, 0.0005537642, 0.0005537632, 0.0005537649, 
    0.0005537648, 0.0005537644, 0.0005537636, 0.0005537641, 0.0005537636, 
    0.0005537646, 0.0005537652, 0.0005537653, 0.0005537656, 0.0005537653, 
    0.0005537654, 0.0005537651, 0.0005537652, 0.0005537646, 0.0005537649, 
    0.0005537639, 0.0005537636, 0.0005537626, 0.000553762, 0.0005537614, 
    0.0005537611, 0.000553761, 0.000553761,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342137e-07, 1.342135e-07, 1.342136e-07, 1.342135e-07, 1.342135e-07, 
    1.342134e-07, 1.342136e-07, 1.342135e-07, 1.342136e-07, 1.342137e-07, 
    1.342132e-07, 1.342135e-07, 1.34213e-07, 1.342132e-07, 1.342128e-07, 
    1.34213e-07, 1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342127e-07, 
    1.342125e-07, 1.342127e-07, 1.342124e-07, 1.342126e-07, 1.342125e-07, 
    1.342127e-07, 1.342134e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 
    1.342134e-07, 1.342135e-07, 1.342136e-07, 1.342137e-07, 1.342137e-07, 
    1.342136e-07, 1.342134e-07, 1.342135e-07, 1.342133e-07, 1.342133e-07, 
    1.342131e-07, 1.342132e-07, 1.342129e-07, 1.34213e-07, 1.342127e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 1.342128e-07, 
    1.342128e-07, 1.342129e-07, 1.342132e-07, 1.342131e-07, 1.342134e-07, 
    1.342135e-07, 1.342136e-07, 1.342137e-07, 1.342137e-07, 1.342137e-07, 
    1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 1.342128e-07, 
    1.342127e-07, 1.342129e-07, 1.342129e-07, 1.342133e-07, 1.342134e-07, 
    1.342135e-07, 1.342136e-07, 1.342137e-07, 1.342136e-07, 1.342136e-07, 
    1.342136e-07, 1.342135e-07, 1.342135e-07, 1.342133e-07, 1.342134e-07, 
    1.34213e-07, 1.342132e-07, 1.342128e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342125e-07, 1.342128e-07, 1.342127e-07, 1.342135e-07, 
    1.342135e-07, 1.342135e-07, 1.342136e-07, 1.342136e-07, 1.342137e-07, 
    1.342136e-07, 1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342132e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 
    1.342129e-07, 1.342128e-07, 1.342129e-07, 1.342129e-07, 1.342126e-07, 
    1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342135e-07, 1.342135e-07, 1.342136e-07, 1.342136e-07, 1.342137e-07, 
    1.342136e-07, 1.342136e-07, 1.342134e-07, 1.342134e-07, 1.342133e-07, 
    1.342133e-07, 1.342132e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342128e-07, 1.342128e-07, 1.342128e-07, 1.342128e-07, 
    1.342127e-07, 1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 
    1.342126e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 
    1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342129e-07, 1.342131e-07, 1.342128e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342134e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342133e-07, 1.342132e-07, 1.34213e-07, 1.342131e-07, 
    1.342129e-07, 1.342129e-07, 1.342131e-07, 1.34213e-07, 1.342133e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.34213e-07, 1.342132e-07, 
    1.342129e-07, 1.34213e-07, 1.342127e-07, 1.342128e-07, 1.342125e-07, 
    1.342124e-07, 1.342123e-07, 1.342122e-07, 1.342133e-07, 1.342134e-07, 
    1.342133e-07, 1.342132e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 
    1.342129e-07, 1.342129e-07, 1.342128e-07, 1.342129e-07, 1.342128e-07, 
    1.342133e-07, 1.34213e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342124e-07, 1.342127e-07, 1.342121e-07, 1.342122e-07, 1.342134e-07, 
    1.342133e-07, 1.342131e-07, 1.342132e-07, 1.34213e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342128e-07, 
    1.342127e-07, 1.34213e-07, 1.342129e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.34213e-07, 1.342124e-07, 1.342128e-07, 
    1.342133e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342129e-07, 
    1.34213e-07, 1.342127e-07, 1.342128e-07, 1.342127e-07, 1.342128e-07, 
    1.342128e-07, 1.342128e-07, 1.342129e-07, 1.34213e-07, 1.342131e-07, 
    1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342131e-07, 1.342128e-07, 1.342131e-07, 1.342131e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 1.342128e-07, 
    1.342129e-07, 1.342129e-07, 1.34213e-07, 1.34213e-07, 1.342131e-07, 
    1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342128e-07, 
    1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 1.342124e-07, 
    1.342126e-07, 1.342123e-07, 1.342128e-07, 1.342126e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342127e-07, 1.342128e-07, 1.342127e-07, 
    1.342129e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342129e-07, 1.34213e-07, 
    1.342128e-07, 1.342127e-07, 1.342124e-07, 1.342123e-07, 1.342121e-07, 
    1.342121e-07, 1.342121e-07, 1.34212e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  7.720352e-26, -7.597807e-26, 5.024356e-26, -1.225453e-27, -5.024356e-26, 
    9.803622e-26, 8.087988e-26, 9.803622e-26, 1.470543e-26, 8.82326e-26, 
    -1.347998e-26, 8.945805e-26, 7.352717e-26, 5.391992e-26, 4.043994e-26, 
    -3.186177e-26, 6.862535e-26, 4.901811e-26, 7.230172e-26, 7.652491e-42, 
    1.225453e-26, -4.166539e-26, 7.352717e-26, -8.945805e-26, 7.107626e-26, 
    -9.681077e-26, -5.759628e-26, 9.803622e-27, -1.225453e-27, 1.495052e-25, 
    -2.205815e-26, 8.333079e-26, 4.65672e-26, -7.597807e-26, 6.127264e-27, 
    -1.960724e-26, -1.960724e-26, -9.926167e-26, -5.637083e-26, 
    -4.901811e-26, -8.333079e-26, -1.372507e-25, -7.842898e-26, 4.043994e-26, 
    -1.225453e-26, -4.166539e-26, -6.372354e-26, -5.759628e-26, 4.043994e-26, 
    -1.960724e-26, 4.534175e-26, 9.803622e-27, -7.107626e-26, 4.289085e-26, 
    7.652491e-42, -2.08327e-26, 4.534175e-26, -9.558531e-26, -3.308722e-26, 
    -3.553813e-26, -8.087988e-26, -6.98508e-26, 3.798904e-26, 3.676358e-26, 
    -7.597807e-26, -2.32836e-26, -9.068351e-26, -5.269447e-26, -7.652491e-42, 
    3.676358e-27, 1.43378e-25, 8.578169e-26, -2.08327e-26, -6.4949e-26, 
    5.759628e-26, 5.759628e-26, 2.695996e-26, -1.347998e-26, -4.901811e-27, 
    -3.431268e-26, 6.004719e-26, 3.431268e-26, 8.210533e-26, -2.941087e-26, 
    2.32836e-26, -6.862535e-26, -3.063632e-26, -4.779266e-26, 4.901811e-27, 
    -3.798904e-26, -2.132288e-25, -8.210533e-26, 3.676358e-27, -4.901811e-27, 
    1.262216e-25, -1.225453e-27, -4.166539e-26, -4.779266e-26, 9.803622e-26, 
    7.107626e-26, -4.166539e-26, -1.115162e-25, -5.024356e-26, -8.578169e-27, 
    -5.024356e-26, -4.166539e-26, -6.98508e-26, -1.200944e-25, -7.965443e-26, 
    -4.043994e-26, -7.352717e-27, 9.803622e-27, 3.676358e-27, 7.352717e-27, 
    -8.945805e-26, -1.715634e-26, -2.450905e-26, 2.058761e-25, 7.475262e-26, 
    1.225453e-26, 1.053889e-25, 5.024356e-26, -3.676358e-27, 2.205815e-26, 
    6.004719e-26, -1.188689e-25, -2.08327e-26, -9.803622e-27, 8.700715e-26, 
    1.960724e-26, -1.102908e-26, -1.041635e-25, 1.102908e-26, -2.695996e-26, 
    5.024356e-26, -1.127417e-25, -1.335744e-25, -5.024356e-26, -2.941087e-26, 
    3.676358e-26, 1.16418e-25, 1.225453e-26, 8.945805e-26, 4.779266e-26, 
    -7.965443e-26, 5.391992e-26, -1.715634e-26, -3.676358e-27, -3.676358e-27, 
    1.102908e-26, 1.593089e-26, 1.274471e-25, 1.347998e-26, -3.798904e-26, 
    4.166539e-26, -1.225453e-26, 7.230172e-26, -1.838179e-26, -2.695996e-26, 
    4.901811e-26, -5.759628e-26, 2.573451e-26, 4.41163e-26, 1.960724e-26, 
    4.901811e-26, -6.73999e-26, 1.923961e-25, -3.063632e-26, 9.435986e-26, 
    6.4949e-26, 5.269447e-26, -5.146902e-26, 5.391992e-26, -9.558531e-26, 
    2.205815e-26, -6.372354e-26, -1.053889e-25, 1.139671e-25, 2.32836e-26, 
    -2.573451e-26, 2.08327e-26, -1.053889e-25, -1.54407e-25, -9.681077e-26, 
    -2.695996e-26, 6.4949e-26, 3.308722e-26, 4.166539e-26, -5.146902e-26, 
    -9.068351e-26, 9.558531e-26, -2.695996e-26, 4.779266e-26, -5.882173e-26, 
    -4.901811e-27, 1.54407e-25, 4.289085e-26, 5.882173e-26, 7.720352e-26, 
    1.02938e-25, -3.431268e-26, 1.225453e-27, -7.720352e-26, 2.08327e-26, 
    9.926167e-26, 4.534175e-26, -8.82326e-26, 1.249962e-25, -2.818541e-26, 
    -1.347998e-26, -3.676358e-27, 7.230172e-26, 8.087988e-26, 5.391992e-26, 
    -1.090653e-25, 1.311234e-25, 1.593089e-26, -7.352717e-27, -2.818541e-26, 
    -1.262216e-25, -4.41163e-26, 1.960724e-26, -4.65672e-26, -3.798904e-26, 
    -1.115162e-25, -1.225453e-26, 1.200944e-25, -1.225453e-27, 9.190896e-26, 
    -2.941087e-26, 8.578169e-26, 3.921449e-26, 7.352717e-27, 8.82326e-26, 
    3.553813e-26, -1.176435e-25, -7.230172e-26, 7.107626e-26, 1.053889e-25, 
    -1.090653e-25, -1.482798e-25, 2.08327e-26, 6.127264e-27, 6.004719e-26, 
    7.475262e-26, -1.347998e-26, -2.573451e-26, -7.352717e-27, 4.901811e-26, 
    -2.941087e-26, -1.102908e-26, -8.945805e-26, 1.789161e-25, -3.676358e-26, 
    2.818541e-26, 3.308722e-26, 3.186177e-26, -8.210533e-26, 2.695996e-26, 
    -7.352717e-27, 4.779266e-26, -6.372354e-26, -4.779266e-26, 8.455624e-26, 
    1.593089e-26, -4.534175e-26, 1.286725e-25, 5.882173e-26, 7.842898e-26, 
    3.826946e-42, 8.578169e-26, -2.450905e-26, 9.803622e-27, 2.818541e-26, 
    7.965443e-26, -7.352717e-27, -1.617598e-25, -1.335744e-25, -3.676358e-27, 
    4.043994e-26, 1.102908e-26, 6.617445e-26, -1.470543e-26, -1.593089e-25, 
    9.435986e-26, -7.720352e-26, -4.65672e-26, 6.4949e-26, 7.842898e-26, 
    1.593089e-26, 1.470543e-26, 1.311234e-25, 3.431268e-26, 3.676358e-26, 
    2.08327e-26, 4.41163e-26, -4.779266e-26, -5.146902e-26, 3.798904e-26, 
    9.803622e-27, 2.573451e-26, 6.617445e-26, 9.190896e-26, -3.676358e-27, 
    5.759628e-26, 6.617445e-26, 1.347998e-26, -1.446034e-25, -2.08327e-26, 0, 
    8.945805e-26, -9.190896e-26, -7.965443e-26, -5.024356e-26, -3.553813e-26, 
    -8.578169e-27, -6.862535e-26, -8.82326e-26, 1.02938e-25, -3.063632e-26, 
    -3.308722e-26, 1.053889e-25, -2.08327e-26, 8.578169e-27, -7.352717e-27, 
    1.102908e-25, 2.818541e-26, 7.352717e-27, 8.700715e-26, 6.127264e-27, 
    3.063632e-26, 4.901811e-27, 7.230172e-26, 4.043994e-26, 5.637083e-26, 
    7.352717e-26, 1.262216e-25, 2.08327e-26,
  1.33813e-32, 1.338128e-32, 1.338129e-32, 1.338128e-32, 1.338128e-32, 
    1.338128e-32, 1.33813e-32, 1.338128e-32, 1.338129e-32, 1.33813e-32, 
    1.338125e-32, 1.338128e-32, 1.338123e-32, 1.338125e-32, 1.338121e-32, 
    1.338124e-32, 1.338121e-32, 1.338121e-32, 1.33812e-32, 1.33812e-32, 
    1.338118e-32, 1.33812e-32, 1.338117e-32, 1.338119e-32, 1.338118e-32, 
    1.33812e-32, 1.338127e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 
    1.338127e-32, 1.338128e-32, 1.338129e-32, 1.33813e-32, 1.33813e-32, 
    1.338129e-32, 1.338127e-32, 1.338128e-32, 1.338126e-32, 1.338126e-32, 
    1.338124e-32, 1.338125e-32, 1.338122e-32, 1.338123e-32, 1.33812e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338121e-32, 
    1.338121e-32, 1.338122e-32, 1.338125e-32, 1.338124e-32, 1.338127e-32, 
    1.338128e-32, 1.33813e-32, 1.33813e-32, 1.33813e-32, 1.33813e-32, 
    1.338129e-32, 1.338128e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338121e-32, 
    1.33812e-32, 1.338122e-32, 1.338122e-32, 1.338126e-32, 1.338127e-32, 
    1.338128e-32, 1.338129e-32, 1.33813e-32, 1.338129e-32, 1.33813e-32, 
    1.338129e-32, 1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338127e-32, 
    1.338124e-32, 1.338125e-32, 1.338121e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338119e-32, 1.338121e-32, 1.33812e-32, 1.338128e-32, 
    1.338128e-32, 1.338128e-32, 1.338129e-32, 1.338129e-32, 1.33813e-32, 
    1.338129e-32, 1.338129e-32, 1.338128e-32, 1.338128e-32, 1.338127e-32, 
    1.338126e-32, 1.338125e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 
    1.338122e-32, 1.338121e-32, 1.338122e-32, 1.338122e-32, 1.338119e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338128e-32, 1.338129e-32, 1.338129e-32, 1.338129e-32, 1.33813e-32, 
    1.338129e-32, 1.338129e-32, 1.338127e-32, 1.338127e-32, 1.338126e-32, 
    1.338126e-32, 1.338125e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.338121e-32, 1.338121e-32, 1.338121e-32, 1.338121e-32, 
    1.33812e-32, 1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 
    1.338119e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 
    1.338128e-32, 1.338127e-32, 1.338126e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338122e-32, 1.338124e-32, 1.338121e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338127e-32, 1.338127e-32, 1.338127e-32, 
    1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338123e-32, 1.338124e-32, 
    1.338123e-32, 1.338122e-32, 1.338124e-32, 1.338123e-32, 1.338126e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338124e-32, 1.338125e-32, 
    1.338122e-32, 1.338123e-32, 1.33812e-32, 1.338121e-32, 1.338119e-32, 
    1.338117e-32, 1.338116e-32, 1.338115e-32, 1.338126e-32, 1.338127e-32, 
    1.338126e-32, 1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338122e-32, 1.338121e-32, 
    1.338126e-32, 1.338123e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338123e-32, 
    1.338118e-32, 1.33812e-32, 1.338114e-32, 1.338115e-32, 1.338127e-32, 
    1.338126e-32, 1.338124e-32, 1.338125e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338121e-32, 1.33812e-32, 1.338121e-32, 
    1.338121e-32, 1.338123e-32, 1.338122e-32, 1.338125e-32, 1.338124e-32, 
    1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338123e-32, 1.338117e-32, 1.338121e-32, 
    1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338122e-32, 
    1.338123e-32, 1.33812e-32, 1.338121e-32, 1.33812e-32, 1.338121e-32, 
    1.338121e-32, 1.338121e-32, 1.338122e-32, 1.338123e-32, 1.338124e-32, 
    1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.338124e-32, 1.338121e-32, 1.338124e-32, 1.338124e-32, 
    1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 1.338121e-32, 
    1.338122e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 1.338124e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338121e-32, 
    1.33812e-32, 1.33812e-32, 1.338118e-32, 1.338119e-32, 1.338117e-32, 
    1.338119e-32, 1.338116e-32, 1.338121e-32, 1.338119e-32, 1.338123e-32, 
    1.338123e-32, 1.338122e-32, 1.33812e-32, 1.338121e-32, 1.33812e-32, 
    1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 
    1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338116e-32, 1.338114e-32, 
    1.338114e-32, 1.338114e-32, 1.338114e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.655938e-15, 1.660414e-15, 1.659545e-15, 1.663152e-15, 1.661152e-15, 
    1.663512e-15, 1.656847e-15, 1.660591e-15, 1.658202e-15, 1.656342e-15, 
    1.67014e-15, 1.663312e-15, 1.677226e-15, 1.672879e-15, 1.68379e-15, 
    1.676549e-15, 1.685249e-15, 1.683583e-15, 1.688599e-15, 1.687163e-15, 
    1.693568e-15, 1.689262e-15, 1.696887e-15, 1.692541e-15, 1.693221e-15, 
    1.689119e-15, 1.664689e-15, 1.66929e-15, 1.664416e-15, 1.665072e-15, 
    1.664778e-15, 1.661193e-15, 1.659384e-15, 1.655597e-15, 1.656285e-15, 
    1.659066e-15, 1.665367e-15, 1.663231e-15, 1.668617e-15, 1.668495e-15, 
    1.674482e-15, 1.671784e-15, 1.681835e-15, 1.678981e-15, 1.687223e-15, 
    1.685151e-15, 1.687125e-15, 1.686527e-15, 1.687133e-15, 1.684095e-15, 
    1.685397e-15, 1.682723e-15, 1.672289e-15, 1.675358e-15, 1.666198e-15, 
    1.660678e-15, 1.657011e-15, 1.654406e-15, 1.654774e-15, 1.655476e-15, 
    1.659083e-15, 1.662472e-15, 1.665053e-15, 1.666778e-15, 1.668478e-15, 
    1.673614e-15, 1.676332e-15, 1.682411e-15, 1.681316e-15, 1.683171e-15, 
    1.684945e-15, 1.68792e-15, 1.687431e-15, 1.68874e-15, 1.683123e-15, 
    1.686857e-15, 1.680691e-15, 1.682379e-15, 1.668935e-15, 1.663807e-15, 
    1.661622e-15, 1.659712e-15, 1.655057e-15, 1.658272e-15, 1.657005e-15, 
    1.66002e-15, 1.661933e-15, 1.660987e-15, 1.666825e-15, 1.664556e-15, 
    1.676493e-15, 1.671356e-15, 1.684738e-15, 1.681541e-15, 1.685505e-15, 
    1.683483e-15, 1.686946e-15, 1.683829e-15, 1.689228e-15, 1.690402e-15, 
    1.6896e-15, 1.692683e-15, 1.683656e-15, 1.687125e-15, 1.66096e-15, 
    1.661115e-15, 1.661834e-15, 1.658671e-15, 1.658477e-15, 1.655578e-15, 
    1.658158e-15, 1.659257e-15, 1.662045e-15, 1.663692e-15, 1.665258e-15, 
    1.668698e-15, 1.672537e-15, 1.677899e-15, 1.681748e-15, 1.684325e-15, 
    1.682745e-15, 1.68414e-15, 1.682581e-15, 1.68185e-15, 1.689962e-15, 
    1.685409e-15, 1.69224e-15, 1.691862e-15, 1.688772e-15, 1.691905e-15, 
    1.661223e-15, 1.660335e-15, 1.657248e-15, 1.659664e-15, 1.655262e-15, 
    1.657726e-15, 1.659142e-15, 1.664603e-15, 1.665803e-15, 1.666914e-15, 
    1.669108e-15, 1.671922e-15, 1.676853e-15, 1.681139e-15, 1.685049e-15, 
    1.684763e-15, 1.684863e-15, 1.685736e-15, 1.683574e-15, 1.68609e-15, 
    1.686512e-15, 1.685409e-15, 1.691811e-15, 1.689983e-15, 1.691854e-15, 
    1.690664e-15, 1.660624e-15, 1.662118e-15, 1.661311e-15, 1.662829e-15, 
    1.661759e-15, 1.666513e-15, 1.667938e-15, 1.674597e-15, 1.671866e-15, 
    1.676212e-15, 1.672308e-15, 1.673e-15, 1.676352e-15, 1.67252e-15, 
    1.680902e-15, 1.675219e-15, 1.685769e-15, 1.6801e-15, 1.686124e-15, 
    1.685032e-15, 1.686841e-15, 1.68846e-15, 1.690497e-15, 1.694251e-15, 
    1.693383e-15, 1.696521e-15, 1.664346e-15, 1.666282e-15, 1.666112e-15, 
    1.668139e-15, 1.669636e-15, 1.672881e-15, 1.678079e-15, 1.676125e-15, 
    1.679712e-15, 1.680432e-15, 1.674983e-15, 1.678328e-15, 1.667578e-15, 
    1.669316e-15, 1.668282e-15, 1.664498e-15, 1.676575e-15, 1.670381e-15, 
    1.681811e-15, 1.678462e-15, 1.688229e-15, 1.683374e-15, 1.692904e-15, 
    1.696968e-15, 1.700794e-15, 1.705254e-15, 1.667339e-15, 1.666024e-15, 
    1.66838e-15, 1.671635e-15, 1.674655e-15, 1.678666e-15, 1.679076e-15, 
    1.679827e-15, 1.681772e-15, 1.683405e-15, 1.680064e-15, 1.683815e-15, 
    1.669717e-15, 1.677112e-15, 1.665526e-15, 1.669017e-15, 1.671443e-15, 
    1.67038e-15, 1.675902e-15, 1.677202e-15, 1.682481e-15, 1.679754e-15, 
    1.695965e-15, 1.688801e-15, 1.70865e-15, 1.703113e-15, 1.665564e-15, 
    1.667335e-15, 1.673492e-15, 1.670564e-15, 1.678934e-15, 1.680991e-15, 
    1.682663e-15, 1.684799e-15, 1.68503e-15, 1.686294e-15, 1.684222e-15, 
    1.686213e-15, 1.678674e-15, 1.682045e-15, 1.67279e-15, 1.675044e-15, 
    1.674007e-15, 1.672869e-15, 1.67638e-15, 1.680116e-15, 1.680197e-15, 
    1.681394e-15, 1.684762e-15, 1.678968e-15, 1.696886e-15, 1.685828e-15, 
    1.669266e-15, 1.672671e-15, 1.673159e-15, 1.67184e-15, 1.680785e-15, 
    1.677546e-15, 1.686264e-15, 1.68391e-15, 1.687766e-15, 1.68585e-15, 
    1.685568e-15, 1.683106e-15, 1.681572e-15, 1.677694e-15, 1.674537e-15, 
    1.672031e-15, 1.672614e-15, 1.675366e-15, 1.680345e-15, 1.68505e-15, 
    1.68402e-15, 1.687473e-15, 1.678328e-15, 1.682165e-15, 1.680682e-15, 
    1.684547e-15, 1.676073e-15, 1.683287e-15, 1.674227e-15, 1.675022e-15, 
    1.677482e-15, 1.682424e-15, 1.683518e-15, 1.684684e-15, 1.683965e-15, 
    1.680471e-15, 1.679899e-15, 1.677422e-15, 1.676738e-15, 1.674849e-15, 
    1.673285e-15, 1.674714e-15, 1.676214e-15, 1.680473e-15, 1.684307e-15, 
    1.688483e-15, 1.689505e-15, 1.694374e-15, 1.690409e-15, 1.696947e-15, 
    1.691386e-15, 1.701009e-15, 1.683706e-15, 1.691225e-15, 1.677594e-15, 
    1.679065e-15, 1.681723e-15, 1.687816e-15, 1.684529e-15, 1.688373e-15, 
    1.679877e-15, 1.67546e-15, 1.674318e-15, 1.672184e-15, 1.674367e-15, 
    1.674189e-15, 1.676277e-15, 1.675606e-15, 1.680615e-15, 1.677925e-15, 
    1.685561e-15, 1.688343e-15, 1.696191e-15, 1.700994e-15, 1.705878e-15, 
    1.708031e-15, 1.708686e-15, 1.70896e-15 ;

 LITR3N_vr =
  7.66374e-06, 7.663732e-06, 7.663733e-06, 7.663727e-06, 7.663731e-06, 
    7.663726e-06, 7.663738e-06, 7.663732e-06, 7.663735e-06, 7.663739e-06, 
    7.663714e-06, 7.663726e-06, 7.663702e-06, 7.66371e-06, 7.663691e-06, 
    7.663703e-06, 7.663688e-06, 7.663691e-06, 7.663682e-06, 7.663685e-06, 
    7.663673e-06, 7.663682e-06, 7.663668e-06, 7.663675e-06, 7.663674e-06, 
    7.663682e-06, 7.663724e-06, 7.663716e-06, 7.663724e-06, 7.663723e-06, 
    7.663724e-06, 7.66373e-06, 7.663733e-06, 7.66374e-06, 7.663739e-06, 
    7.663734e-06, 7.663722e-06, 7.663727e-06, 7.663717e-06, 7.663717e-06, 
    7.663707e-06, 7.663712e-06, 7.663694e-06, 7.663699e-06, 7.663684e-06, 
    7.663688e-06, 7.663685e-06, 7.663686e-06, 7.663685e-06, 7.66369e-06, 
    7.663688e-06, 7.663692e-06, 7.663711e-06, 7.663705e-06, 7.663722e-06, 
    7.663731e-06, 7.663737e-06, 7.663742e-06, 7.663742e-06, 7.66374e-06, 
    7.663733e-06, 7.663728e-06, 7.663723e-06, 7.663721e-06, 7.663717e-06, 
    7.663709e-06, 7.663703e-06, 7.663693e-06, 7.663695e-06, 7.663692e-06, 
    7.663689e-06, 7.663683e-06, 7.663684e-06, 7.663682e-06, 7.663692e-06, 
    7.663685e-06, 7.663696e-06, 7.663693e-06, 7.663717e-06, 7.663725e-06, 
    7.66373e-06, 7.663733e-06, 7.663741e-06, 7.663735e-06, 7.663737e-06, 
    7.663733e-06, 7.663729e-06, 7.663731e-06, 7.663721e-06, 7.663724e-06, 
    7.663703e-06, 7.663712e-06, 7.663689e-06, 7.663694e-06, 7.663688e-06, 
    7.663692e-06, 7.663685e-06, 7.663691e-06, 7.663682e-06, 7.663679e-06, 
    7.663681e-06, 7.663675e-06, 7.663691e-06, 7.663685e-06, 7.663731e-06, 
    7.663731e-06, 7.663729e-06, 7.663734e-06, 7.663735e-06, 7.66374e-06, 
    7.663735e-06, 7.663733e-06, 7.663729e-06, 7.663726e-06, 7.663723e-06, 
    7.663717e-06, 7.663711e-06, 7.663701e-06, 7.663694e-06, 7.66369e-06, 
    7.663692e-06, 7.66369e-06, 7.663692e-06, 7.663694e-06, 7.66368e-06, 
    7.663688e-06, 7.663676e-06, 7.663677e-06, 7.663682e-06, 7.663676e-06, 
    7.66373e-06, 7.663732e-06, 7.663737e-06, 7.663733e-06, 7.663741e-06, 
    7.663736e-06, 7.663733e-06, 7.663724e-06, 7.663722e-06, 7.66372e-06, 
    7.663716e-06, 7.663712e-06, 7.663702e-06, 7.663695e-06, 7.663689e-06, 
    7.663689e-06, 7.663689e-06, 7.663687e-06, 7.663691e-06, 7.663687e-06, 
    7.663686e-06, 7.663688e-06, 7.663677e-06, 7.66368e-06, 7.663677e-06, 
    7.663679e-06, 7.663732e-06, 7.663729e-06, 7.66373e-06, 7.663727e-06, 
    7.663729e-06, 7.663721e-06, 7.663718e-06, 7.663707e-06, 7.663712e-06, 
    7.663704e-06, 7.663711e-06, 7.66371e-06, 7.663703e-06, 7.663711e-06, 
    7.663696e-06, 7.663706e-06, 7.663687e-06, 7.663697e-06, 7.663687e-06, 
    7.663689e-06, 7.663685e-06, 7.663682e-06, 7.663679e-06, 7.663672e-06, 
    7.663674e-06, 7.663669e-06, 7.663724e-06, 7.663722e-06, 7.663722e-06, 
    7.663718e-06, 7.663715e-06, 7.66371e-06, 7.663701e-06, 7.663704e-06, 
    7.663698e-06, 7.663697e-06, 7.663706e-06, 7.663701e-06, 7.663719e-06, 
    7.663716e-06, 7.663718e-06, 7.663724e-06, 7.663703e-06, 7.663714e-06, 
    7.663694e-06, 7.6637e-06, 7.663683e-06, 7.663692e-06, 7.663675e-06, 
    7.663668e-06, 7.663661e-06, 7.663653e-06, 7.66372e-06, 7.663722e-06, 
    7.663718e-06, 7.663712e-06, 7.663707e-06, 7.6637e-06, 7.663699e-06, 
    7.663698e-06, 7.663694e-06, 7.663692e-06, 7.663697e-06, 7.663691e-06, 
    7.663715e-06, 7.663702e-06, 7.663722e-06, 7.663716e-06, 7.663712e-06, 
    7.663714e-06, 7.663704e-06, 7.663702e-06, 7.663693e-06, 7.663698e-06, 
    7.66367e-06, 7.663682e-06, 7.663647e-06, 7.663657e-06, 7.663722e-06, 
    7.66372e-06, 7.663709e-06, 7.663713e-06, 7.663699e-06, 7.663695e-06, 
    7.663692e-06, 7.663689e-06, 7.663689e-06, 7.663686e-06, 7.66369e-06, 
    7.663686e-06, 7.6637e-06, 7.663693e-06, 7.66371e-06, 7.663706e-06, 
    7.663708e-06, 7.66371e-06, 7.663703e-06, 7.663697e-06, 7.663697e-06, 
    7.663695e-06, 7.663689e-06, 7.663699e-06, 7.663668e-06, 7.663687e-06, 
    7.663716e-06, 7.66371e-06, 7.663709e-06, 7.663712e-06, 7.663696e-06, 
    7.663702e-06, 7.663686e-06, 7.663691e-06, 7.663683e-06, 7.663687e-06, 
    7.663688e-06, 7.663692e-06, 7.663694e-06, 7.663702e-06, 7.663707e-06, 
    7.663712e-06, 7.663711e-06, 7.663705e-06, 7.663697e-06, 7.663689e-06, 
    7.663691e-06, 7.663684e-06, 7.663701e-06, 7.663693e-06, 7.663696e-06, 
    7.66369e-06, 7.663704e-06, 7.663692e-06, 7.663707e-06, 7.663706e-06, 
    7.663702e-06, 7.663693e-06, 7.663692e-06, 7.663689e-06, 7.663691e-06, 
    7.663696e-06, 7.663698e-06, 7.663702e-06, 7.663703e-06, 7.663706e-06, 
    7.663709e-06, 7.663706e-06, 7.663704e-06, 7.663696e-06, 7.66369e-06, 
    7.663682e-06, 7.663681e-06, 7.663672e-06, 7.663679e-06, 7.663668e-06, 
    7.663677e-06, 7.663661e-06, 7.663691e-06, 7.663678e-06, 7.663702e-06, 
    7.663699e-06, 7.663694e-06, 7.663683e-06, 7.66369e-06, 7.663682e-06, 
    7.663698e-06, 7.663705e-06, 7.663707e-06, 7.663711e-06, 7.663707e-06, 
    7.663708e-06, 7.663703e-06, 7.663705e-06, 7.663696e-06, 7.663701e-06, 
    7.663688e-06, 7.663682e-06, 7.663669e-06, 7.663661e-06, 7.663652e-06, 
    7.663649e-06, 7.663647e-06, 7.663647e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.982752e-14, 5.998923e-14, 5.995782e-14, 6.008813e-14, 6.001588e-14, 
    6.010117e-14, 5.986034e-14, 5.999564e-14, 5.990929e-14, 5.984211e-14, 
    6.034062e-14, 6.009395e-14, 6.059662e-14, 6.043959e-14, 6.08338e-14, 
    6.057217e-14, 6.08865e-14, 6.08263e-14, 6.100752e-14, 6.095563e-14, 
    6.118706e-14, 6.103146e-14, 6.130695e-14, 6.114994e-14, 6.117449e-14, 
    6.102632e-14, 6.014367e-14, 6.030992e-14, 6.01338e-14, 6.015752e-14, 
    6.014689e-14, 6.001735e-14, 5.9952e-14, 5.981518e-14, 5.984005e-14, 
    5.994054e-14, 6.016819e-14, 6.009098e-14, 6.028558e-14, 6.028119e-14, 
    6.04975e-14, 6.040001e-14, 6.076313e-14, 6.066003e-14, 6.09578e-14, 
    6.088297e-14, 6.095427e-14, 6.093266e-14, 6.095456e-14, 6.08448e-14, 
    6.089183e-14, 6.079522e-14, 6.041826e-14, 6.052914e-14, 6.019818e-14, 
    5.999876e-14, 5.986627e-14, 5.977215e-14, 5.978546e-14, 5.981082e-14, 
    5.994113e-14, 6.006359e-14, 6.015683e-14, 6.021916e-14, 6.028056e-14, 
    6.046612e-14, 6.056434e-14, 6.078394e-14, 6.074438e-14, 6.081144e-14, 
    6.087552e-14, 6.0983e-14, 6.096532e-14, 6.101264e-14, 6.080969e-14, 
    6.094459e-14, 6.072183e-14, 6.078279e-14, 6.029708e-14, 6.011182e-14, 
    6.003287e-14, 5.996385e-14, 5.979569e-14, 5.991183e-14, 5.986605e-14, 
    5.997497e-14, 6.004412e-14, 6.000993e-14, 6.022086e-14, 6.013889e-14, 
    6.057016e-14, 6.038455e-14, 6.086805e-14, 6.07525e-14, 6.089573e-14, 
    6.082267e-14, 6.094782e-14, 6.083519e-14, 6.103026e-14, 6.107267e-14, 
    6.104369e-14, 6.115507e-14, 6.082895e-14, 6.095426e-14, 6.000896e-14, 
    6.001454e-14, 6.004053e-14, 5.992625e-14, 5.991926e-14, 5.98145e-14, 
    5.990773e-14, 5.994741e-14, 6.004814e-14, 6.010766e-14, 6.016423e-14, 
    6.028853e-14, 6.042721e-14, 6.062095e-14, 6.076e-14, 6.085312e-14, 
    6.079603e-14, 6.084644e-14, 6.079009e-14, 6.076368e-14, 6.105677e-14, 
    6.089226e-14, 6.113905e-14, 6.112541e-14, 6.101376e-14, 6.112695e-14, 
    6.001846e-14, 5.998637e-14, 5.987484e-14, 5.996213e-14, 5.980309e-14, 
    5.989211e-14, 5.994326e-14, 6.014057e-14, 6.018392e-14, 6.022406e-14, 
    6.030334e-14, 6.0405e-14, 6.058316e-14, 6.073802e-14, 6.087925e-14, 
    6.086891e-14, 6.087255e-14, 6.090407e-14, 6.082596e-14, 6.091689e-14, 
    6.093213e-14, 6.089226e-14, 6.112358e-14, 6.105754e-14, 6.112512e-14, 
    6.108213e-14, 5.99968e-14, 6.00508e-14, 6.002162e-14, 6.007648e-14, 
    6.003782e-14, 6.020959e-14, 6.026105e-14, 6.050164e-14, 6.040299e-14, 
    6.056001e-14, 6.041896e-14, 6.044395e-14, 6.056506e-14, 6.04266e-14, 
    6.072945e-14, 6.052413e-14, 6.090529e-14, 6.070045e-14, 6.091812e-14, 
    6.087864e-14, 6.094401e-14, 6.100251e-14, 6.10761e-14, 6.121174e-14, 
    6.118035e-14, 6.129373e-14, 6.013128e-14, 6.020123e-14, 6.019511e-14, 
    6.026831e-14, 6.032241e-14, 6.043965e-14, 6.062745e-14, 6.055687e-14, 
    6.068645e-14, 6.071244e-14, 6.051558e-14, 6.063645e-14, 6.024806e-14, 
    6.031085e-14, 6.027349e-14, 6.013678e-14, 6.057309e-14, 6.034932e-14, 
    6.076229e-14, 6.064127e-14, 6.099416e-14, 6.081875e-14, 6.116306e-14, 
    6.13099e-14, 6.144811e-14, 6.160927e-14, 6.023943e-14, 6.019191e-14, 
    6.027702e-14, 6.039463e-14, 6.050375e-14, 6.064865e-14, 6.066348e-14, 
    6.06906e-14, 6.076086e-14, 6.081989e-14, 6.069915e-14, 6.083469e-14, 
    6.032535e-14, 6.059252e-14, 6.017391e-14, 6.030005e-14, 6.038771e-14, 
    6.03493e-14, 6.05488e-14, 6.059577e-14, 6.078648e-14, 6.068795e-14, 
    6.127365e-14, 6.101482e-14, 6.173194e-14, 6.153191e-14, 6.017529e-14, 
    6.023928e-14, 6.046172e-14, 6.035593e-14, 6.065833e-14, 6.073266e-14, 
    6.079308e-14, 6.087023e-14, 6.087858e-14, 6.092426e-14, 6.084938e-14, 
    6.092132e-14, 6.064896e-14, 6.077074e-14, 6.043635e-14, 6.051779e-14, 
    6.048034e-14, 6.043922e-14, 6.056607e-14, 6.070104e-14, 6.070397e-14, 
    6.074721e-14, 6.086891e-14, 6.065956e-14, 6.130693e-14, 6.09074e-14, 
    6.030902e-14, 6.043207e-14, 6.044969e-14, 6.040203e-14, 6.072521e-14, 
    6.060819e-14, 6.092316e-14, 6.083811e-14, 6.097744e-14, 6.090822e-14, 
    6.089803e-14, 6.080908e-14, 6.075365e-14, 6.061355e-14, 6.049946e-14, 
    6.040895e-14, 6.043001e-14, 6.052941e-14, 6.07093e-14, 6.087931e-14, 
    6.084208e-14, 6.096686e-14, 6.063643e-14, 6.077505e-14, 6.072147e-14, 
    6.086115e-14, 6.055498e-14, 6.081559e-14, 6.048827e-14, 6.051701e-14, 
    6.060586e-14, 6.078442e-14, 6.082397e-14, 6.086609e-14, 6.084011e-14, 
    6.071388e-14, 6.069321e-14, 6.060372e-14, 6.057898e-14, 6.051076e-14, 
    6.045423e-14, 6.050587e-14, 6.056006e-14, 6.071395e-14, 6.085246e-14, 
    6.100333e-14, 6.104025e-14, 6.121616e-14, 6.107291e-14, 6.130914e-14, 
    6.110823e-14, 6.145589e-14, 6.083075e-14, 6.110242e-14, 6.060992e-14, 
    6.066308e-14, 6.075911e-14, 6.097923e-14, 6.086049e-14, 6.099937e-14, 
    6.06924e-14, 6.053282e-14, 6.049156e-14, 6.041445e-14, 6.049332e-14, 
    6.048691e-14, 6.056234e-14, 6.053811e-14, 6.071906e-14, 6.062189e-14, 
    6.089776e-14, 6.099828e-14, 6.128183e-14, 6.145533e-14, 6.163179e-14, 
    6.170959e-14, 6.173327e-14, 6.174316e-14 ;

 LITTERC =
  5.976256e-05, 5.976241e-05, 5.976244e-05, 5.976232e-05, 5.976239e-05, 
    5.976231e-05, 5.976253e-05, 5.976241e-05, 5.976249e-05, 5.976254e-05, 
    5.976209e-05, 5.976231e-05, 5.976186e-05, 5.9762e-05, 5.976164e-05, 
    5.976188e-05, 5.976159e-05, 5.976165e-05, 5.976148e-05, 5.976153e-05, 
    5.976132e-05, 5.976146e-05, 5.976121e-05, 5.976135e-05, 5.976133e-05, 
    5.976146e-05, 5.976227e-05, 5.976212e-05, 5.976228e-05, 5.976226e-05, 
    5.976227e-05, 5.976238e-05, 5.976245e-05, 5.976257e-05, 5.976255e-05, 
    5.976246e-05, 5.976225e-05, 5.976232e-05, 5.976214e-05, 5.976214e-05, 
    5.976195e-05, 5.976203e-05, 5.97617e-05, 5.97618e-05, 5.976153e-05, 
    5.976159e-05, 5.976153e-05, 5.976155e-05, 5.976153e-05, 5.976163e-05, 
    5.976159e-05, 5.976167e-05, 5.976202e-05, 5.976192e-05, 5.976222e-05, 
    5.97624e-05, 5.976252e-05, 5.976261e-05, 5.97626e-05, 5.976257e-05, 
    5.976246e-05, 5.976234e-05, 5.976226e-05, 5.97622e-05, 5.976214e-05, 
    5.976198e-05, 5.976189e-05, 5.976169e-05, 5.976172e-05, 5.976166e-05, 
    5.97616e-05, 5.97615e-05, 5.976152e-05, 5.976148e-05, 5.976166e-05, 
    5.976154e-05, 5.976174e-05, 5.976169e-05, 5.976213e-05, 5.97623e-05, 
    5.976237e-05, 5.976243e-05, 5.976259e-05, 5.976248e-05, 5.976252e-05, 
    5.976242e-05, 5.976236e-05, 5.976239e-05, 5.97622e-05, 5.976227e-05, 
    5.976188e-05, 5.976205e-05, 5.976161e-05, 5.976171e-05, 5.976158e-05, 
    5.976165e-05, 5.976154e-05, 5.976164e-05, 5.976146e-05, 5.976142e-05, 
    5.976145e-05, 5.976135e-05, 5.976165e-05, 5.976153e-05, 5.976239e-05, 
    5.976239e-05, 5.976237e-05, 5.976247e-05, 5.976247e-05, 5.976257e-05, 
    5.976249e-05, 5.976245e-05, 5.976236e-05, 5.97623e-05, 5.976225e-05, 
    5.976214e-05, 5.976201e-05, 5.976183e-05, 5.976171e-05, 5.976162e-05, 
    5.976167e-05, 5.976163e-05, 5.976168e-05, 5.97617e-05, 5.976144e-05, 
    5.976159e-05, 5.976136e-05, 5.976137e-05, 5.976147e-05, 5.976137e-05, 
    5.976238e-05, 5.976241e-05, 5.976251e-05, 5.976243e-05, 5.976258e-05, 
    5.97625e-05, 5.976245e-05, 5.976227e-05, 5.976223e-05, 5.97622e-05, 
    5.976213e-05, 5.976203e-05, 5.976187e-05, 5.976173e-05, 5.97616e-05, 
    5.976161e-05, 5.976161e-05, 5.976158e-05, 5.976165e-05, 5.976157e-05, 
    5.976155e-05, 5.976159e-05, 5.976138e-05, 5.976143e-05, 5.976137e-05, 
    5.976141e-05, 5.976241e-05, 5.976235e-05, 5.976238e-05, 5.976233e-05, 
    5.976237e-05, 5.976221e-05, 5.976216e-05, 5.976194e-05, 5.976203e-05, 
    5.976189e-05, 5.976202e-05, 5.976199e-05, 5.976189e-05, 5.976201e-05, 
    5.976174e-05, 5.976192e-05, 5.976158e-05, 5.976176e-05, 5.976156e-05, 
    5.97616e-05, 5.976154e-05, 5.976149e-05, 5.976142e-05, 5.97613e-05, 
    5.976133e-05, 5.976122e-05, 5.976228e-05, 5.976222e-05, 5.976222e-05, 
    5.976215e-05, 5.976211e-05, 5.9762e-05, 5.976183e-05, 5.976189e-05, 
    5.976178e-05, 5.976175e-05, 5.976193e-05, 5.976182e-05, 5.976218e-05, 
    5.976212e-05, 5.976215e-05, 5.976227e-05, 5.976188e-05, 5.976208e-05, 
    5.976171e-05, 5.976182e-05, 5.976149e-05, 5.976165e-05, 5.976134e-05, 
    5.976121e-05, 5.976108e-05, 5.976093e-05, 5.976218e-05, 5.976223e-05, 
    5.976215e-05, 5.976204e-05, 5.976194e-05, 5.976181e-05, 5.976179e-05, 
    5.976177e-05, 5.976171e-05, 5.976165e-05, 5.976176e-05, 5.976164e-05, 
    5.97621e-05, 5.976186e-05, 5.976224e-05, 5.976213e-05, 5.976205e-05, 
    5.976208e-05, 5.97619e-05, 5.976186e-05, 5.976168e-05, 5.976177e-05, 
    5.976124e-05, 5.976147e-05, 5.976082e-05, 5.9761e-05, 5.976224e-05, 
    5.976218e-05, 5.976198e-05, 5.976207e-05, 5.97618e-05, 5.976173e-05, 
    5.976168e-05, 5.976161e-05, 5.97616e-05, 5.976156e-05, 5.976163e-05, 
    5.976156e-05, 5.976181e-05, 5.97617e-05, 5.9762e-05, 5.976193e-05, 
    5.976196e-05, 5.9762e-05, 5.976189e-05, 5.976176e-05, 5.976176e-05, 
    5.976172e-05, 5.976161e-05, 5.97618e-05, 5.976121e-05, 5.976157e-05, 
    5.976212e-05, 5.976201e-05, 5.976199e-05, 5.976203e-05, 5.976174e-05, 
    5.976185e-05, 5.976156e-05, 5.976163e-05, 5.976151e-05, 5.976157e-05, 
    5.976158e-05, 5.976166e-05, 5.976171e-05, 5.976184e-05, 5.976194e-05, 
    5.976203e-05, 5.976201e-05, 5.976192e-05, 5.976175e-05, 5.97616e-05, 
    5.976163e-05, 5.976152e-05, 5.976182e-05, 5.976169e-05, 5.976174e-05, 
    5.976162e-05, 5.97619e-05, 5.976166e-05, 5.976195e-05, 5.976193e-05, 
    5.976185e-05, 5.976169e-05, 5.976165e-05, 5.976161e-05, 5.976163e-05, 
    5.976175e-05, 5.976177e-05, 5.976185e-05, 5.976187e-05, 5.976194e-05, 
    5.976199e-05, 5.976194e-05, 5.976189e-05, 5.976175e-05, 5.976162e-05, 
    5.976149e-05, 5.976145e-05, 5.976129e-05, 5.976142e-05, 5.976121e-05, 
    5.976139e-05, 5.976107e-05, 5.976164e-05, 5.976139e-05, 5.976185e-05, 
    5.976179e-05, 5.976171e-05, 5.976151e-05, 5.976162e-05, 5.976149e-05, 
    5.976177e-05, 5.976191e-05, 5.976195e-05, 5.976202e-05, 5.976195e-05, 
    5.976196e-05, 5.976189e-05, 5.976191e-05, 5.976174e-05, 5.976183e-05, 
    5.976158e-05, 5.976149e-05, 5.976123e-05, 5.976107e-05, 5.976091e-05, 
    5.976084e-05, 5.976082e-05, 5.976081e-05 ;

 LITTERC_HR =
  9.652399e-13, 9.678468e-13, 9.673404e-13, 9.69441e-13, 9.682762e-13, 
    9.696512e-13, 9.65769e-13, 9.679499e-13, 9.665581e-13, 9.654752e-13, 
    9.735113e-13, 9.695348e-13, 9.776379e-13, 9.751066e-13, 9.814612e-13, 
    9.772438e-13, 9.823108e-13, 9.813404e-13, 9.842616e-13, 9.834251e-13, 
    9.871558e-13, 9.846476e-13, 9.890884e-13, 9.865574e-13, 9.869532e-13, 
    9.845646e-13, 9.703362e-13, 9.730164e-13, 9.701772e-13, 9.705597e-13, 
    9.703883e-13, 9.683001e-13, 9.672466e-13, 9.650411e-13, 9.654418e-13, 
    9.670618e-13, 9.707316e-13, 9.69487e-13, 9.726239e-13, 9.725531e-13, 
    9.760401e-13, 9.744686e-13, 9.803222e-13, 9.786601e-13, 9.834602e-13, 
    9.822538e-13, 9.834034e-13, 9.830549e-13, 9.834079e-13, 9.816385e-13, 
    9.823967e-13, 9.808393e-13, 9.747628e-13, 9.765501e-13, 9.712151e-13, 
    9.680003e-13, 9.658645e-13, 9.643473e-13, 9.645619e-13, 9.649706e-13, 
    9.670714e-13, 9.690454e-13, 9.705484e-13, 9.715532e-13, 9.725429e-13, 
    9.755342e-13, 9.771176e-13, 9.806576e-13, 9.800199e-13, 9.811007e-13, 
    9.821338e-13, 9.838663e-13, 9.835813e-13, 9.843441e-13, 9.810728e-13, 
    9.832472e-13, 9.796564e-13, 9.80639e-13, 9.728094e-13, 9.69823e-13, 
    9.685502e-13, 9.674376e-13, 9.647268e-13, 9.66599e-13, 9.658611e-13, 
    9.676169e-13, 9.687315e-13, 9.681804e-13, 9.715807e-13, 9.702592e-13, 
    9.772114e-13, 9.742194e-13, 9.820133e-13, 9.801509e-13, 9.824597e-13, 
    9.812819e-13, 9.832993e-13, 9.814838e-13, 9.846282e-13, 9.85312e-13, 
    9.848446e-13, 9.866401e-13, 9.813831e-13, 9.83403e-13, 9.681649e-13, 
    9.682548e-13, 9.686737e-13, 9.668314e-13, 9.667188e-13, 9.650299e-13, 
    9.66533e-13, 9.671725e-13, 9.687963e-13, 9.697559e-13, 9.706678e-13, 
    9.726715e-13, 9.74907e-13, 9.7803e-13, 9.802715e-13, 9.817727e-13, 
    9.808526e-13, 9.816649e-13, 9.807566e-13, 9.803309e-13, 9.850556e-13, 
    9.824036e-13, 9.86382e-13, 9.861621e-13, 9.843621e-13, 9.861868e-13, 
    9.683179e-13, 9.678006e-13, 9.660028e-13, 9.674099e-13, 9.64846e-13, 
    9.662811e-13, 9.671057e-13, 9.702864e-13, 9.709851e-13, 9.716322e-13, 
    9.729102e-13, 9.74549e-13, 9.774209e-13, 9.799172e-13, 9.82194e-13, 
    9.820273e-13, 9.820859e-13, 9.82594e-13, 9.813349e-13, 9.828006e-13, 
    9.830463e-13, 9.824036e-13, 9.861326e-13, 9.850679e-13, 9.861574e-13, 
    9.854643e-13, 9.679688e-13, 9.688393e-13, 9.683689e-13, 9.692532e-13, 
    9.6863e-13, 9.71399e-13, 9.722285e-13, 9.761069e-13, 9.745166e-13, 
    9.770478e-13, 9.747741e-13, 9.75177e-13, 9.771292e-13, 9.748971e-13, 
    9.797791e-13, 9.764694e-13, 9.826137e-13, 9.793118e-13, 9.828205e-13, 
    9.821842e-13, 9.832379e-13, 9.841808e-13, 9.853672e-13, 9.875536e-13, 
    9.870476e-13, 9.888752e-13, 9.701366e-13, 9.712643e-13, 9.711655e-13, 
    9.723455e-13, 9.732176e-13, 9.751076e-13, 9.781349e-13, 9.769971e-13, 
    9.790861e-13, 9.79505e-13, 9.763315e-13, 9.782801e-13, 9.720191e-13, 
    9.730312e-13, 9.724291e-13, 9.702253e-13, 9.772586e-13, 9.736515e-13, 
    9.803085e-13, 9.783578e-13, 9.840464e-13, 9.812186e-13, 9.867688e-13, 
    9.891361e-13, 9.913638e-13, 9.939616e-13, 9.7188e-13, 9.71114e-13, 
    9.724859e-13, 9.743818e-13, 9.761409e-13, 9.784767e-13, 9.787158e-13, 
    9.79153e-13, 9.802855e-13, 9.81237e-13, 9.792907e-13, 9.814755e-13, 
    9.73265e-13, 9.775718e-13, 9.708239e-13, 9.728572e-13, 9.742703e-13, 
    9.73651e-13, 9.768671e-13, 9.776243e-13, 9.806985e-13, 9.791101e-13, 
    9.885516e-13, 9.843794e-13, 9.959391e-13, 9.927146e-13, 9.708461e-13, 
    9.718776e-13, 9.754633e-13, 9.73758e-13, 9.786328e-13, 9.798309e-13, 
    9.808048e-13, 9.820484e-13, 9.821831e-13, 9.829196e-13, 9.817124e-13, 
    9.828721e-13, 9.784816e-13, 9.804448e-13, 9.750543e-13, 9.763672e-13, 
    9.757635e-13, 9.751008e-13, 9.771456e-13, 9.793212e-13, 9.793685e-13, 
    9.800655e-13, 9.820272e-13, 9.786526e-13, 9.89088e-13, 9.826478e-13, 
    9.730018e-13, 9.749854e-13, 9.752695e-13, 9.745013e-13, 9.797108e-13, 
    9.778245e-13, 9.829017e-13, 9.815308e-13, 9.837768e-13, 9.826609e-13, 
    9.824966e-13, 9.810628e-13, 9.801694e-13, 9.779108e-13, 9.760718e-13, 
    9.746128e-13, 9.749522e-13, 9.765546e-13, 9.794544e-13, 9.821949e-13, 
    9.815947e-13, 9.836062e-13, 9.782796e-13, 9.805143e-13, 9.796506e-13, 
    9.819021e-13, 9.769667e-13, 9.811677e-13, 9.758914e-13, 9.763546e-13, 
    9.77787e-13, 9.806652e-13, 9.813027e-13, 9.819817e-13, 9.815629e-13, 
    9.795281e-13, 9.791949e-13, 9.777524e-13, 9.773535e-13, 9.762538e-13, 
    9.753425e-13, 9.76175e-13, 9.770486e-13, 9.795293e-13, 9.817621e-13, 
    9.841942e-13, 9.847893e-13, 9.876248e-13, 9.853158e-13, 9.891237e-13, 
    9.85885e-13, 9.914891e-13, 9.814121e-13, 9.857913e-13, 9.778525e-13, 
    9.787092e-13, 9.802573e-13, 9.838056e-13, 9.818915e-13, 9.841302e-13, 
    9.791819e-13, 9.766094e-13, 9.759444e-13, 9.747013e-13, 9.759728e-13, 
    9.758695e-13, 9.770854e-13, 9.766947e-13, 9.796117e-13, 9.780453e-13, 
    9.824923e-13, 9.841127e-13, 9.886835e-13, 9.914802e-13, 9.943246e-13, 
    9.955787e-13, 9.959604e-13, 9.961199e-13 ;

 LITTERC_LOSS =
  1.787615e-12, 1.792443e-12, 1.791505e-12, 1.795395e-12, 1.793238e-12, 
    1.795785e-12, 1.788595e-12, 1.792634e-12, 1.790056e-12, 1.788051e-12, 
    1.802934e-12, 1.795569e-12, 1.810576e-12, 1.805888e-12, 1.817657e-12, 
    1.809846e-12, 1.819231e-12, 1.817433e-12, 1.822843e-12, 1.821294e-12, 
    1.828203e-12, 1.823558e-12, 1.831783e-12, 1.827095e-12, 1.827828e-12, 
    1.823405e-12, 1.797053e-12, 1.802017e-12, 1.796759e-12, 1.797467e-12, 
    1.79715e-12, 1.793282e-12, 1.791331e-12, 1.787247e-12, 1.787989e-12, 
    1.790989e-12, 1.797786e-12, 1.795481e-12, 1.80129e-12, 1.801159e-12, 
    1.807617e-12, 1.804706e-12, 1.815547e-12, 1.812469e-12, 1.821359e-12, 
    1.819125e-12, 1.821254e-12, 1.820609e-12, 1.821262e-12, 1.817985e-12, 
    1.819389e-12, 1.816505e-12, 1.805251e-12, 1.808562e-12, 1.798681e-12, 
    1.792727e-12, 1.788772e-12, 1.785962e-12, 1.786359e-12, 1.787116e-12, 
    1.791007e-12, 1.794663e-12, 1.797446e-12, 1.799307e-12, 1.80114e-12, 
    1.80668e-12, 1.809613e-12, 1.816169e-12, 1.814988e-12, 1.816989e-12, 
    1.818903e-12, 1.822111e-12, 1.821583e-12, 1.822996e-12, 1.816937e-12, 
    1.820965e-12, 1.814314e-12, 1.816134e-12, 1.801634e-12, 1.796103e-12, 
    1.793746e-12, 1.791685e-12, 1.786664e-12, 1.790132e-12, 1.788765e-12, 
    1.792017e-12, 1.794081e-12, 1.793061e-12, 1.799358e-12, 1.796911e-12, 
    1.809786e-12, 1.804245e-12, 1.81868e-12, 1.81523e-12, 1.819506e-12, 
    1.817325e-12, 1.821061e-12, 1.817699e-12, 1.823522e-12, 1.824789e-12, 
    1.823923e-12, 1.827248e-12, 1.817512e-12, 1.821253e-12, 1.793032e-12, 
    1.793198e-12, 1.793974e-12, 1.790562e-12, 1.790354e-12, 1.787226e-12, 
    1.79001e-12, 1.791194e-12, 1.794201e-12, 1.795978e-12, 1.797667e-12, 
    1.801378e-12, 1.805519e-12, 1.811303e-12, 1.815454e-12, 1.818234e-12, 
    1.81653e-12, 1.818034e-12, 1.816352e-12, 1.815564e-12, 1.824314e-12, 
    1.819402e-12, 1.82677e-12, 1.826363e-12, 1.82303e-12, 1.826409e-12, 
    1.793315e-12, 1.792357e-12, 1.789028e-12, 1.791634e-12, 1.786885e-12, 
    1.789543e-12, 1.79107e-12, 1.796961e-12, 1.798255e-12, 1.799453e-12, 
    1.80182e-12, 1.804855e-12, 1.810174e-12, 1.814797e-12, 1.819014e-12, 
    1.818705e-12, 1.818814e-12, 1.819755e-12, 1.817423e-12, 1.820138e-12, 
    1.820593e-12, 1.819402e-12, 1.826309e-12, 1.824337e-12, 1.826354e-12, 
    1.825071e-12, 1.792669e-12, 1.794281e-12, 1.79341e-12, 1.795048e-12, 
    1.793893e-12, 1.799021e-12, 1.800558e-12, 1.807741e-12, 1.804795e-12, 
    1.809483e-12, 1.805272e-12, 1.806018e-12, 1.809634e-12, 1.8055e-12, 
    1.814542e-12, 1.808412e-12, 1.819791e-12, 1.813676e-12, 1.820174e-12, 
    1.818996e-12, 1.820947e-12, 1.822694e-12, 1.824891e-12, 1.82894e-12, 
    1.828003e-12, 1.831388e-12, 1.796684e-12, 1.798772e-12, 1.798589e-12, 
    1.800774e-12, 1.80239e-12, 1.80589e-12, 1.811497e-12, 1.809389e-12, 
    1.813258e-12, 1.814034e-12, 1.808157e-12, 1.811765e-12, 1.80017e-12, 
    1.802045e-12, 1.800929e-12, 1.796848e-12, 1.809874e-12, 1.803193e-12, 
    1.815522e-12, 1.811909e-12, 1.822445e-12, 1.817208e-12, 1.827487e-12, 
    1.831871e-12, 1.835997e-12, 1.840808e-12, 1.799913e-12, 1.798494e-12, 
    1.801035e-12, 1.804546e-12, 1.807804e-12, 1.81213e-12, 1.812572e-12, 
    1.813382e-12, 1.81548e-12, 1.817242e-12, 1.813637e-12, 1.817683e-12, 
    1.802477e-12, 1.810454e-12, 1.797956e-12, 1.801722e-12, 1.804339e-12, 
    1.803192e-12, 1.809149e-12, 1.810551e-12, 1.816245e-12, 1.813303e-12, 
    1.830789e-12, 1.823061e-12, 1.844471e-12, 1.838499e-12, 1.797998e-12, 
    1.799908e-12, 1.806549e-12, 1.803391e-12, 1.812419e-12, 1.814638e-12, 
    1.816441e-12, 1.818745e-12, 1.818994e-12, 1.820358e-12, 1.818122e-12, 
    1.82027e-12, 1.812139e-12, 1.815775e-12, 1.805791e-12, 1.808223e-12, 
    1.807105e-12, 1.805877e-12, 1.809664e-12, 1.813694e-12, 1.813781e-12, 
    1.815072e-12, 1.818705e-12, 1.812455e-12, 1.831782e-12, 1.819855e-12, 
    1.80199e-12, 1.805664e-12, 1.80619e-12, 1.804767e-12, 1.814415e-12, 
    1.810922e-12, 1.820325e-12, 1.817786e-12, 1.821945e-12, 1.819879e-12, 
    1.819575e-12, 1.816919e-12, 1.815265e-12, 1.811082e-12, 1.807676e-12, 
    1.804974e-12, 1.805602e-12, 1.80857e-12, 1.81394e-12, 1.819016e-12, 
    1.817904e-12, 1.821629e-12, 1.811765e-12, 1.815903e-12, 1.814304e-12, 
    1.818474e-12, 1.809333e-12, 1.817114e-12, 1.807341e-12, 1.8082e-12, 
    1.810852e-12, 1.816183e-12, 1.817363e-12, 1.818621e-12, 1.817845e-12, 
    1.814077e-12, 1.81346e-12, 1.810788e-12, 1.81005e-12, 1.808013e-12, 
    1.806325e-12, 1.807867e-12, 1.809485e-12, 1.814079e-12, 1.818214e-12, 
    1.822719e-12, 1.823821e-12, 1.829072e-12, 1.824796e-12, 1.831848e-12, 
    1.82585e-12, 1.836229e-12, 1.817566e-12, 1.825676e-12, 1.810973e-12, 
    1.81256e-12, 1.815427e-12, 1.821999e-12, 1.818454e-12, 1.8226e-12, 
    1.813436e-12, 1.808671e-12, 1.80744e-12, 1.805138e-12, 1.807492e-12, 
    1.807301e-12, 1.809553e-12, 1.808829e-12, 1.814232e-12, 1.811331e-12, 
    1.819567e-12, 1.822568e-12, 1.831033e-12, 1.836212e-12, 1.84148e-12, 
    1.843803e-12, 1.84451e-12, 1.844805e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.676328e-18, 1.676591e-18, 1.676541e-18, 1.676751e-18, 1.676636e-18, 
    1.676772e-18, 1.676384e-18, 1.676599e-18, 1.676463e-18, 1.676355e-18, 
    1.677151e-18, 1.676761e-18, 1.67758e-18, 1.677327e-18, 1.677971e-18, 
    1.677538e-18, 1.67806e-18, 1.677964e-18, 1.678265e-18, 1.678179e-18, 
    1.678554e-18, 1.678305e-18, 1.678757e-18, 1.678497e-18, 1.678536e-18, 
    1.678296e-18, 1.676844e-18, 1.677101e-18, 1.676828e-18, 1.676865e-18, 
    1.676849e-18, 1.676637e-18, 1.676527e-18, 1.676311e-18, 1.676351e-18, 
    1.676511e-18, 1.676881e-18, 1.676759e-18, 1.677077e-18, 1.67707e-18, 
    1.677422e-18, 1.677263e-18, 1.677859e-18, 1.677691e-18, 1.678183e-18, 
    1.678058e-18, 1.678176e-18, 1.678141e-18, 1.678176e-18, 1.677994e-18, 
    1.678072e-18, 1.677913e-18, 1.677292e-18, 1.677473e-18, 1.676932e-18, 
    1.6766e-18, 1.676392e-18, 1.676241e-18, 1.676262e-18, 1.676302e-18, 
    1.676512e-18, 1.676714e-18, 1.676867e-18, 1.676968e-18, 1.677069e-18, 
    1.677361e-18, 1.677527e-18, 1.677891e-18, 1.67783e-18, 1.677937e-18, 
    1.678046e-18, 1.678223e-18, 1.678194e-18, 1.678271e-18, 1.677937e-18, 
    1.678158e-18, 1.677794e-18, 1.677893e-18, 1.677079e-18, 1.676793e-18, 
    1.676656e-18, 1.67655e-18, 1.676279e-18, 1.676465e-18, 1.676391e-18, 
    1.676571e-18, 1.676682e-18, 1.676628e-18, 1.676971e-18, 1.676837e-18, 
    1.677537e-18, 1.677235e-18, 1.678033e-18, 1.677843e-18, 1.678079e-18, 
    1.677959e-18, 1.678164e-18, 1.67798e-18, 1.678301e-18, 1.67837e-18, 
    1.678323e-18, 1.678509e-18, 1.677969e-18, 1.678174e-18, 1.676626e-18, 
    1.676634e-18, 1.676677e-18, 1.676488e-18, 1.676478e-18, 1.676309e-18, 
    1.676461e-18, 1.676524e-18, 1.67669e-18, 1.676786e-18, 1.676878e-18, 
    1.677081e-18, 1.677304e-18, 1.677623e-18, 1.677855e-18, 1.67801e-18, 
    1.677916e-18, 1.677998e-18, 1.677905e-18, 1.677862e-18, 1.678343e-18, 
    1.678071e-18, 1.678482e-18, 1.67846e-18, 1.678273e-18, 1.678462e-18, 
    1.676641e-18, 1.67659e-18, 1.676407e-18, 1.67655e-18, 1.676291e-18, 
    1.676434e-18, 1.676515e-18, 1.676836e-18, 1.676911e-18, 1.676975e-18, 
    1.677106e-18, 1.677271e-18, 1.677561e-18, 1.677817e-18, 1.678053e-18, 
    1.678036e-18, 1.678042e-18, 1.678093e-18, 1.677964e-18, 1.678114e-18, 
    1.678137e-18, 1.678073e-18, 1.678457e-18, 1.678347e-18, 1.678459e-18, 
    1.678389e-18, 1.676607e-18, 1.676694e-18, 1.676646e-18, 1.676734e-18, 
    1.676671e-18, 1.676948e-18, 1.677031e-18, 1.677424e-18, 1.677267e-18, 
    1.677522e-18, 1.677294e-18, 1.677334e-18, 1.677523e-18, 1.677308e-18, 
    1.677799e-18, 1.677459e-18, 1.678095e-18, 1.677748e-18, 1.678116e-18, 
    1.678052e-18, 1.67816e-18, 1.678255e-18, 1.678378e-18, 1.6786e-18, 
    1.678549e-18, 1.678738e-18, 1.676825e-18, 1.676936e-18, 1.67693e-18, 
    1.677048e-18, 1.677136e-18, 1.677329e-18, 1.677636e-18, 1.677521e-18, 
    1.677735e-18, 1.677777e-18, 1.677454e-18, 1.677649e-18, 1.677013e-18, 
    1.677112e-18, 1.677056e-18, 1.676832e-18, 1.677543e-18, 1.677176e-18, 
    1.677858e-18, 1.677659e-18, 1.678241e-18, 1.677948e-18, 1.67852e-18, 
    1.678757e-18, 1.678996e-18, 1.679258e-18, 1.677e-18, 1.676924e-18, 
    1.677064e-18, 1.67725e-18, 1.677433e-18, 1.677671e-18, 1.677697e-18, 
    1.67774e-18, 1.677858e-18, 1.677954e-18, 1.677751e-18, 1.677979e-18, 
    1.677129e-18, 1.677576e-18, 1.676893e-18, 1.677094e-18, 1.677241e-18, 
    1.67718e-18, 1.677509e-18, 1.677586e-18, 1.677896e-18, 1.677737e-18, 
    1.678696e-18, 1.67827e-18, 1.679468e-18, 1.67913e-18, 1.676897e-18, 
    1.677002e-18, 1.677362e-18, 1.677191e-18, 1.677688e-18, 1.677809e-18, 
    1.677911e-18, 1.678035e-18, 1.678051e-18, 1.678125e-18, 1.678003e-18, 
    1.678122e-18, 1.677671e-18, 1.677873e-18, 1.677324e-18, 1.677456e-18, 
    1.677396e-18, 1.677329e-18, 1.677537e-18, 1.677753e-18, 1.677763e-18, 
    1.677832e-18, 1.678016e-18, 1.67769e-18, 1.678741e-18, 1.678082e-18, 
    1.677116e-18, 1.67731e-18, 1.677344e-18, 1.677268e-18, 1.677797e-18, 
    1.677604e-18, 1.678124e-18, 1.677985e-18, 1.678215e-18, 1.6781e-18, 
    1.678083e-18, 1.677937e-18, 1.677844e-18, 1.677612e-18, 1.677425e-18, 
    1.67728e-18, 1.677314e-18, 1.677474e-18, 1.677768e-18, 1.67805e-18, 
    1.677988e-18, 1.678197e-18, 1.677652e-18, 1.677878e-18, 1.677789e-18, 
    1.678022e-18, 1.677517e-18, 1.677931e-18, 1.677409e-18, 1.677456e-18, 
    1.677601e-18, 1.677889e-18, 1.677961e-18, 1.678029e-18, 1.677988e-18, 
    1.677776e-18, 1.677744e-18, 1.677598e-18, 1.677556e-18, 1.677446e-18, 
    1.677354e-18, 1.677437e-18, 1.677524e-18, 1.677779e-18, 1.678006e-18, 
    1.678256e-18, 1.678319e-18, 1.678598e-18, 1.678364e-18, 1.678744e-18, 
    1.678409e-18, 1.678994e-18, 1.677963e-18, 1.67841e-18, 1.677609e-18, 
    1.677696e-18, 1.677849e-18, 1.678211e-18, 1.678021e-18, 1.678246e-18, 
    1.677743e-18, 1.677477e-18, 1.677414e-18, 1.677287e-18, 1.677417e-18, 
    1.677407e-18, 1.677531e-18, 1.677492e-18, 1.677787e-18, 1.677628e-18, 
    1.678081e-18, 1.678245e-18, 1.678716e-18, 1.679002e-18, 1.679303e-18, 
    1.679433e-18, 1.679473e-18, 1.679489e-18 ;

 MEG_acetic_acid =
  2.514492e-19, 2.514887e-19, 2.514812e-19, 2.515126e-19, 2.514954e-19, 
    2.515158e-19, 2.514575e-19, 2.514899e-19, 2.514694e-19, 2.514532e-19, 
    2.515727e-19, 2.515141e-19, 2.51637e-19, 2.51599e-19, 2.516957e-19, 
    2.516306e-19, 2.517089e-19, 2.516945e-19, 2.517397e-19, 2.517268e-19, 
    2.517831e-19, 2.517457e-19, 2.518136e-19, 2.517746e-19, 2.517804e-19, 
    2.517443e-19, 2.515266e-19, 2.515652e-19, 2.515241e-19, 2.515297e-19, 
    2.515274e-19, 2.514955e-19, 2.51479e-19, 2.514467e-19, 2.514527e-19, 
    2.514767e-19, 2.515322e-19, 2.515139e-19, 2.515616e-19, 2.515605e-19, 
    2.516133e-19, 2.515895e-19, 2.516789e-19, 2.516536e-19, 2.517274e-19, 
    2.517087e-19, 2.517264e-19, 2.517211e-19, 2.517264e-19, 2.516991e-19, 
    2.517108e-19, 2.516869e-19, 2.515938e-19, 2.516209e-19, 2.515398e-19, 
    2.514899e-19, 2.514588e-19, 2.514362e-19, 2.514394e-19, 2.514453e-19, 
    2.514768e-19, 2.515072e-19, 2.515301e-19, 2.515453e-19, 2.515604e-19, 
    2.516042e-19, 2.516291e-19, 2.516836e-19, 2.516744e-19, 2.516905e-19, 
    2.517069e-19, 2.517334e-19, 2.517292e-19, 2.517407e-19, 2.516906e-19, 
    2.517236e-19, 2.51669e-19, 2.516839e-19, 2.515619e-19, 2.515189e-19, 
    2.514984e-19, 2.514825e-19, 2.514418e-19, 2.514698e-19, 2.514586e-19, 
    2.514856e-19, 2.515024e-19, 2.514942e-19, 2.515457e-19, 2.515256e-19, 
    2.516305e-19, 2.515853e-19, 2.51705e-19, 2.516764e-19, 2.517119e-19, 
    2.516939e-19, 2.517246e-19, 2.51697e-19, 2.517452e-19, 2.517554e-19, 
    2.517484e-19, 2.517763e-19, 2.516954e-19, 2.517261e-19, 2.514938e-19, 
    2.514951e-19, 2.515016e-19, 2.514732e-19, 2.514716e-19, 2.514464e-19, 
    2.514691e-19, 2.514785e-19, 2.515035e-19, 2.515179e-19, 2.515317e-19, 
    2.515621e-19, 2.515956e-19, 2.516434e-19, 2.516782e-19, 2.517014e-19, 
    2.516874e-19, 2.516998e-19, 2.516858e-19, 2.516794e-19, 2.517514e-19, 
    2.517107e-19, 2.517723e-19, 2.51769e-19, 2.517409e-19, 2.517694e-19, 
    2.514961e-19, 2.514884e-19, 2.51461e-19, 2.514825e-19, 2.514437e-19, 
    2.514651e-19, 2.514772e-19, 2.515254e-19, 2.515366e-19, 2.515462e-19, 
    2.515658e-19, 2.515907e-19, 2.516342e-19, 2.516725e-19, 2.517079e-19, 
    2.517054e-19, 2.517063e-19, 2.517139e-19, 2.516946e-19, 2.517171e-19, 
    2.517206e-19, 2.51711e-19, 2.517685e-19, 2.517521e-19, 2.517689e-19, 
    2.517583e-19, 2.51491e-19, 2.51504e-19, 2.514969e-19, 2.515101e-19, 
    2.515006e-19, 2.515421e-19, 2.515546e-19, 2.516137e-19, 2.515901e-19, 
    2.516284e-19, 2.515941e-19, 2.516001e-19, 2.516285e-19, 2.515962e-19, 
    2.516699e-19, 2.516189e-19, 2.517142e-19, 2.516621e-19, 2.517174e-19, 
    2.517078e-19, 2.51724e-19, 2.517383e-19, 2.517567e-19, 2.5179e-19, 
    2.517824e-19, 2.518107e-19, 2.515237e-19, 2.515404e-19, 2.515394e-19, 
    2.515573e-19, 2.515703e-19, 2.515993e-19, 2.516453e-19, 2.516282e-19, 
    2.516602e-19, 2.516665e-19, 2.516181e-19, 2.516473e-19, 2.51552e-19, 
    2.515668e-19, 2.515583e-19, 2.515248e-19, 2.516314e-19, 2.515763e-19, 
    2.516787e-19, 2.516488e-19, 2.517361e-19, 2.516922e-19, 2.517781e-19, 
    2.518136e-19, 2.518494e-19, 2.518886e-19, 2.515501e-19, 2.515387e-19, 
    2.515595e-19, 2.515875e-19, 2.516149e-19, 2.516506e-19, 2.516545e-19, 
    2.51661e-19, 2.516786e-19, 2.516932e-19, 2.516626e-19, 2.516969e-19, 
    2.515693e-19, 2.516365e-19, 2.515339e-19, 2.515641e-19, 2.515861e-19, 
    2.515769e-19, 2.516263e-19, 2.516378e-19, 2.516844e-19, 2.516606e-19, 
    2.518044e-19, 2.517406e-19, 2.519202e-19, 2.518695e-19, 2.515346e-19, 
    2.515503e-19, 2.516042e-19, 2.515786e-19, 2.516532e-19, 2.516714e-19, 
    2.516866e-19, 2.517053e-19, 2.517077e-19, 2.517188e-19, 2.517005e-19, 
    2.517183e-19, 2.516507e-19, 2.516809e-19, 2.515986e-19, 2.516183e-19, 
    2.516094e-19, 2.515993e-19, 2.516305e-19, 2.51663e-19, 2.516645e-19, 
    2.516748e-19, 2.517024e-19, 2.516535e-19, 2.518112e-19, 2.517123e-19, 
    2.515673e-19, 2.515965e-19, 2.516017e-19, 2.515902e-19, 2.516695e-19, 
    2.516406e-19, 2.517186e-19, 2.516977e-19, 2.517322e-19, 2.51715e-19, 
    2.517124e-19, 2.516905e-19, 2.516767e-19, 2.516418e-19, 2.516138e-19, 
    2.515919e-19, 2.515971e-19, 2.516211e-19, 2.516652e-19, 2.517075e-19, 
    2.516981e-19, 2.517296e-19, 2.516478e-19, 2.516816e-19, 2.516683e-19, 
    2.517033e-19, 2.516275e-19, 2.516896e-19, 2.516114e-19, 2.516184e-19, 
    2.516401e-19, 2.516834e-19, 2.516942e-19, 2.517043e-19, 2.516982e-19, 
    2.516664e-19, 2.516616e-19, 2.516397e-19, 2.516333e-19, 2.51617e-19, 
    2.51603e-19, 2.516156e-19, 2.516285e-19, 2.516668e-19, 2.517008e-19, 
    2.517383e-19, 2.517478e-19, 2.517897e-19, 2.517545e-19, 2.518116e-19, 
    2.517614e-19, 2.518491e-19, 2.516944e-19, 2.517615e-19, 2.516413e-19, 
    2.516545e-19, 2.516773e-19, 2.517316e-19, 2.517031e-19, 2.517368e-19, 
    2.516615e-19, 2.516215e-19, 2.516122e-19, 2.515931e-19, 2.516126e-19, 
    2.51611e-19, 2.516297e-19, 2.516237e-19, 2.51668e-19, 2.516443e-19, 
    2.517121e-19, 2.517368e-19, 2.518074e-19, 2.518503e-19, 2.518954e-19, 
    2.519149e-19, 2.519209e-19, 2.519234e-19 ;

 MEG_acetone =
  8.435572e-17, 8.436433e-17, 8.436269e-17, 8.436956e-17, 8.436581e-17, 
    8.437026e-17, 8.435754e-17, 8.436461e-17, 8.436014e-17, 8.43566e-17, 
    8.438267e-17, 8.436988e-17, 8.43967e-17, 8.43884e-17, 8.44095e-17, 
    8.439531e-17, 8.44124e-17, 8.440926e-17, 8.441913e-17, 8.441631e-17, 
    8.442859e-17, 8.442043e-17, 8.443525e-17, 8.442673e-17, 8.4428e-17, 
    8.442013e-17, 8.437261e-17, 8.438103e-17, 8.437208e-17, 8.437328e-17, 
    8.437278e-17, 8.436583e-17, 8.436222e-17, 8.435518e-17, 8.435649e-17, 
    8.436172e-17, 8.437383e-17, 8.436983e-17, 8.438025e-17, 8.438002e-17, 
    8.439153e-17, 8.438633e-17, 8.440585e-17, 8.440033e-17, 8.441643e-17, 
    8.441235e-17, 8.441621e-17, 8.441506e-17, 8.441622e-17, 8.441025e-17, 
    8.44128e-17, 8.440761e-17, 8.438727e-17, 8.439319e-17, 8.437548e-17, 
    8.436461e-17, 8.435782e-17, 8.435288e-17, 8.435358e-17, 8.435487e-17, 
    8.436175e-17, 8.436837e-17, 8.437337e-17, 8.437668e-17, 8.437999e-17, 
    8.438954e-17, 8.439497e-17, 8.440688e-17, 8.440487e-17, 8.440839e-17, 
    8.441196e-17, 8.441775e-17, 8.441682e-17, 8.441934e-17, 8.44084e-17, 
    8.441561e-17, 8.44037e-17, 8.440693e-17, 8.43803e-17, 8.437093e-17, 
    8.436647e-17, 8.436299e-17, 8.43541e-17, 8.436021e-17, 8.435778e-17, 
    8.436367e-17, 8.436733e-17, 8.436554e-17, 8.437678e-17, 8.437238e-17, 
    8.439529e-17, 8.438542e-17, 8.441154e-17, 8.44053e-17, 8.441305e-17, 
    8.440912e-17, 8.441581e-17, 8.440979e-17, 8.442033e-17, 8.442256e-17, 
    8.442101e-17, 8.442712e-17, 8.440945e-17, 8.441616e-17, 8.436546e-17, 
    8.436575e-17, 8.436715e-17, 8.436096e-17, 8.436062e-17, 8.435512e-17, 
    8.436006e-17, 8.436212e-17, 8.436759e-17, 8.437071e-17, 8.437372e-17, 
    8.438035e-17, 8.438768e-17, 8.43981e-17, 8.440569e-17, 8.441076e-17, 
    8.440769e-17, 8.44104e-17, 8.440736e-17, 8.440595e-17, 8.442168e-17, 
    8.441279e-17, 8.442624e-17, 8.442551e-17, 8.441937e-17, 8.442559e-17, 
    8.436596e-17, 8.436429e-17, 8.435829e-17, 8.436299e-17, 8.435452e-17, 
    8.435919e-17, 8.436183e-17, 8.437235e-17, 8.43748e-17, 8.43769e-17, 
    8.438118e-17, 8.43866e-17, 8.439609e-17, 8.440445e-17, 8.441219e-17, 
    8.441163e-17, 8.441182e-17, 8.441349e-17, 8.440928e-17, 8.441419e-17, 
    8.441495e-17, 8.441286e-17, 8.442541e-17, 8.442183e-17, 8.442549e-17, 
    8.442318e-17, 8.436485e-17, 8.436769e-17, 8.436614e-17, 8.436902e-17, 
    8.436695e-17, 8.4376e-17, 8.437872e-17, 8.439161e-17, 8.438646e-17, 
    8.439482e-17, 8.438735e-17, 8.438864e-17, 8.439485e-17, 8.438779e-17, 
    8.440388e-17, 8.439275e-17, 8.441356e-17, 8.440219e-17, 8.441425e-17, 
    8.441215e-17, 8.441569e-17, 8.44188e-17, 8.442283e-17, 8.443009e-17, 
    8.442843e-17, 8.443461e-17, 8.437199e-17, 8.437563e-17, 8.437541e-17, 
    8.43793e-17, 8.438216e-17, 8.438848e-17, 8.439852e-17, 8.439478e-17, 
    8.440177e-17, 8.440313e-17, 8.439258e-17, 8.439895e-17, 8.437815e-17, 
    8.438139e-17, 8.437954e-17, 8.437221e-17, 8.439549e-17, 8.438346e-17, 
    8.44058e-17, 8.439929e-17, 8.441835e-17, 8.440875e-17, 8.442749e-17, 
    8.443525e-17, 8.444307e-17, 8.445164e-17, 8.437773e-17, 8.437524e-17, 
    8.437979e-17, 8.43859e-17, 8.439188e-17, 8.439967e-17, 8.440053e-17, 
    8.440195e-17, 8.440579e-17, 8.440896e-17, 8.44023e-17, 8.440977e-17, 
    8.438193e-17, 8.439658e-17, 8.43742e-17, 8.438079e-17, 8.438558e-17, 
    8.438359e-17, 8.439438e-17, 8.439688e-17, 8.440704e-17, 8.440185e-17, 
    8.443324e-17, 8.441931e-17, 8.445854e-17, 8.444746e-17, 8.437435e-17, 
    8.437778e-17, 8.438956e-17, 8.438396e-17, 8.440024e-17, 8.440421e-17, 
    8.440753e-17, 8.441161e-17, 8.441213e-17, 8.441456e-17, 8.441057e-17, 
    8.441444e-17, 8.439968e-17, 8.440629e-17, 8.438834e-17, 8.439263e-17, 
    8.439069e-17, 8.438848e-17, 8.439529e-17, 8.440238e-17, 8.44027e-17, 
    8.440495e-17, 8.441097e-17, 8.440032e-17, 8.443472e-17, 8.441313e-17, 
    8.43815e-17, 8.438787e-17, 8.438899e-17, 8.438648e-17, 8.440381e-17, 
    8.43975e-17, 8.441452e-17, 8.440996e-17, 8.441749e-17, 8.441373e-17, 
    8.441317e-17, 8.440838e-17, 8.440536e-17, 8.439775e-17, 8.439163e-17, 
    8.438687e-17, 8.438799e-17, 8.439323e-17, 8.440285e-17, 8.44121e-17, 
    8.441005e-17, 8.441692e-17, 8.439906e-17, 8.440645e-17, 8.440353e-17, 
    8.441117e-17, 8.439464e-17, 8.440818e-17, 8.439112e-17, 8.439265e-17, 
    8.439738e-17, 8.440683e-17, 8.440918e-17, 8.441139e-17, 8.441006e-17, 
    8.440313e-17, 8.440207e-17, 8.43973e-17, 8.43959e-17, 8.439233e-17, 
    8.438929e-17, 8.439202e-17, 8.439486e-17, 8.44032e-17, 8.441064e-17, 
    8.441882e-17, 8.44209e-17, 8.443004e-17, 8.442235e-17, 8.443481e-17, 
    8.442385e-17, 8.444301e-17, 8.440923e-17, 8.442389e-17, 8.439765e-17, 
    8.440051e-17, 8.44055e-17, 8.441735e-17, 8.441113e-17, 8.441849e-17, 
    8.440204e-17, 8.439332e-17, 8.439128e-17, 8.438713e-17, 8.439138e-17, 
    8.439104e-17, 8.43951e-17, 8.43938e-17, 8.440348e-17, 8.439829e-17, 
    8.441311e-17, 8.441848e-17, 8.44339e-17, 8.444328e-17, 8.445312e-17, 
    8.445738e-17, 8.445869e-17, 8.445923e-17 ;

 MEG_carene_3 =
  3.259777e-17, 3.260117e-17, 3.260052e-17, 3.260323e-17, 3.260176e-17, 
    3.260351e-17, 3.259848e-17, 3.260128e-17, 3.259951e-17, 3.259811e-17, 
    3.260842e-17, 3.260336e-17, 3.261397e-17, 3.261069e-17, 3.261903e-17, 
    3.261342e-17, 3.262017e-17, 3.261893e-17, 3.262283e-17, 3.262172e-17, 
    3.262657e-17, 3.262334e-17, 3.26292e-17, 3.262584e-17, 3.262634e-17, 
    3.262323e-17, 3.260444e-17, 3.260777e-17, 3.260423e-17, 3.260471e-17, 
    3.260451e-17, 3.260176e-17, 3.260033e-17, 3.259755e-17, 3.259807e-17, 
    3.260014e-17, 3.260493e-17, 3.260334e-17, 3.260746e-17, 3.260737e-17, 
    3.261192e-17, 3.260987e-17, 3.261758e-17, 3.26154e-17, 3.262177e-17, 
    3.262015e-17, 3.262168e-17, 3.262122e-17, 3.262168e-17, 3.261932e-17, 
    3.262033e-17, 3.261828e-17, 3.261024e-17, 3.261258e-17, 3.260558e-17, 
    3.260128e-17, 3.25986e-17, 3.259664e-17, 3.259691e-17, 3.259743e-17, 
    3.260015e-17, 3.260276e-17, 3.260474e-17, 3.260605e-17, 3.260736e-17, 
    3.261113e-17, 3.261328e-17, 3.261799e-17, 3.26172e-17, 3.261858e-17, 
    3.262e-17, 3.262229e-17, 3.262192e-17, 3.262291e-17, 3.261859e-17, 
    3.262144e-17, 3.261673e-17, 3.261801e-17, 3.260748e-17, 3.260378e-17, 
    3.260201e-17, 3.260064e-17, 3.259712e-17, 3.259954e-17, 3.259858e-17, 
    3.260091e-17, 3.260235e-17, 3.260165e-17, 3.260609e-17, 3.260435e-17, 
    3.261341e-17, 3.26095e-17, 3.261983e-17, 3.261736e-17, 3.262043e-17, 
    3.261887e-17, 3.262152e-17, 3.261914e-17, 3.262331e-17, 3.262419e-17, 
    3.262358e-17, 3.262599e-17, 3.2619e-17, 3.262166e-17, 3.260162e-17, 
    3.260173e-17, 3.260228e-17, 3.259984e-17, 3.25997e-17, 3.259752e-17, 
    3.259948e-17, 3.26003e-17, 3.260245e-17, 3.260369e-17, 3.260488e-17, 
    3.26075e-17, 3.26104e-17, 3.261452e-17, 3.261752e-17, 3.261953e-17, 
    3.261831e-17, 3.261938e-17, 3.261818e-17, 3.261762e-17, 3.262384e-17, 
    3.262033e-17, 3.262564e-17, 3.262536e-17, 3.262293e-17, 3.262539e-17, 
    3.260181e-17, 3.260115e-17, 3.259878e-17, 3.260064e-17, 3.259729e-17, 
    3.259914e-17, 3.260018e-17, 3.260434e-17, 3.260531e-17, 3.260614e-17, 
    3.260783e-17, 3.260997e-17, 3.261372e-17, 3.261703e-17, 3.262009e-17, 
    3.261987e-17, 3.261994e-17, 3.26206e-17, 3.261894e-17, 3.262088e-17, 
    3.262118e-17, 3.262035e-17, 3.262532e-17, 3.26239e-17, 3.262535e-17, 
    3.262443e-17, 3.260137e-17, 3.26025e-17, 3.260188e-17, 3.260302e-17, 
    3.26022e-17, 3.260578e-17, 3.260685e-17, 3.261195e-17, 3.260991e-17, 
    3.261322e-17, 3.261027e-17, 3.261078e-17, 3.261323e-17, 3.261044e-17, 
    3.26168e-17, 3.26124e-17, 3.262063e-17, 3.261614e-17, 3.26209e-17, 
    3.262007e-17, 3.262147e-17, 3.26227e-17, 3.262429e-17, 3.262717e-17, 
    3.262651e-17, 3.262895e-17, 3.260419e-17, 3.260563e-17, 3.260555e-17, 
    3.260709e-17, 3.260821e-17, 3.261072e-17, 3.261468e-17, 3.26132e-17, 
    3.261597e-17, 3.261651e-17, 3.261234e-17, 3.261485e-17, 3.260663e-17, 
    3.260791e-17, 3.260718e-17, 3.260428e-17, 3.261349e-17, 3.260873e-17, 
    3.261756e-17, 3.261499e-17, 3.262252e-17, 3.261873e-17, 3.262614e-17, 
    3.26292e-17, 3.26323e-17, 3.263568e-17, 3.260647e-17, 3.260548e-17, 
    3.260728e-17, 3.26097e-17, 3.261206e-17, 3.261514e-17, 3.261548e-17, 
    3.261604e-17, 3.261756e-17, 3.261881e-17, 3.261618e-17, 3.261913e-17, 
    3.260812e-17, 3.261392e-17, 3.260507e-17, 3.260767e-17, 3.260957e-17, 
    3.260878e-17, 3.261305e-17, 3.261404e-17, 3.261805e-17, 3.2616e-17, 
    3.262841e-17, 3.26229e-17, 3.263841e-17, 3.263403e-17, 3.260513e-17, 
    3.260648e-17, 3.261114e-17, 3.260893e-17, 3.261537e-17, 3.261694e-17, 
    3.261825e-17, 3.261986e-17, 3.262007e-17, 3.262103e-17, 3.261945e-17, 
    3.262098e-17, 3.261514e-17, 3.261776e-17, 3.261066e-17, 3.261236e-17, 
    3.261159e-17, 3.261072e-17, 3.261341e-17, 3.261621e-17, 3.261634e-17, 
    3.261722e-17, 3.261961e-17, 3.261539e-17, 3.262899e-17, 3.262046e-17, 
    3.260796e-17, 3.261047e-17, 3.261092e-17, 3.260993e-17, 3.261677e-17, 
    3.261428e-17, 3.262101e-17, 3.261921e-17, 3.262218e-17, 3.26207e-17, 
    3.262048e-17, 3.261858e-17, 3.261739e-17, 3.261438e-17, 3.261196e-17, 
    3.261008e-17, 3.261052e-17, 3.261259e-17, 3.26164e-17, 3.262005e-17, 
    3.261924e-17, 3.262196e-17, 3.26149e-17, 3.261782e-17, 3.261666e-17, 
    3.261969e-17, 3.261315e-17, 3.26185e-17, 3.261176e-17, 3.261236e-17, 
    3.261423e-17, 3.261797e-17, 3.26189e-17, 3.261977e-17, 3.261925e-17, 
    3.261651e-17, 3.261609e-17, 3.261421e-17, 3.261365e-17, 3.261224e-17, 
    3.261104e-17, 3.261212e-17, 3.261324e-17, 3.261654e-17, 3.261947e-17, 
    3.262271e-17, 3.262353e-17, 3.262715e-17, 3.262411e-17, 3.262903e-17, 
    3.26247e-17, 3.263227e-17, 3.261892e-17, 3.262471e-17, 3.261434e-17, 
    3.261547e-17, 3.261745e-17, 3.262213e-17, 3.261967e-17, 3.262258e-17, 
    3.261608e-17, 3.261263e-17, 3.261182e-17, 3.261018e-17, 3.261186e-17, 
    3.261173e-17, 3.261333e-17, 3.261282e-17, 3.261665e-17, 3.261459e-17, 
    3.262045e-17, 3.262257e-17, 3.262867e-17, 3.263237e-17, 3.263627e-17, 
    3.263795e-17, 3.263847e-17, 3.263868e-17 ;

 MEG_ethanol =
  1.676328e-18, 1.676591e-18, 1.676541e-18, 1.676751e-18, 1.676636e-18, 
    1.676772e-18, 1.676384e-18, 1.676599e-18, 1.676463e-18, 1.676355e-18, 
    1.677151e-18, 1.676761e-18, 1.67758e-18, 1.677327e-18, 1.677971e-18, 
    1.677538e-18, 1.67806e-18, 1.677964e-18, 1.678265e-18, 1.678179e-18, 
    1.678554e-18, 1.678305e-18, 1.678757e-18, 1.678497e-18, 1.678536e-18, 
    1.678296e-18, 1.676844e-18, 1.677101e-18, 1.676828e-18, 1.676865e-18, 
    1.676849e-18, 1.676637e-18, 1.676527e-18, 1.676311e-18, 1.676351e-18, 
    1.676511e-18, 1.676881e-18, 1.676759e-18, 1.677077e-18, 1.67707e-18, 
    1.677422e-18, 1.677263e-18, 1.677859e-18, 1.677691e-18, 1.678183e-18, 
    1.678058e-18, 1.678176e-18, 1.678141e-18, 1.678176e-18, 1.677994e-18, 
    1.678072e-18, 1.677913e-18, 1.677292e-18, 1.677473e-18, 1.676932e-18, 
    1.6766e-18, 1.676392e-18, 1.676241e-18, 1.676262e-18, 1.676302e-18, 
    1.676512e-18, 1.676714e-18, 1.676867e-18, 1.676968e-18, 1.677069e-18, 
    1.677361e-18, 1.677527e-18, 1.677891e-18, 1.67783e-18, 1.677937e-18, 
    1.678046e-18, 1.678223e-18, 1.678194e-18, 1.678271e-18, 1.677937e-18, 
    1.678158e-18, 1.677794e-18, 1.677893e-18, 1.677079e-18, 1.676793e-18, 
    1.676656e-18, 1.67655e-18, 1.676279e-18, 1.676465e-18, 1.676391e-18, 
    1.676571e-18, 1.676682e-18, 1.676628e-18, 1.676971e-18, 1.676837e-18, 
    1.677537e-18, 1.677235e-18, 1.678033e-18, 1.677843e-18, 1.678079e-18, 
    1.677959e-18, 1.678164e-18, 1.67798e-18, 1.678301e-18, 1.67837e-18, 
    1.678323e-18, 1.678509e-18, 1.677969e-18, 1.678174e-18, 1.676626e-18, 
    1.676634e-18, 1.676677e-18, 1.676488e-18, 1.676478e-18, 1.676309e-18, 
    1.676461e-18, 1.676524e-18, 1.67669e-18, 1.676786e-18, 1.676878e-18, 
    1.677081e-18, 1.677304e-18, 1.677623e-18, 1.677855e-18, 1.67801e-18, 
    1.677916e-18, 1.677998e-18, 1.677905e-18, 1.677862e-18, 1.678343e-18, 
    1.678071e-18, 1.678482e-18, 1.67846e-18, 1.678273e-18, 1.678462e-18, 
    1.676641e-18, 1.67659e-18, 1.676407e-18, 1.67655e-18, 1.676291e-18, 
    1.676434e-18, 1.676515e-18, 1.676836e-18, 1.676911e-18, 1.676975e-18, 
    1.677106e-18, 1.677271e-18, 1.677561e-18, 1.677817e-18, 1.678053e-18, 
    1.678036e-18, 1.678042e-18, 1.678093e-18, 1.677964e-18, 1.678114e-18, 
    1.678137e-18, 1.678073e-18, 1.678457e-18, 1.678347e-18, 1.678459e-18, 
    1.678389e-18, 1.676607e-18, 1.676694e-18, 1.676646e-18, 1.676734e-18, 
    1.676671e-18, 1.676948e-18, 1.677031e-18, 1.677424e-18, 1.677267e-18, 
    1.677522e-18, 1.677294e-18, 1.677334e-18, 1.677523e-18, 1.677308e-18, 
    1.677799e-18, 1.677459e-18, 1.678095e-18, 1.677748e-18, 1.678116e-18, 
    1.678052e-18, 1.67816e-18, 1.678255e-18, 1.678378e-18, 1.6786e-18, 
    1.678549e-18, 1.678738e-18, 1.676825e-18, 1.676936e-18, 1.67693e-18, 
    1.677048e-18, 1.677136e-18, 1.677329e-18, 1.677636e-18, 1.677521e-18, 
    1.677735e-18, 1.677777e-18, 1.677454e-18, 1.677649e-18, 1.677013e-18, 
    1.677112e-18, 1.677056e-18, 1.676832e-18, 1.677543e-18, 1.677176e-18, 
    1.677858e-18, 1.677659e-18, 1.678241e-18, 1.677948e-18, 1.67852e-18, 
    1.678757e-18, 1.678996e-18, 1.679258e-18, 1.677e-18, 1.676924e-18, 
    1.677064e-18, 1.67725e-18, 1.677433e-18, 1.677671e-18, 1.677697e-18, 
    1.67774e-18, 1.677858e-18, 1.677954e-18, 1.677751e-18, 1.677979e-18, 
    1.677129e-18, 1.677576e-18, 1.676893e-18, 1.677094e-18, 1.677241e-18, 
    1.67718e-18, 1.677509e-18, 1.677586e-18, 1.677896e-18, 1.677737e-18, 
    1.678696e-18, 1.67827e-18, 1.679468e-18, 1.67913e-18, 1.676897e-18, 
    1.677002e-18, 1.677362e-18, 1.677191e-18, 1.677688e-18, 1.677809e-18, 
    1.677911e-18, 1.678035e-18, 1.678051e-18, 1.678125e-18, 1.678003e-18, 
    1.678122e-18, 1.677671e-18, 1.677873e-18, 1.677324e-18, 1.677456e-18, 
    1.677396e-18, 1.677329e-18, 1.677537e-18, 1.677753e-18, 1.677763e-18, 
    1.677832e-18, 1.678016e-18, 1.67769e-18, 1.678741e-18, 1.678082e-18, 
    1.677116e-18, 1.67731e-18, 1.677344e-18, 1.677268e-18, 1.677797e-18, 
    1.677604e-18, 1.678124e-18, 1.677985e-18, 1.678215e-18, 1.6781e-18, 
    1.678083e-18, 1.677937e-18, 1.677844e-18, 1.677612e-18, 1.677425e-18, 
    1.67728e-18, 1.677314e-18, 1.677474e-18, 1.677768e-18, 1.67805e-18, 
    1.677988e-18, 1.678197e-18, 1.677652e-18, 1.677878e-18, 1.677789e-18, 
    1.678022e-18, 1.677517e-18, 1.677931e-18, 1.677409e-18, 1.677456e-18, 
    1.677601e-18, 1.677889e-18, 1.677961e-18, 1.678029e-18, 1.677988e-18, 
    1.677776e-18, 1.677744e-18, 1.677598e-18, 1.677556e-18, 1.677446e-18, 
    1.677354e-18, 1.677437e-18, 1.677524e-18, 1.677779e-18, 1.678006e-18, 
    1.678256e-18, 1.678319e-18, 1.678598e-18, 1.678364e-18, 1.678744e-18, 
    1.678409e-18, 1.678994e-18, 1.677963e-18, 1.67841e-18, 1.677609e-18, 
    1.677696e-18, 1.677849e-18, 1.678211e-18, 1.678021e-18, 1.678246e-18, 
    1.677743e-18, 1.677477e-18, 1.677414e-18, 1.677287e-18, 1.677417e-18, 
    1.677407e-18, 1.677531e-18, 1.677492e-18, 1.677787e-18, 1.677628e-18, 
    1.678081e-18, 1.678245e-18, 1.678716e-18, 1.679002e-18, 1.679303e-18, 
    1.679433e-18, 1.679473e-18, 1.679489e-18 ;

 MEG_formaldehyde =
  3.352656e-19, 3.353182e-19, 3.353082e-19, 3.353501e-19, 3.353273e-19, 
    3.353544e-19, 3.352767e-19, 3.353199e-19, 3.352926e-19, 3.352709e-19, 
    3.354303e-19, 3.353521e-19, 3.35516e-19, 3.354653e-19, 3.355942e-19, 
    3.355075e-19, 3.356119e-19, 3.355927e-19, 3.35653e-19, 3.356358e-19, 
    3.357108e-19, 3.356609e-19, 3.357514e-19, 3.356994e-19, 3.357071e-19, 
    3.356591e-19, 3.353688e-19, 3.354202e-19, 3.353655e-19, 3.353729e-19, 
    3.353698e-19, 3.353274e-19, 3.353053e-19, 3.352623e-19, 3.352703e-19, 
    3.353023e-19, 3.353763e-19, 3.353518e-19, 3.354155e-19, 3.354141e-19, 
    3.354844e-19, 3.354527e-19, 3.355718e-19, 3.355382e-19, 3.356365e-19, 
    3.356116e-19, 3.356352e-19, 3.356281e-19, 3.356353e-19, 3.355988e-19, 
    3.356143e-19, 3.355826e-19, 3.354584e-19, 3.354945e-19, 3.353864e-19, 
    3.353199e-19, 3.352784e-19, 3.352482e-19, 3.352525e-19, 3.352604e-19, 
    3.353024e-19, 3.353429e-19, 3.353734e-19, 3.353937e-19, 3.354138e-19, 
    3.354722e-19, 3.355054e-19, 3.355782e-19, 3.355659e-19, 3.355874e-19, 
    3.356091e-19, 3.356446e-19, 3.356388e-19, 3.356543e-19, 3.355874e-19, 
    3.356315e-19, 3.355587e-19, 3.355785e-19, 3.354158e-19, 3.353586e-19, 
    3.353312e-19, 3.3531e-19, 3.352557e-19, 3.35293e-19, 3.352782e-19, 
    3.353142e-19, 3.353365e-19, 3.353256e-19, 3.353943e-19, 3.353674e-19, 
    3.355074e-19, 3.35447e-19, 3.356066e-19, 3.355685e-19, 3.356159e-19, 
    3.355919e-19, 3.356327e-19, 3.35596e-19, 3.356603e-19, 3.356739e-19, 
    3.356645e-19, 3.357018e-19, 3.355938e-19, 3.356348e-19, 3.353251e-19, 
    3.353269e-19, 3.353355e-19, 3.352976e-19, 3.352955e-19, 3.352619e-19, 
    3.352921e-19, 3.353047e-19, 3.353381e-19, 3.353572e-19, 3.353756e-19, 
    3.354161e-19, 3.354608e-19, 3.355245e-19, 3.355709e-19, 3.356019e-19, 
    3.355831e-19, 3.355997e-19, 3.35581e-19, 3.355725e-19, 3.356686e-19, 
    3.356143e-19, 3.356964e-19, 3.35692e-19, 3.356545e-19, 3.356925e-19, 
    3.353282e-19, 3.353179e-19, 3.352813e-19, 3.3531e-19, 3.352583e-19, 
    3.352868e-19, 3.353029e-19, 3.353672e-19, 3.353822e-19, 3.35395e-19, 
    3.354211e-19, 3.354543e-19, 3.355122e-19, 3.355633e-19, 3.356106e-19, 
    3.356072e-19, 3.356083e-19, 3.356185e-19, 3.355928e-19, 3.356228e-19, 
    3.356275e-19, 3.356147e-19, 3.356913e-19, 3.356695e-19, 3.356919e-19, 
    3.356777e-19, 3.353213e-19, 3.353387e-19, 3.353293e-19, 3.353469e-19, 
    3.353342e-19, 3.353895e-19, 3.354061e-19, 3.354849e-19, 3.354534e-19, 
    3.355045e-19, 3.354589e-19, 3.354667e-19, 3.355047e-19, 3.354615e-19, 
    3.355599e-19, 3.354918e-19, 3.356189e-19, 3.355495e-19, 3.356232e-19, 
    3.356104e-19, 3.35632e-19, 3.35651e-19, 3.356756e-19, 3.3572e-19, 
    3.357098e-19, 3.357475e-19, 3.35365e-19, 3.353872e-19, 3.353859e-19, 
    3.354097e-19, 3.354271e-19, 3.354658e-19, 3.355271e-19, 3.355042e-19, 
    3.355469e-19, 3.355553e-19, 3.354908e-19, 3.355297e-19, 3.354026e-19, 
    3.354224e-19, 3.354111e-19, 3.353663e-19, 3.355086e-19, 3.354351e-19, 
    3.355716e-19, 3.355318e-19, 3.356482e-19, 3.355896e-19, 3.357041e-19, 
    3.357515e-19, 3.357992e-19, 3.358515e-19, 3.354001e-19, 3.353849e-19, 
    3.354127e-19, 3.3545e-19, 3.354865e-19, 3.355341e-19, 3.355393e-19, 
    3.355481e-19, 3.355715e-19, 3.355909e-19, 3.355502e-19, 3.355958e-19, 
    3.354257e-19, 3.355153e-19, 3.353785e-19, 3.354188e-19, 3.354481e-19, 
    3.354359e-19, 3.355018e-19, 3.355171e-19, 3.355792e-19, 3.355474e-19, 
    3.357392e-19, 3.356541e-19, 3.358936e-19, 3.35826e-19, 3.353794e-19, 
    3.354003e-19, 3.354723e-19, 3.354382e-19, 3.355376e-19, 3.355619e-19, 
    3.355822e-19, 3.356071e-19, 3.356102e-19, 3.356251e-19, 3.356007e-19, 
    3.356244e-19, 3.355342e-19, 3.355746e-19, 3.354649e-19, 3.354911e-19, 
    3.354793e-19, 3.354658e-19, 3.355074e-19, 3.355506e-19, 3.355526e-19, 
    3.355664e-19, 3.356031e-19, 3.355381e-19, 3.357482e-19, 3.356164e-19, 
    3.354231e-19, 3.35462e-19, 3.354689e-19, 3.354536e-19, 3.355594e-19, 
    3.355209e-19, 3.356249e-19, 3.355969e-19, 3.35643e-19, 3.3562e-19, 
    3.356166e-19, 3.355873e-19, 3.355689e-19, 3.355224e-19, 3.35485e-19, 
    3.354559e-19, 3.354628e-19, 3.354948e-19, 3.355535e-19, 3.3561e-19, 
    3.355975e-19, 3.356395e-19, 3.355304e-19, 3.355755e-19, 3.355577e-19, 
    3.356044e-19, 3.355034e-19, 3.355861e-19, 3.354819e-19, 3.354912e-19, 
    3.355201e-19, 3.355779e-19, 3.355922e-19, 3.356057e-19, 3.355976e-19, 
    3.355553e-19, 3.355488e-19, 3.355197e-19, 3.355111e-19, 3.354893e-19, 
    3.354707e-19, 3.354874e-19, 3.355047e-19, 3.355557e-19, 3.356011e-19, 
    3.356511e-19, 3.356638e-19, 3.357197e-19, 3.356727e-19, 3.357488e-19, 
    3.356819e-19, 3.357989e-19, 3.355925e-19, 3.35682e-19, 3.355218e-19, 
    3.355393e-19, 3.355698e-19, 3.356421e-19, 3.356042e-19, 3.356491e-19, 
    3.355486e-19, 3.354953e-19, 3.354829e-19, 3.354575e-19, 3.354835e-19, 
    3.354814e-19, 3.355062e-19, 3.354983e-19, 3.355574e-19, 3.355257e-19, 
    3.356162e-19, 3.35649e-19, 3.357432e-19, 3.358004e-19, 3.358605e-19, 
    3.358866e-19, 3.358946e-19, 3.358979e-19 ;

 MEG_isoprene =
  2.294623e-19, 2.295062e-19, 2.294979e-19, 2.295328e-19, 2.295137e-19, 
    2.295364e-19, 2.294716e-19, 2.295076e-19, 2.294848e-19, 2.294668e-19, 
    2.295996e-19, 2.295345e-19, 2.29671e-19, 2.296288e-19, 2.297361e-19, 
    2.296639e-19, 2.297509e-19, 2.297349e-19, 2.297851e-19, 2.297707e-19, 
    2.298332e-19, 2.297917e-19, 2.29867e-19, 2.298237e-19, 2.298302e-19, 
    2.297902e-19, 2.295484e-19, 2.295912e-19, 2.295456e-19, 2.295518e-19, 
    2.295492e-19, 2.295138e-19, 2.294954e-19, 2.294596e-19, 2.294662e-19, 
    2.294929e-19, 2.295546e-19, 2.295342e-19, 2.295872e-19, 2.295861e-19, 
    2.296447e-19, 2.296182e-19, 2.297175e-19, 2.296894e-19, 2.297713e-19, 
    2.297506e-19, 2.297702e-19, 2.297644e-19, 2.297703e-19, 2.297399e-19, 
    2.297529e-19, 2.297265e-19, 2.29623e-19, 2.296531e-19, 2.29563e-19, 
    2.295076e-19, 2.29473e-19, 2.294479e-19, 2.294514e-19, 2.29458e-19, 
    2.294931e-19, 2.295267e-19, 2.295522e-19, 2.295691e-19, 2.295859e-19, 
    2.296345e-19, 2.296622e-19, 2.297228e-19, 2.297126e-19, 2.297304e-19, 
    2.297486e-19, 2.297781e-19, 2.297733e-19, 2.297861e-19, 2.297305e-19, 
    2.297672e-19, 2.297066e-19, 2.29723e-19, 2.295875e-19, 2.295398e-19, 
    2.295171e-19, 2.294993e-19, 2.294541e-19, 2.294852e-19, 2.294729e-19, 
    2.295028e-19, 2.295214e-19, 2.295124e-19, 2.295696e-19, 2.295472e-19, 
    2.296638e-19, 2.296136e-19, 2.297465e-19, 2.297147e-19, 2.297542e-19, 
    2.297342e-19, 2.297682e-19, 2.297376e-19, 2.297911e-19, 2.298025e-19, 
    2.297947e-19, 2.298257e-19, 2.297358e-19, 2.297699e-19, 2.29512e-19, 
    2.295134e-19, 2.295206e-19, 2.29489e-19, 2.294873e-19, 2.294593e-19, 
    2.294844e-19, 2.294949e-19, 2.295227e-19, 2.295387e-19, 2.29554e-19, 
    2.295878e-19, 2.296251e-19, 2.296781e-19, 2.297167e-19, 2.297425e-19, 
    2.297269e-19, 2.297407e-19, 2.297252e-19, 2.29718e-19, 2.29798e-19, 
    2.297528e-19, 2.298212e-19, 2.298175e-19, 2.297863e-19, 2.298179e-19, 
    2.295145e-19, 2.29506e-19, 2.294755e-19, 2.294993e-19, 2.294562e-19, 
    2.2948e-19, 2.294935e-19, 2.29547e-19, 2.295595e-19, 2.295702e-19, 
    2.295919e-19, 2.296195e-19, 2.296679e-19, 2.297104e-19, 2.297498e-19, 
    2.297469e-19, 2.297479e-19, 2.297564e-19, 2.297349e-19, 2.297599e-19, 
    2.297638e-19, 2.297532e-19, 2.29817e-19, 2.297988e-19, 2.298175e-19, 
    2.298056e-19, 2.295088e-19, 2.295233e-19, 2.295154e-19, 2.295301e-19, 
    2.295195e-19, 2.295656e-19, 2.295795e-19, 2.296451e-19, 2.296188e-19, 
    2.296614e-19, 2.296234e-19, 2.2963e-19, 2.296616e-19, 2.296256e-19, 
    2.297075e-19, 2.296509e-19, 2.297567e-19, 2.296989e-19, 2.297603e-19, 
    2.297496e-19, 2.297676e-19, 2.297834e-19, 2.298039e-19, 2.298408e-19, 
    2.298324e-19, 2.298638e-19, 2.295452e-19, 2.295637e-19, 2.295626e-19, 
    2.295824e-19, 2.29597e-19, 2.296291e-19, 2.296802e-19, 2.296612e-19, 
    2.296968e-19, 2.297037e-19, 2.2965e-19, 2.296824e-19, 2.295765e-19, 
    2.295931e-19, 2.295836e-19, 2.295463e-19, 2.296648e-19, 2.296036e-19, 
    2.297173e-19, 2.296841e-19, 2.297811e-19, 2.297323e-19, 2.298276e-19, 
    2.298671e-19, 2.299068e-19, 2.299503e-19, 2.295744e-19, 2.295617e-19, 
    2.295849e-19, 2.29616e-19, 2.296464e-19, 2.296861e-19, 2.296904e-19, 
    2.296977e-19, 2.297172e-19, 2.297334e-19, 2.296995e-19, 2.297375e-19, 
    2.295958e-19, 2.296704e-19, 2.295565e-19, 2.2959e-19, 2.296144e-19, 
    2.296042e-19, 2.296591e-19, 2.296719e-19, 2.297236e-19, 2.296972e-19, 
    2.298568e-19, 2.29786e-19, 2.299853e-19, 2.299291e-19, 2.295572e-19, 
    2.295746e-19, 2.296346e-19, 2.296061e-19, 2.29689e-19, 2.297092e-19, 
    2.297261e-19, 2.297468e-19, 2.297495e-19, 2.297618e-19, 2.297415e-19, 
    2.297612e-19, 2.296861e-19, 2.297198e-19, 2.296284e-19, 2.296503e-19, 
    2.296404e-19, 2.296292e-19, 2.296638e-19, 2.296999e-19, 2.297015e-19, 
    2.297129e-19, 2.297436e-19, 2.296894e-19, 2.298644e-19, 2.297546e-19, 
    2.295936e-19, 2.29626e-19, 2.296317e-19, 2.29619e-19, 2.297071e-19, 
    2.29675e-19, 2.297616e-19, 2.297384e-19, 2.297767e-19, 2.297576e-19, 
    2.297547e-19, 2.297304e-19, 2.29715e-19, 2.296764e-19, 2.296452e-19, 
    2.296209e-19, 2.296267e-19, 2.296533e-19, 2.297023e-19, 2.297493e-19, 
    2.297389e-19, 2.297738e-19, 2.29683e-19, 2.297206e-19, 2.297057e-19, 
    2.297446e-19, 2.296605e-19, 2.297294e-19, 2.296426e-19, 2.296504e-19, 
    2.296744e-19, 2.297225e-19, 2.297345e-19, 2.297457e-19, 2.297389e-19, 
    2.297037e-19, 2.296983e-19, 2.29674e-19, 2.296669e-19, 2.296487e-19, 
    2.296333e-19, 2.296472e-19, 2.296616e-19, 2.29704e-19, 2.297419e-19, 
    2.297835e-19, 2.29794e-19, 2.298406e-19, 2.298015e-19, 2.298648e-19, 
    2.298091e-19, 2.299065e-19, 2.297347e-19, 2.298093e-19, 2.296758e-19, 
    2.296904e-19, 2.297158e-19, 2.29776e-19, 2.297444e-19, 2.297818e-19, 
    2.296982e-19, 2.296538e-19, 2.296434e-19, 2.296223e-19, 2.296439e-19, 
    2.296422e-19, 2.296628e-19, 2.296563e-19, 2.297055e-19, 2.296791e-19, 
    2.297544e-19, 2.297818e-19, 2.298602e-19, 2.299078e-19, 2.299578e-19, 
    2.299794e-19, 2.299861e-19, 2.299889e-19 ;

 MEG_methanol =
  5.798236e-17, 5.798805e-17, 5.798697e-17, 5.79915e-17, 5.798903e-17, 
    5.799197e-17, 5.798356e-17, 5.798823e-17, 5.798527e-17, 5.798294e-17, 
    5.800016e-17, 5.799171e-17, 5.800943e-17, 5.800395e-17, 5.801787e-17, 
    5.800851e-17, 5.801978e-17, 5.801771e-17, 5.802422e-17, 5.802236e-17, 
    5.803046e-17, 5.802508e-17, 5.803485e-17, 5.802923e-17, 5.803007e-17, 
    5.802488e-17, 5.799352e-17, 5.799907e-17, 5.799316e-17, 5.799396e-17, 
    5.799363e-17, 5.798904e-17, 5.798665e-17, 5.7982e-17, 5.798287e-17, 
    5.798633e-17, 5.799432e-17, 5.799168e-17, 5.799856e-17, 5.799841e-17, 
    5.800601e-17, 5.800258e-17, 5.801546e-17, 5.801182e-17, 5.802244e-17, 
    5.801975e-17, 5.802229e-17, 5.802154e-17, 5.802231e-17, 5.801837e-17, 
    5.802005e-17, 5.801662e-17, 5.80032e-17, 5.800711e-17, 5.799541e-17, 
    5.798823e-17, 5.798375e-17, 5.798048e-17, 5.798094e-17, 5.79818e-17, 
    5.798634e-17, 5.799071e-17, 5.799402e-17, 5.799621e-17, 5.799838e-17, 
    5.80047e-17, 5.800828e-17, 5.801614e-17, 5.801482e-17, 5.801713e-17, 
    5.801949e-17, 5.802331e-17, 5.80227e-17, 5.802436e-17, 5.801714e-17, 
    5.80219e-17, 5.801404e-17, 5.801618e-17, 5.79986e-17, 5.799241e-17, 
    5.798946e-17, 5.798716e-17, 5.798129e-17, 5.798532e-17, 5.798373e-17, 
    5.798761e-17, 5.799003e-17, 5.798885e-17, 5.799627e-17, 5.799337e-17, 
    5.80085e-17, 5.800198e-17, 5.801922e-17, 5.801509e-17, 5.802022e-17, 
    5.801762e-17, 5.802203e-17, 5.801806e-17, 5.802501e-17, 5.802648e-17, 
    5.802546e-17, 5.802949e-17, 5.801783e-17, 5.802226e-17, 5.79888e-17, 
    5.798899e-17, 5.798991e-17, 5.798582e-17, 5.798559e-17, 5.798196e-17, 
    5.798523e-17, 5.798659e-17, 5.79902e-17, 5.799226e-17, 5.799425e-17, 
    5.799863e-17, 5.800347e-17, 5.801035e-17, 5.801536e-17, 5.801871e-17, 
    5.801667e-17, 5.801846e-17, 5.801645e-17, 5.801552e-17, 5.802591e-17, 
    5.802004e-17, 5.802891e-17, 5.802843e-17, 5.802438e-17, 5.802849e-17, 
    5.798913e-17, 5.798802e-17, 5.798406e-17, 5.798716e-17, 5.798157e-17, 
    5.798465e-17, 5.798639e-17, 5.799335e-17, 5.799496e-17, 5.799635e-17, 
    5.799917e-17, 5.800275e-17, 5.800902e-17, 5.801454e-17, 5.801964e-17, 
    5.801928e-17, 5.80194e-17, 5.80205e-17, 5.801772e-17, 5.802096e-17, 
    5.802147e-17, 5.802008e-17, 5.802837e-17, 5.8026e-17, 5.802842e-17, 
    5.802689e-17, 5.798839e-17, 5.799026e-17, 5.798925e-17, 5.799114e-17, 
    5.798977e-17, 5.799576e-17, 5.799755e-17, 5.800606e-17, 5.800266e-17, 
    5.800818e-17, 5.800325e-17, 5.80041e-17, 5.80082e-17, 5.800354e-17, 
    5.801416e-17, 5.800681e-17, 5.802055e-17, 5.801304e-17, 5.8021e-17, 
    5.801962e-17, 5.802196e-17, 5.802401e-17, 5.802666e-17, 5.803145e-17, 
    5.803036e-17, 5.803443e-17, 5.79931e-17, 5.799551e-17, 5.799537e-17, 
    5.799793e-17, 5.799982e-17, 5.8004e-17, 5.801062e-17, 5.800815e-17, 
    5.801276e-17, 5.801367e-17, 5.80067e-17, 5.801091e-17, 5.799717e-17, 
    5.799932e-17, 5.799809e-17, 5.799325e-17, 5.800862e-17, 5.800069e-17, 
    5.801543e-17, 5.801113e-17, 5.80237e-17, 5.801737e-17, 5.802974e-17, 
    5.803485e-17, 5.804001e-17, 5.804565e-17, 5.79969e-17, 5.799525e-17, 
    5.799826e-17, 5.800229e-17, 5.800624e-17, 5.801138e-17, 5.801194e-17, 
    5.801289e-17, 5.801542e-17, 5.801752e-17, 5.801311e-17, 5.801804e-17, 
    5.799967e-17, 5.800935e-17, 5.799457e-17, 5.799892e-17, 5.800209e-17, 
    5.800077e-17, 5.800789e-17, 5.800954e-17, 5.801625e-17, 5.801282e-17, 
    5.803353e-17, 5.802434e-17, 5.80502e-17, 5.80429e-17, 5.799467e-17, 
    5.799693e-17, 5.80047e-17, 5.800101e-17, 5.801176e-17, 5.801438e-17, 
    5.801657e-17, 5.801926e-17, 5.801961e-17, 5.802121e-17, 5.801857e-17, 
    5.802113e-17, 5.801139e-17, 5.801575e-17, 5.80039e-17, 5.800674e-17, 
    5.800546e-17, 5.8004e-17, 5.800849e-17, 5.801317e-17, 5.801339e-17, 
    5.801486e-17, 5.801884e-17, 5.80118e-17, 5.80345e-17, 5.802027e-17, 
    5.799939e-17, 5.800359e-17, 5.800433e-17, 5.800268e-17, 5.801411e-17, 
    5.800995e-17, 5.802118e-17, 5.801817e-17, 5.802314e-17, 5.802066e-17, 
    5.802029e-17, 5.801713e-17, 5.801513e-17, 5.801012e-17, 5.800608e-17, 
    5.800293e-17, 5.800367e-17, 5.800713e-17, 5.801348e-17, 5.801958e-17, 
    5.801823e-17, 5.802276e-17, 5.801098e-17, 5.801585e-17, 5.801393e-17, 
    5.801897e-17, 5.800806e-17, 5.8017e-17, 5.800574e-17, 5.800675e-17, 
    5.800987e-17, 5.801611e-17, 5.801766e-17, 5.801911e-17, 5.801824e-17, 
    5.801366e-17, 5.801297e-17, 5.800982e-17, 5.80089e-17, 5.800654e-17, 
    5.800453e-17, 5.800634e-17, 5.800821e-17, 5.801372e-17, 5.801862e-17, 
    5.802402e-17, 5.802538e-17, 5.803142e-17, 5.802635e-17, 5.803456e-17, 
    5.802734e-17, 5.803997e-17, 5.801769e-17, 5.802736e-17, 5.801005e-17, 
    5.801194e-17, 5.801523e-17, 5.802305e-17, 5.801894e-17, 5.80238e-17, 
    5.801295e-17, 5.800719e-17, 5.800585e-17, 5.80031e-17, 5.800591e-17, 
    5.800569e-17, 5.800837e-17, 5.800751e-17, 5.80139e-17, 5.801047e-17, 
    5.802025e-17, 5.802379e-17, 5.803396e-17, 5.804014e-17, 5.804663e-17, 
    5.804944e-17, 5.80503e-17, 5.805066e-17 ;

 MEG_pinene_a =
  4.796219e-17, 4.796741e-17, 4.796642e-17, 4.797057e-17, 4.796831e-17, 
    4.7971e-17, 4.796329e-17, 4.796758e-17, 4.796487e-17, 4.796272e-17, 
    4.797852e-17, 4.797077e-17, 4.798702e-17, 4.798199e-17, 4.799477e-17, 
    4.798618e-17, 4.799653e-17, 4.799463e-17, 4.80006e-17, 4.799889e-17, 
    4.800633e-17, 4.800139e-17, 4.801036e-17, 4.800521e-17, 4.800597e-17, 
    4.800121e-17, 4.797243e-17, 4.797752e-17, 4.79721e-17, 4.797283e-17, 
    4.797253e-17, 4.796832e-17, 4.796613e-17, 4.796186e-17, 4.796265e-17, 
    4.796583e-17, 4.797316e-17, 4.797074e-17, 4.797705e-17, 4.797691e-17, 
    4.798388e-17, 4.798074e-17, 4.799256e-17, 4.798922e-17, 4.799896e-17, 
    4.79965e-17, 4.799883e-17, 4.799814e-17, 4.799884e-17, 4.799523e-17, 
    4.799677e-17, 4.799362e-17, 4.798131e-17, 4.798489e-17, 4.797416e-17, 
    4.796758e-17, 4.796346e-17, 4.796047e-17, 4.796089e-17, 4.796168e-17, 
    4.796584e-17, 4.796985e-17, 4.797288e-17, 4.797489e-17, 4.797689e-17, 
    4.798268e-17, 4.798597e-17, 4.799318e-17, 4.799197e-17, 4.799409e-17, 
    4.799626e-17, 4.799977e-17, 4.79992e-17, 4.800073e-17, 4.79941e-17, 
    4.799847e-17, 4.799125e-17, 4.799321e-17, 4.797708e-17, 4.797141e-17, 
    4.79687e-17, 4.79666e-17, 4.796121e-17, 4.796491e-17, 4.796344e-17, 
    4.796701e-17, 4.796922e-17, 4.796814e-17, 4.797495e-17, 4.797229e-17, 
    4.798616e-17, 4.798018e-17, 4.7996e-17, 4.799222e-17, 4.799692e-17, 
    4.799454e-17, 4.799859e-17, 4.799495e-17, 4.800132e-17, 4.800267e-17, 
    4.800174e-17, 4.800544e-17, 4.799474e-17, 4.79988e-17, 4.796809e-17, 
    4.796827e-17, 4.796912e-17, 4.796537e-17, 4.796516e-17, 4.796182e-17, 
    4.796482e-17, 4.796607e-17, 4.796938e-17, 4.797127e-17, 4.797309e-17, 
    4.797711e-17, 4.798155e-17, 4.798786e-17, 4.799246e-17, 4.799554e-17, 
    4.799367e-17, 4.799532e-17, 4.799347e-17, 4.799262e-17, 4.800214e-17, 
    4.799676e-17, 4.80049e-17, 4.800447e-17, 4.800075e-17, 4.800452e-17, 
    4.79684e-17, 4.796738e-17, 4.796375e-17, 4.796659e-17, 4.796147e-17, 
    4.796429e-17, 4.796589e-17, 4.797227e-17, 4.797375e-17, 4.797502e-17, 
    4.797761e-17, 4.79809e-17, 4.798664e-17, 4.799171e-17, 4.799639e-17, 
    4.799606e-17, 4.799617e-17, 4.799718e-17, 4.799463e-17, 4.799761e-17, 
    4.799807e-17, 4.79968e-17, 4.80044e-17, 4.800223e-17, 4.800446e-17, 
    4.800305e-17, 4.796772e-17, 4.796944e-17, 4.79685e-17, 4.797025e-17, 
    4.796899e-17, 4.797448e-17, 4.797612e-17, 4.798393e-17, 4.798081e-17, 
    4.798588e-17, 4.798135e-17, 4.798213e-17, 4.79859e-17, 4.798162e-17, 
    4.799136e-17, 4.798462e-17, 4.799722e-17, 4.799034e-17, 4.799765e-17, 
    4.799637e-17, 4.799852e-17, 4.80004e-17, 4.800284e-17, 4.800724e-17, 
    4.800623e-17, 4.800998e-17, 4.797205e-17, 4.797425e-17, 4.797412e-17, 
    4.797648e-17, 4.797821e-17, 4.798204e-17, 4.798812e-17, 4.798585e-17, 
    4.799009e-17, 4.799091e-17, 4.798452e-17, 4.798838e-17, 4.797578e-17, 
    4.797774e-17, 4.797662e-17, 4.797218e-17, 4.798628e-17, 4.7979e-17, 
    4.799253e-17, 4.798859e-17, 4.800013e-17, 4.799431e-17, 4.800567e-17, 
    4.801036e-17, 4.80151e-17, 4.802029e-17, 4.797553e-17, 4.797402e-17, 
    4.797678e-17, 4.798047e-17, 4.79841e-17, 4.798881e-17, 4.798933e-17, 
    4.79902e-17, 4.799252e-17, 4.799445e-17, 4.799041e-17, 4.799493e-17, 
    4.797807e-17, 4.798695e-17, 4.797339e-17, 4.797738e-17, 4.798028e-17, 
    4.797908e-17, 4.798561e-17, 4.798713e-17, 4.799328e-17, 4.799014e-17, 
    4.800915e-17, 4.800071e-17, 4.802446e-17, 4.801776e-17, 4.797348e-17, 
    4.797555e-17, 4.798269e-17, 4.79793e-17, 4.798916e-17, 4.799157e-17, 
    4.799358e-17, 4.799605e-17, 4.799636e-17, 4.799783e-17, 4.799541e-17, 
    4.799776e-17, 4.798882e-17, 4.799282e-17, 4.798195e-17, 4.798455e-17, 
    4.798338e-17, 4.798204e-17, 4.798616e-17, 4.799045e-17, 4.799065e-17, 
    4.799201e-17, 4.799566e-17, 4.79892e-17, 4.801004e-17, 4.799697e-17, 
    4.797781e-17, 4.798167e-17, 4.798235e-17, 4.798083e-17, 4.799132e-17, 
    4.79875e-17, 4.799781e-17, 4.799504e-17, 4.799961e-17, 4.799733e-17, 
    4.799699e-17, 4.799409e-17, 4.799226e-17, 4.798766e-17, 4.798395e-17, 
    4.798106e-17, 4.798174e-17, 4.798491e-17, 4.799074e-17, 4.799634e-17, 
    4.79951e-17, 4.799926e-17, 4.798844e-17, 4.799292e-17, 4.799115e-17, 
    4.799578e-17, 4.798577e-17, 4.799397e-17, 4.798364e-17, 4.798457e-17, 
    4.798743e-17, 4.799315e-17, 4.799458e-17, 4.799591e-17, 4.799511e-17, 
    4.799091e-17, 4.799027e-17, 4.798738e-17, 4.798653e-17, 4.798437e-17, 
    4.798253e-17, 4.798418e-17, 4.79859e-17, 4.799095e-17, 4.799546e-17, 
    4.800041e-17, 4.800167e-17, 4.800721e-17, 4.800255e-17, 4.801009e-17, 
    4.800346e-17, 4.801506e-17, 4.79946e-17, 4.800348e-17, 4.798759e-17, 
    4.798933e-17, 4.799235e-17, 4.799952e-17, 4.799576e-17, 4.800022e-17, 
    4.799025e-17, 4.798497e-17, 4.798373e-17, 4.798122e-17, 4.798379e-17, 
    4.798359e-17, 4.798605e-17, 4.798526e-17, 4.799112e-17, 4.798798e-17, 
    4.799695e-17, 4.800021e-17, 4.800955e-17, 4.801522e-17, 4.802118e-17, 
    4.802376e-17, 4.802455e-17, 4.802488e-17 ;

 MEG_thujene_a =
  1.210192e-18, 1.210318e-18, 1.210294e-18, 1.210395e-18, 1.21034e-18, 
    1.210405e-18, 1.210219e-18, 1.210322e-18, 1.210257e-18, 1.210205e-18, 
    1.210588e-18, 1.2104e-18, 1.210793e-18, 1.210672e-18, 1.210981e-18, 
    1.210773e-18, 1.211024e-18, 1.210978e-18, 1.211123e-18, 1.211081e-18, 
    1.211261e-18, 1.211142e-18, 1.211359e-18, 1.211234e-18, 1.211253e-18, 
    1.211137e-18, 1.21044e-18, 1.210563e-18, 1.210432e-18, 1.21045e-18, 
    1.210442e-18, 1.21034e-18, 1.210287e-18, 1.210184e-18, 1.210203e-18, 
    1.21028e-18, 1.210458e-18, 1.210399e-18, 1.210552e-18, 1.210549e-18, 
    1.210718e-18, 1.210641e-18, 1.210928e-18, 1.210847e-18, 1.211083e-18, 
    1.211023e-18, 1.21108e-18, 1.211063e-18, 1.21108e-18, 1.210992e-18, 
    1.21103e-18, 1.210954e-18, 1.210655e-18, 1.210742e-18, 1.210482e-18, 
    1.210323e-18, 1.210223e-18, 1.21015e-18, 1.21016e-18, 1.21018e-18, 
    1.210281e-18, 1.210378e-18, 1.210451e-18, 1.2105e-18, 1.210548e-18, 
    1.210688e-18, 1.210768e-18, 1.210943e-18, 1.210913e-18, 1.210965e-18, 
    1.211017e-18, 1.211102e-18, 1.211089e-18, 1.211126e-18, 1.210965e-18, 
    1.211071e-18, 1.210896e-18, 1.210944e-18, 1.210553e-18, 1.210415e-18, 
    1.21035e-18, 1.210299e-18, 1.210168e-18, 1.210258e-18, 1.210222e-18, 
    1.210309e-18, 1.210362e-18, 1.210336e-18, 1.210501e-18, 1.210437e-18, 
    1.210773e-18, 1.210628e-18, 1.211011e-18, 1.21092e-18, 1.211033e-18, 
    1.210976e-18, 1.211074e-18, 1.210986e-18, 1.21114e-18, 1.211173e-18, 
    1.21115e-18, 1.21124e-18, 1.210981e-18, 1.211079e-18, 1.210335e-18, 
    1.210339e-18, 1.21036e-18, 1.210269e-18, 1.210264e-18, 1.210183e-18, 
    1.210256e-18, 1.210286e-18, 1.210366e-18, 1.210412e-18, 1.210456e-18, 
    1.210553e-18, 1.210661e-18, 1.210814e-18, 1.210925e-18, 1.211e-18, 
    1.210955e-18, 1.210995e-18, 1.21095e-18, 1.210929e-18, 1.21116e-18, 
    1.21103e-18, 1.211227e-18, 1.211216e-18, 1.211126e-18, 1.211218e-18, 
    1.210342e-18, 1.210318e-18, 1.21023e-18, 1.210299e-18, 1.210174e-18, 
    1.210243e-18, 1.210282e-18, 1.210436e-18, 1.210472e-18, 1.210503e-18, 
    1.210566e-18, 1.210645e-18, 1.210784e-18, 1.210907e-18, 1.211021e-18, 
    1.211013e-18, 1.211015e-18, 1.21104e-18, 1.210978e-18, 1.21105e-18, 
    1.211061e-18, 1.211031e-18, 1.211215e-18, 1.211162e-18, 1.211216e-18, 
    1.211182e-18, 1.210326e-18, 1.210368e-18, 1.210345e-18, 1.210387e-18, 
    1.210357e-18, 1.21049e-18, 1.21053e-18, 1.210719e-18, 1.210643e-18, 
    1.210766e-18, 1.210656e-18, 1.210675e-18, 1.210766e-18, 1.210663e-18, 
    1.210899e-18, 1.210735e-18, 1.211041e-18, 1.210874e-18, 1.211051e-18, 
    1.21102e-18, 1.211072e-18, 1.211118e-18, 1.211177e-18, 1.211283e-18, 
    1.211259e-18, 1.21135e-18, 1.210431e-18, 1.210484e-18, 1.210481e-18, 
    1.210538e-18, 1.21058e-18, 1.210673e-18, 1.21082e-18, 1.210765e-18, 
    1.210868e-18, 1.210888e-18, 1.210733e-18, 1.210827e-18, 1.210521e-18, 
    1.210569e-18, 1.210542e-18, 1.210434e-18, 1.210776e-18, 1.210599e-18, 
    1.210927e-18, 1.210831e-18, 1.211111e-18, 1.21097e-18, 1.211245e-18, 
    1.211359e-18, 1.211474e-18, 1.2116e-18, 1.210515e-18, 1.210479e-18, 
    1.210545e-18, 1.210635e-18, 1.210723e-18, 1.210837e-18, 1.21085e-18, 
    1.210871e-18, 1.210927e-18, 1.210973e-18, 1.210876e-18, 1.210985e-18, 
    1.210577e-18, 1.210792e-18, 1.210463e-18, 1.21056e-18, 1.21063e-18, 
    1.210601e-18, 1.210759e-18, 1.210796e-18, 1.210945e-18, 1.210869e-18, 
    1.21133e-18, 1.211125e-18, 1.211701e-18, 1.211538e-18, 1.210465e-18, 
    1.210516e-18, 1.210689e-18, 1.210607e-18, 1.210845e-18, 1.210904e-18, 
    1.210953e-18, 1.211012e-18, 1.21102e-18, 1.211056e-18, 1.210997e-18, 
    1.211054e-18, 1.210837e-18, 1.210934e-18, 1.210671e-18, 1.210734e-18, 
    1.210705e-18, 1.210673e-18, 1.210773e-18, 1.210877e-18, 1.210882e-18, 
    1.210914e-18, 1.211003e-18, 1.210847e-18, 1.211351e-18, 1.211035e-18, 
    1.21057e-18, 1.210664e-18, 1.21068e-18, 1.210644e-18, 1.210898e-18, 
    1.210805e-18, 1.211055e-18, 1.210988e-18, 1.211099e-18, 1.211043e-18, 
    1.211035e-18, 1.210965e-18, 1.210921e-18, 1.210809e-18, 1.210719e-18, 
    1.210649e-18, 1.210666e-18, 1.210743e-18, 1.210884e-18, 1.211019e-18, 
    1.210989e-18, 1.21109e-18, 1.210828e-18, 1.210936e-18, 1.210894e-18, 
    1.211006e-18, 1.210763e-18, 1.210962e-18, 1.210712e-18, 1.210734e-18, 
    1.210803e-18, 1.210942e-18, 1.210977e-18, 1.211009e-18, 1.21099e-18, 
    1.210888e-18, 1.210872e-18, 1.210802e-18, 1.210782e-18, 1.210729e-18, 
    1.210685e-18, 1.210725e-18, 1.210766e-18, 1.210889e-18, 1.210998e-18, 
    1.211118e-18, 1.211149e-18, 1.211283e-18, 1.21117e-18, 1.211353e-18, 
    1.211192e-18, 1.211473e-18, 1.210977e-18, 1.211192e-18, 1.210807e-18, 
    1.210849e-18, 1.210923e-18, 1.211097e-18, 1.211005e-18, 1.211113e-18, 
    1.210872e-18, 1.210744e-18, 1.210714e-18, 1.210653e-18, 1.210715e-18, 
    1.21071e-18, 1.21077e-18, 1.210751e-18, 1.210893e-18, 1.210817e-18, 
    1.211034e-18, 1.211113e-18, 1.211339e-18, 1.211477e-18, 1.211621e-18, 
    1.211684e-18, 1.211703e-18, 1.211711e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -2.3075e-25, -1.510863e-25, 3.049198e-25, -1.730625e-25, 1.867978e-25, 
    4.66995e-26, -9.065174e-26, -3.296421e-26, 1.208692e-25, 2.389912e-25, 
    -4.367769e-25, 5.219355e-26, -1.813036e-25, -3.40631e-25, 3.021735e-26, 
    2.527264e-25, -8.240992e-27, -1.730625e-25, -7.966364e-26, -3.323899e-25, 
    1.455924e-25, 4.120545e-26, -2.032798e-25, 2.747033e-26, -4.312828e-25, 
    1.648223e-26, 3.21402e-25, -6.647799e-25, -1.648207e-26, 1.758097e-25, 
    2.14268e-25, 2.911847e-25, -7.197204e-25, 2.554734e-25, 4.120545e-26, 
    2.472323e-25, 1.538335e-25, -2.747024e-25, -4.999584e-25, 4.395241e-25, 
    -1.730625e-25, -2.911845e-25, 8.241083e-26, 6.015985e-25, -6.318148e-26, 
    -4.642471e-25, -8.241066e-26, 5.76876e-26, -3.681012e-25, -2.417381e-25, 
    -2.746942e-27, -1.950387e-25, 7.087325e-25, -2.417381e-25, -3.708483e-25, 
    8.515785e-26, -1.098802e-26, -4.038125e-25, -4.53259e-25, 2.032799e-25, 
    1.648223e-26, -2.884375e-25, -2.994256e-25, 3.516192e-25, -2.25256e-25, 
    -1.895446e-25, -1.291101e-25, -2.28003e-25, 4.395248e-26, -3.076667e-25, 
    2.14268e-25, -3.021719e-26, 1.126281e-25, -3.46125e-25, 4.202949e-25, 
    1.648216e-25, -2.060268e-25, -2.747016e-26, -3.626072e-25, -2.36244e-25, 
    -3.021719e-26, -4.340298e-25, -5.493967e-27, 4.175478e-25, 8.515785e-26, 
    7.96638e-26, 6.318165e-26, 4.532592e-25, -3.653542e-25, 1.153751e-25, 
    -3.735953e-25, -1.620744e-25, 1.895448e-25, 2.225091e-25, 3.323901e-25, 
    3.296438e-26, -5.081995e-25, 5.494132e-27, -1.895446e-25, 2.334972e-25, 
    3.296438e-26, 2.499793e-25, -2.417381e-25, -1.373512e-25, 4.28536e-25, 
    -4.148007e-25, -2.417381e-25, -5.494041e-26, -1.23616e-25, 1.455924e-25, 
    1.208692e-25, -2.856905e-25, -2.032798e-25, -1.565803e-25, -3.351369e-25, 
    1.126281e-25, -3.845826e-26, 3.708484e-25, 2.197628e-26, 9.339892e-26, 
    -3.845834e-25, -3.159078e-25, -6.318148e-26, -5.109465e-25, 
    -1.895446e-25, -2.582203e-25, 8.241083e-26, 2.032799e-25, -4.834763e-25, 
    2.994258e-25, -1.455922e-25, 2.389912e-25, 3.296438e-26, -1.922909e-26, 
    9.06519e-26, -1.950387e-25, -8.241066e-26, 1.922926e-26, -3.214018e-25, 
    4.395248e-26, -6.78515e-25, 1.922918e-25, 2.747026e-25, -1.098809e-25, 
    8.790487e-26, -2.225089e-25, -2.3075e-25, -1.538333e-25, 1.703156e-25, 
    -1.373504e-26, -1.15375e-25, -1.016398e-25, -2.884375e-25, 3.571133e-25, 
    -2.032798e-25, -1.620744e-25, -7.691661e-26, -1.455922e-25, 5.494058e-26, 
    8.241157e-27, 5.796223e-25, -5.493967e-27, 3.57114e-26, -1.098809e-25, 
    2.08774e-25, -5.246816e-25, 7.96638e-26, -2.389911e-25, -3.790893e-25, 
    3.18655e-25, -1.565803e-25, -1.538333e-25, -1.950387e-25, 4.175478e-25, 
    -3.845834e-25, -1.455922e-25, -6.592851e-26, 7.801551e-25, -9.614578e-26, 
    1.483394e-25, -1.703155e-25, 2.609674e-25, -2.637143e-25, -4.148007e-25, 
    -1.510863e-25, -5.521519e-25, 1.373521e-26, 5.494132e-27, -1.703155e-25, 
    -1.346041e-25, -2.801964e-25, 1.236162e-25, -1.18122e-25, -4.395239e-25, 
    2.14268e-25, 2.966788e-25, -2.664613e-25, 1.318573e-25, 7.416975e-26, 
    -8.515768e-26, 3.104139e-25, 8.241083e-26, -2.142679e-25, 1.04387e-25, 
    -2.554732e-25, -2.582203e-25, 2.08774e-25, -1.18122e-25, -1.593274e-25, 
    1.977859e-25, -3.900774e-25, -4.038125e-25, -1.071339e-25, 1.04387e-25, 
    8.25756e-32, 4.395248e-26, 3.378841e-25, 3.24149e-25, 3.57114e-26, 
    -1.675684e-25, -8.240992e-27, 1.620745e-25, 7.691677e-26, -4.889703e-25, 
    3.433782e-25, 1.648223e-26, -3.049197e-25, -2.747016e-26, -1.373512e-25, 
    -1.648207e-26, -3.296421e-26, -3.076667e-25, 6.043463e-26, 3.57114e-26, 
    8.241083e-26, -1.950387e-25, -3.021727e-25, -2.25256e-25, -7.142256e-26, 
    2.389912e-25, 5.494132e-27, 1.730626e-25, 1.703156e-25, 1.208692e-25, 
    -1.098809e-25, -5.329227e-25, -1.263631e-25, -1.977857e-25, 
    -3.543661e-25, 4.065598e-25, -3.708483e-25, 3.57114e-26, -3.983185e-25, 
    6.86757e-26, -8.240992e-27, 3.049198e-25, -2.25256e-25, -2.472321e-25, 
    -4.175477e-25, -1.895446e-25, 2.197628e-26, -8.240992e-27, -2.664613e-25, 
    3.735955e-25, 3.461252e-25, 2.747033e-26, -3.076667e-25, 5.494058e-26, 
    3.076668e-25, 4.944653e-26, 1.510864e-25, -1.703155e-25, 5.494132e-27, 
    -3.516191e-25, 2.032799e-25, -1.098802e-26, -4.615001e-25, 1.263632e-25, 
    -2.637143e-25, 8.790487e-26, 4.889705e-25, -7.416958e-26, -4.093066e-25, 
    -3.268959e-25, 1.620745e-25, -3.104137e-25, -1.593274e-25, -1.126279e-25, 
    -1.895446e-25, -1.23616e-25, 1.291103e-25, -6.318148e-26, 2.966788e-25, 
    -2.3075e-25, -4.53259e-25, -1.346041e-25, -1.291101e-25, -4.615001e-25, 
    9.06519e-26, 1.977859e-25, 2.197621e-25, 2.554734e-25, -1.867976e-25, 
    -5.851162e-25, 8.241157e-27, -3.928245e-25, -1.23616e-25, -3.626072e-25, 
    2.08774e-25, -2.499792e-25, 2.307502e-25, -7.966364e-26, -2.746942e-27, 
    -5.768744e-26, -3.955715e-25, -6.318148e-26, -4.999584e-25, 2.747107e-27, 
    2.856907e-25, -9.614578e-26, 1.208692e-25, -3.708483e-25, -2.389911e-25, 
    -2.911845e-25, -5.356697e-25, -6.592851e-26, -2.609673e-25, 1.318573e-25, 
    -1.648214e-25, 2.692085e-25, 1.0164e-25, -7.966364e-26, 2.472331e-26, 
    5.76876e-26, -1.565803e-25, 5.301759e-25, -2.197619e-25, -2.801964e-25 ;

 M_LITR2C_TO_LEACHING =
  -1.098805e-26, 3.3239e-25, 1.07134e-25, -1.648214e-25, -6.867557e-26, 
    1.703156e-25, -1.867976e-25, -1.373507e-26, -1.15375e-25, 9.614592e-26, 
    -2.170149e-25, -2.472322e-25, 1.153751e-25, 2.74703e-26, -9.614581e-26, 
    -1.098805e-26, -2.197614e-26, 1.64822e-26, 2.747078e-27, -2.197619e-25, 
    1.922918e-25, 5.219352e-26, -4.944639e-26, -5.494044e-26, 9.889295e-26, 
    -6.867557e-26, 1.922923e-26, -1.346042e-25, -1.043869e-25, 3.84584e-26, 
    7.691675e-26, -1.428452e-25, -2.554732e-25, -1.016399e-25, 2.472323e-25, 
    5.494055e-26, -1.318571e-25, -2.994256e-25, -2.884375e-25, 7.14227e-26, 
    3.076668e-25, -8.241069e-26, -1.510863e-25, 1.098815e-26, 5.219352e-26, 
    -3.35137e-25, 1.126281e-25, -1.455923e-25, -4.944639e-26, 1.09881e-25, 
    1.098815e-26, 2.472328e-26, -1.043869e-25, 2.801966e-25, 2.19762e-25, 
    2.252561e-25, -2.747024e-25, 4.669947e-26, -7.142259e-26, -1.15375e-25, 
    -2.472322e-25, 8.515782e-26, 8.515782e-26, -3.021722e-26, -1.620744e-25, 
    -8.790474e-26, -3.461251e-25, -1.098805e-26, -2.939316e-25, 
    -1.510863e-25, 1.208691e-25, 1.153751e-25, -3.186548e-25, -2.719554e-25, 
    3.021733e-26, 6.04346e-26, -2.527262e-25, -4.944639e-26, 1.703156e-25, 
    7.966377e-26, -1.785566e-25, 2.527263e-25, -1.922917e-25, -9.339879e-26, 
    1.126281e-25, 2.637144e-25, 8.790485e-26, -2.719554e-25, -3.076667e-25, 
    -1.703155e-25, -3.021722e-26, 9.339889e-26, -1.373512e-25, 2.74703e-26, 
    4.120543e-26, -2.499792e-25, -1.648214e-25, -1.538333e-25, 2.197625e-26, 
    -3.461251e-25, 2.472328e-26, -1.922917e-25, -2.225089e-25, -4.395234e-26, 
    1.455924e-25, -1.318571e-25, -2.25256e-25, -2.801965e-25, -3.296424e-26, 
    2.389912e-25, 1.153751e-25, -2.746971e-27, 6.04346e-26, -1.895447e-25, 
    3.131609e-25, 9.889295e-26, 1.098815e-26, -4.615001e-25, 5.35145e-32, 
    2.197625e-26, 7.416973e-26, 1.703156e-25, 2.74703e-26, -1.043869e-25, 
    3.3239e-25, 1.098815e-26, 1.895448e-25, 8.515782e-26, 1.373518e-26, 
    -1.043869e-25, 1.977858e-25, -2.472317e-26, 1.593275e-25, -1.236161e-25, 
    6.592865e-26, 8.790485e-26, -6.043449e-26, 3.84584e-26, -5.494044e-26, 
    2.362442e-25, -1.373512e-25, -1.016399e-25, 7.14227e-26, -1.071339e-25, 
    6.04346e-26, -1.922912e-26, 1.813037e-25, -1.236161e-25, -9.065177e-26, 
    -1.758095e-25, 7.14227e-26, -2.28003e-25, -5.60393e-25, 1.758096e-25, 
    -1.510863e-25, 1.09881e-25, 1.04387e-25, -1.813036e-25, 3.296435e-26, 
    -4.120532e-26, 7.14227e-26, -6.043449e-26, 3.296435e-26, -2.74702e-26, 
    6.592865e-26, 4.395245e-26, 9.339889e-26, 1.373513e-25, 1.263632e-25, 
    -1.043869e-25, 2.747078e-27, 3.021733e-26, 9.339889e-26, -1.15375e-25, 
    -1.922912e-26, 2.747078e-27, 2.884376e-25, 1.04387e-25, 4.120543e-26, 
    -1.785566e-25, 1.09881e-25, -5.493996e-27, 1.758096e-25, -5.494044e-26, 
    -6.043449e-26, -2.060268e-25, 9.889295e-26, -5.219346e-25, -3.131608e-25, 
    9.614592e-26, 9.614592e-26, -1.565804e-25, 2.197625e-26, -1.565804e-25, 
    -1.977857e-25, 3.049198e-25, -2.747024e-25, -1.455923e-25, -4.697412e-25, 
    1.428453e-25, 1.373518e-26, 1.09881e-25, 1.400983e-25, 3.296435e-26, 
    1.950388e-25, -1.318571e-25, 7.14227e-26, -1.071339e-25, 5.494103e-27, 
    -1.593274e-25, 6.592865e-26, -6.043449e-26, -5.493996e-27, -2.664613e-25, 
    -1.867976e-25, 1.400983e-25, 3.571138e-26, -2.582203e-25, -6.318152e-26, 
    -1.428452e-25, -1.318571e-25, -1.098809e-25, 1.09881e-25, 2.17015e-25, 
    -1.373512e-25, -3.296424e-26, -3.571127e-26, -3.186548e-25, 
    -3.571127e-26, -2.499792e-25, 3.21402e-25, -8.241069e-26, -1.593274e-25, 
    1.098815e-26, -7.691664e-26, -3.571127e-26, 4.395245e-26, -8.241069e-26, 
    7.14227e-26, -1.895447e-25, -2.472322e-25, 6.867567e-26, 7.14227e-26, 
    -2.060268e-25, -2.74702e-26, -5.494044e-26, -2.472317e-26, 1.758096e-25, 
    1.867977e-25, 2.11521e-25, 9.339889e-26, -2.994256e-25, -3.845829e-26, 
    2.197625e-26, -1.236161e-25, -6.318152e-26, -8.515771e-26, -3.571127e-26, 
    -7.416961e-26, 5.351445e-32, -2.197619e-25, -2.005328e-25, 5.494103e-27, 
    -2.746971e-27, -4.395234e-26, -7.691664e-26, -1.071339e-25, -1.15375e-25, 
    -1.373507e-26, -1.236161e-25, -1.263631e-25, -1.565804e-25, 2.74703e-26, 
    2.74703e-26, -9.065177e-26, -1.648209e-26, 1.758096e-25, 4.148008e-25, 
    -1.098809e-25, -1.620744e-25, -7.966367e-26, -4.395234e-26, 
    -3.516191e-25, -1.346042e-25, -1.867976e-25, -1.098809e-25, 
    -1.428452e-25, 1.620745e-25, 1.263632e-25, 1.703156e-25, -2.28003e-25, 
    -2.554732e-25, 5.351447e-32, 2.032799e-25, -6.318152e-26, -9.889284e-26, 
    2.197625e-26, 4.94465e-26, 3.84584e-26, 5.494055e-26, -2.087738e-25, 
    -2.829435e-25, -3.268959e-25, -1.373512e-25, -1.593274e-25, 1.291102e-25, 
    -3.021727e-25, 1.922923e-26, -1.098809e-25, 9.065187e-26, -3.845829e-26, 
    1.64822e-26, -1.483393e-25, 7.691675e-26, -1.977857e-25, -9.889284e-26, 
    5.494055e-26, -1.813036e-25, -5.493996e-27, -8.241069e-26, -6.592854e-26, 
    -8.241069e-26, 8.515782e-26, -1.538333e-25, 6.592865e-26, 1.620745e-25, 
    -2.801965e-25, -1.510863e-25, 1.922923e-26, 8.790485e-26, 1.758096e-25, 
    -1.593274e-25, -2.939316e-25, 2.032799e-25, 4.94465e-26, 2.252561e-25, 
    -1.785566e-25, -1.538333e-25 ;

 M_LITR3C_TO_LEACHING =
  7.691672e-26, 1.153751e-25, -1.09881e-25, -2.060266e-26, -1.922915e-26, 
    -1.922915e-26, -1.648212e-26, 4.944647e-26, -2.747022e-26, -6.043452e-26, 
    4.120564e-27, 2.747028e-26, -1.922915e-26, -1.346042e-25, -9.889287e-26, 
    -2.28003e-25, -1.12628e-25, -3.021725e-26, -6.180803e-26, 5.768755e-26, 
    -2.747022e-26, 1.648217e-26, 2.747052e-27, -6.043452e-26, -5.494023e-27, 
    8.653131e-26, 6.592862e-26, -2.060266e-26, -3.708481e-26, -1.346042e-25, 
    -5.081993e-26, 7.279618e-26, -2.197617e-26, -4.395237e-26, 1.675685e-25, 
    -5.494047e-26, -1.922917e-25, 1.373515e-26, 6.180808e-26, 5.21935e-26, 
    1.373539e-27, -5.219344e-26, -1.236161e-25, -3.159076e-26, 1.552069e-25, 
    -4.120511e-27, -8.241071e-26, -7.691667e-26, -1.922915e-26, 
    -4.944642e-26, -1.469658e-25, 4.395242e-26, -5.494047e-26, -8.241047e-27, 
    1.208691e-25, 1.277367e-25, 3.845837e-26, 4.669945e-26, -9.065179e-26, 
    5.494052e-26, -6.867535e-27, -7.279613e-26, 2.747052e-27, 3.02173e-26, 
    -1.373486e-27, 6.180808e-26, -7.142262e-26, 2.884379e-26, 1.181221e-25, 
    6.867565e-26, 1.593275e-25, 6.455511e-26, -4.669939e-26, 2.67572e-32, 
    -8.10372e-26, -1.043869e-25, 9.889292e-26, -3.57113e-26, 6.867589e-27, 
    -3.433778e-26, -6.318154e-26, -2.197617e-26, -2.334968e-26, 6.180808e-26, 
    4.395242e-26, 4.944647e-26, 8.653131e-26, -2.884373e-26, -4.120511e-27, 
    -6.180803e-26, 7.142267e-26, 5.906106e-26, -6.043452e-26, -2.47232e-26, 
    7.966375e-26, 1.66195e-25, 7.142267e-26, -5.494047e-26, -2.746998e-27, 
    -7.142262e-26, -5.768749e-26, -7.829018e-26, -2.746998e-27, 
    -2.486057e-25, -1.346042e-25, -2.747022e-26, -6.867559e-26, -1.15375e-25, 
    -7.966369e-26, 1.04387e-25, -7.966369e-26, 8.515779e-26, 3.571135e-26, 
    -9.065179e-26, -6.867559e-26, -2.747022e-26, 8.241077e-26, -9.065179e-26, 
    -7.142262e-26, -9.614584e-26, -4.807291e-26, -7.691667e-26, 
    -1.867977e-25, 6.043457e-26, -2.747022e-26, -4.120535e-26, 6.592862e-26, 
    6.592862e-26, -2.747022e-26, 1.648217e-26, -7.966369e-26, -1.09881e-25, 
    -9.889287e-26, -8.241071e-26, -9.339881e-26, -9.339881e-26, 6.592862e-26, 
    5.494076e-27, -1.18122e-25, 1.153751e-25, -1.922915e-26, -1.71689e-25, 
    3.983189e-26, -7.966369e-26, 2.747028e-26, 4.120564e-27, -9.889287e-26, 
    -4.120535e-26, 1.085075e-25, -1.579539e-25, -4.807291e-26, -6.867559e-26, 
    -3.845832e-26, 3.02173e-26, 1.373515e-26, 2.747052e-27, 3.02173e-26, 
    4.669945e-26, -1.016399e-25, -5.494047e-26, 6.730214e-26, -1.030134e-25, 
    -2.47232e-26, -4.120535e-26, 1.387248e-25, 5.494052e-26, -1.400982e-25, 
    -6.318154e-26, -5.219344e-26, 3.708486e-26, -1.648212e-26, -6.318154e-26, 
    -5.494047e-26, -4.669939e-26, -3.159076e-26, 3.296432e-26, -5.768749e-26, 
    -1.373486e-27, 2.472325e-26, -6.043452e-26, 2.747028e-26, -7.554316e-26, 
    -6.180803e-26, -1.442188e-25, -1.263631e-25, -2.884373e-26, 9.065185e-26, 
    -5.631398e-26, -5.768749e-26, -1.373486e-27, 1.400983e-25, -5.356696e-26, 
    -8.241071e-26, -6.318154e-26, 1.648217e-26, -4.532588e-26, -2.746998e-27, 
    6.592862e-26, -4.395237e-26, 1.318572e-25, 2.197622e-26, -1.016399e-25, 
    7.966375e-26, -5.494023e-27, 8.241101e-27, 2.675715e-32, -1.12628e-25, 
    -5.494023e-27, 9.75194e-26, -1.593274e-25, -1.922915e-26, -5.768749e-26, 
    6.31816e-26, -1.098807e-26, -4.807291e-26, -7.416964e-26, -5.631398e-26, 
    -1.15375e-25, -9.065179e-26, -1.071339e-25, -3.983183e-26, -8.927828e-26, 
    -1.37351e-26, -1.510861e-26, -4.257886e-26, -3.708481e-26, -2.334968e-26, 
    1.181221e-25, -1.922915e-26, 5.494076e-27, 9.339887e-26, 1.373539e-27, 
    1.922918e-25, -3.296427e-26, -5.494047e-26, 6.31816e-26, 9.339887e-26, 
    -2.060266e-26, -7.691667e-26, 2.675725e-32, -4.120511e-27, -4.257886e-26, 
    8.103726e-26, -7.00491e-26, 5.081998e-26, -1.043869e-25, -7.00491e-26, 
    -1.222426e-25, -2.417381e-25, -6.867535e-27, 5.21935e-26, -4.395237e-26, 
    -8.378423e-26, -1.785563e-26, -1.922915e-26, -6.592857e-26, 
    -1.236161e-25, 2.197622e-26, -1.648212e-26, 9.065185e-26, -1.09881e-25, 
    -1.37351e-26, 9.065185e-26, -7.554316e-26, 3.708486e-26, 3.159081e-26, 
    -2.403646e-25, -1.016399e-25, -8.515774e-26, 5.906106e-26, 4.669945e-26, 
    2.675723e-32, -2.197617e-26, -3.845832e-26, 8.241101e-27, -8.241047e-27, 
    -9.477233e-26, -1.785563e-26, 4.669945e-26, -1.085074e-25, 6.455511e-26, 
    1.400983e-25, 7.142267e-26, 4.120564e-27, -6.043452e-26, -3.845832e-26, 
    1.304837e-25, 3.159081e-26, 8.241077e-26, 4.807296e-26, -1.15375e-25, 
    -1.826771e-25, -2.47232e-26, 4.944647e-26, 1.648215e-25, 3.159081e-26, 
    1.263632e-25, -1.002664e-25, -3.983183e-26, 7.142267e-26, 2.609676e-26, 
    1.373539e-27, 3.159081e-26, -2.47232e-26, 8.378428e-26, -2.334968e-26, 
    -1.098807e-26, -3.845832e-26, 7.416969e-26, 1.92292e-26, -4.257886e-26, 
    -1.208691e-25, -1.249896e-25, -2.884373e-26, -4.944642e-26, 7.966375e-26, 
    3.845837e-26, -5.081993e-26, 5.494076e-27, 1.194956e-25, -3.57113e-26, 
    -5.494023e-27, -1.400982e-25, 7.416969e-26, 2.197622e-26, -9.339881e-26, 
    -6.318154e-26, -1.922915e-26, -5.219344e-26, -3.159076e-26, 8.241101e-27, 
    8.378428e-26, -3.021725e-26, 4.944647e-26, -2.22509e-25, 4.944647e-26, 
    6.043457e-26, -4.120535e-26 ;

 M_SOIL1C_TO_LEACHING =
  -1.091314e-20, 3.762666e-20, 2.10428e-20, 2.316639e-20, 3.542361e-20, 
    -4.137738e-20, 3.056405e-20, -2.766222e-21, 2.910175e-21, 1.518209e-20, 
    7.475401e-21, -6.28258e-21, 2.110275e-20, 2.936327e-20, 1.290553e-20, 
    5.475366e-21, -1.978268e-20, 1.021422e-20, -2.460266e-20, 7.551744e-21, 
    8.68211e-21, -2.834716e-20, 2.103265e-21, 1.722792e-20, 3.108907e-20, 
    3.395398e-20, -8.317664e-21, -4.200475e-20, 1.814595e-20, 3.564274e-20, 
    1.371537e-21, 1.449534e-20, -4.297233e-21, -2.834376e-20, -3.067059e-21, 
    1.065217e-20, -1.9602e-20, -5.778744e-21, -5.745375e-21, -3.172805e-20, 
    -2.589969e-22, -7.877157e-21, 7.888111e-22, -2.565101e-20, 5.724174e-21, 
    -3.998096e-20, 8.337643e-22, -3.147078e-21, -1.747079e-20, -9.53224e-21, 
    7.38436e-21, 4.482725e-20, 2.949843e-20, 1.548179e-20, 2.663888e-20, 
    1.166322e-20, -2.610596e-20, -2.847665e-20, -5.117989e-21, 3.909659e-20, 
    3.028045e-20, -4.087703e-21, -1.982113e-20, -1.80546e-20, 3.314339e-20, 
    1.751234e-20, -2.366144e-20, 1.085404e-20, -1.415917e-20, 3.303139e-21, 
    -2.124666e-20, 1.923617e-20, 4.255579e-20, 2.77226e-20, -9.350774e-21, 
    8.830839e-21, -1.772624e-22, 3.580732e-20, -1.953527e-20, 3.960634e-20, 
    1.86851e-20, 4.089671e-21, 3.733724e-21, -2.766437e-20, 2.690862e-20, 
    1.957939e-20, 1.079239e-20, 1.107598e-20, 1.020601e-20, -5.973266e-21, 
    1.298187e-20, 2.845656e-20, 2.858041e-20, -3.752799e-20, -3.95707e-20, 
    2.934181e-20, -5.286047e-20, -2.245024e-20, -2.96203e-20, 3.579663e-21, 
    -1.597995e-20, -4.443961e-21, -2.52408e-20, -1.512387e-20, -1.00703e-20, 
    -1.590356e-21, -9.1028e-21, 7.585112e-21, 2.10623e-20, 1.925709e-20, 
    -1.393693e-20, -6.269851e-21, 9.066608e-21, -4.684009e-21, 7.432709e-21, 
    -5.150309e-20, 1.638171e-20, -8.29335e-21, -2.371829e-20, 9.575504e-21, 
    1.228013e-20, 1.634426e-22, -1.140822e-21, 1.420863e-20, -2.567469e-21, 
    -3.285644e-21, -4.808966e-20, 2.956459e-20, -6.435807e-21, -2.355373e-20, 
    -4.318204e-20, 1.622905e-20, -5.350737e-20, -2.4163e-20, 5.083077e-20, 
    1.774306e-20, 8.680054e-22, -5.69713e-22, -2.700531e-20, -1.377805e-20, 
    1.848749e-20, -1.529716e-20, 3.109389e-20, 2.906491e-22, -3.070456e-21, 
    -4.278083e-20, -3.501594e-20, -1.258011e-20, -3.932745e-22, 3.197826e-20, 
    1.55075e-20, -1.258123e-20, 3.921815e-20, 1.168328e-20, 9.737489e-22, 
    4.091538e-20, 1.62833e-20, 2.363487e-20, -8.979535e-21, -2.857334e-20, 
    -1.232763e-20, 1.030638e-20, -9.545541e-21, 1.808006e-20, -2.936076e-20, 
    -7.419434e-21, 1.869049e-20, 6.856204e-21, 6.235349e-21, -3.485079e-20, 
    -2.785662e-20, 1.581879e-20, 4.106778e-20, -2.145023e-20, -1.838592e-21, 
    1.416846e-20, 1.284899e-20, -2.688261e-20, 1.655966e-21, -2.839169e-21, 
    3.499699e-20, -1.071407e-20, 3.209304e-20, -2.446441e-20, 6.798269e-21, 
    2.412484e-20, 5.495354e-20, 2.385117e-20, 8.562536e-21, 4.077825e-21, 
    3.498906e-20, 1.125747e-20, -4.715115e-21, 3.346175e-20, 3.0663e-20, 
    -1.506757e-20, -9.015156e-21, 8.628952e-21, -2.47409e-20, -3.298036e-21, 
    -8.171775e-21, 1.419139e-20, 1.229429e-20, 8.601242e-21, -2.434326e-21, 
    -1.039593e-21, 3.230595e-20, 3.566566e-20, -1.369716e-20, -1.548716e-20, 
    2.821343e-20, -1.326573e-20, -1.3512e-20, 1.678769e-20, -5.449078e-21, 
    4.756861e-20, 1.419676e-20, -1.328814e-22, 2.44398e-20, 1.983637e-20, 
    2.030656e-20, -2.782722e-20, -4.571558e-20, -2.661118e-20, 2.11152e-20, 
    4.229372e-21, -2.953984e-21, 9.710119e-21, -1.402515e-20, 4.23702e-21, 
    -1.599748e-20, 3.607392e-20, 1.070476e-20, 2.870565e-20, -1.590926e-20, 
    1.218993e-20, 1.701532e-20, 1.833509e-20, 7.242718e-21, -2.53895e-20, 
    1.651459e-20, -2.100124e-20, 2.803587e-20, 2.969226e-21, 1.063907e-21, 
    -2.238408e-20, -1.858135e-20, -3.399544e-21, 8.854842e-21, -1.788641e-20, 
    1.253346e-20, 2.665475e-20, 4.43319e-20, 5.442569e-21, 9.288561e-21, 
    -4.425583e-21, 1.389621e-20, -1.51979e-20, -2.012703e-20, 1.373278e-20, 
    -4.267199e-20, -9.539605e-21, -1.346309e-20, 2.937348e-20, 1.230248e-20, 
    -2.035719e-20, 6.432984e-21, -7.709538e-21, 2.397545e-21, -2.598635e-20, 
    -1.389708e-20, 1.611226e-20, -2.665019e-20, 4.13211e-20, 6.153069e-21, 
    -1.665453e-20, -1.354845e-20, 2.219012e-20, 1.05665e-20, -9.096863e-21, 
    6.077553e-20, 4.317468e-20, 1.122216e-20, -9.066018e-21, 2.633079e-21, 
    9.507953e-21, -3.783137e-20, -2.810572e-20, 1.742811e-20, -2.229304e-20, 
    -2.069165e-20, -4.874561e-20, 7.19663e-21, 1.203104e-20, -3.599159e-22, 
    -1.560279e-20, -3.960209e-20, 8.76087e-24, -7.741452e-21, 1.830314e-20, 
    4.232196e-21, -2.564645e-21, 3.268282e-20, -2.548676e-20, -5.567197e-20, 
    3.577762e-20, -6.373595e-21, 2.866042e-20, 2.152147e-20, -3.233112e-20, 
    -3.332538e-21, 1.312466e-20, 1.964612e-20, -1.491687e-20, -3.671598e-20, 
    4.075282e-20, 1.188489e-20, 8.762406e-21, 2.418478e-20, -7.787261e-21, 
    1.461212e-20, -7.984323e-21, 2.138859e-20, 5.16405e-20, 1.39129e-20, 
    -6.857059e-21, 1.319221e-20, -4.589455e-20, 1.45287e-20, -1.067e-20, 
    -1.675407e-20, 1.013194e-20, -2.096162e-21, 2.988126e-20, -6.293593e-21, 
    4.589173e-20, -1.450407e-20, 1.033381e-20 ;

 M_SOIL2C_TO_LEACHING =
  5.272361e-21, -1.951407e-21, 5.726998e-21, -1.245854e-20, 8.591364e-21, 
    1.11677e-21, -5.354069e-21, -2.555408e-20, -3.46874e-20, 1.315997e-20, 
    1.007258e-20, 1.028461e-20, -1.152407e-21, -3.494126e-20, 2.505221e-20, 
    -3.993292e-21, -1.183765e-20, 7.574431e-22, 3.169185e-20, 3.611887e-20, 
    -5.874211e-20, -1.528583e-20, 5.459362e-20, 3.01719e-20, -1.107427e-20, 
    -2.233063e-20, -6.31366e-21, 1.839248e-20, -2.183755e-20, -2.579605e-20, 
    -8.006894e-22, -1.163268e-20, -3.118324e-20, 3.900613e-20, -1.613404e-20, 
    -3.787603e-20, -1.368713e-21, -1.987794e-20, 2.696658e-20, 1.440512e-20, 
    -2.614806e-20, 2.50245e-20, 4.404382e-21, 1.57812e-20, -1.401242e-20, 
    -3.793422e-21, -1.670178e-20, 4.456431e-20, -9.23971e-22, -3.07775e-20, 
    9.067115e-22, 3.655646e-22, 1.866646e-20, -4.277694e-21, 1.477523e-20, 
    -2.535839e-20, -8.006097e-21, -9.663752e-21, 1.229895e-21, -1.713236e-20, 
    -2.495098e-20, -3.056131e-22, -1.743576e-20, 7.736087e-21, 1.578882e-20, 
    -2.783203e-21, -2.558987e-21, 7.574352e-21, -3.993487e-20, 1.759065e-20, 
    2.685744e-20, 1.668283e-20, -1.313567e-20, -9.305805e-21, 6.978634e-21, 
    -9.230596e-21, 2.776416e-20, 2.179035e-20, 1.585159e-20, 2.01868e-21, 
    -8.941947e-21, 3.153308e-21, -1.995655e-20, -3.713967e-21, 1.513233e-20, 
    -3.378408e-20, -1.340258e-20, -1.772242e-20, 3.551268e-20, 2.183812e-21, 
    -3.98888e-20, 1.726042e-20, -1.505654e-20, 1.04093e-20, 1.750358e-20, 
    4.648801e-20, -1.387352e-21, -1.182778e-20, 2.680399e-20, 1.399855e-20, 
    -1.320548e-20, -1.882226e-20, 6.794874e-21, 1.916434e-20, 2.59708e-20, 
    3.899083e-20, 1.70563e-20, 2.356646e-20, -3.872084e-20, -5.496194e-22, 
    3.18861e-20, 2.885889e-20, -7.973284e-21, -7.09371e-21, -2.114346e-20, 
    1.404917e-20, 1.438421e-20, 2.5614e-20, -1.623742e-21, 3.907901e-21, 
    -1.35414e-20, 1.857599e-20, -2.842565e-21, -2.023872e-20, -3.069182e-20, 
    -2.394221e-20, 3.493196e-20, 6.236493e-21, 1.738511e-20, -1.227163e-20, 
    -1.226881e-20, 5.162155e-20, -1.836705e-20, -4.671851e-21, -3.749943e-20, 
    -8.114381e-21, 2.381724e-20, -1.240397e-20, -5.292428e-21, -1.449306e-20, 
    1.583548e-20, -1.873345e-20, -3.225929e-20, -2.022485e-20, -9.750824e-21, 
    1.300505e-20, 1.59005e-20, 7.280617e-21, 2.632706e-20, 9.208686e-22, 
    -1.806539e-20, 3.164859e-20, -2.957641e-21, -2.549609e-20, 8.542425e-21, 
    -1.608455e-20, 7.274942e-21, 2.526681e-20, -1.007655e-20, -2.275703e-21, 
    2.610904e-20, -1.752281e-20, -2.627404e-21, -5.15879e-20, -8.514993e-21, 
    2.708985e-20, 4.846573e-20, -4.254542e-21, -1.279075e-20, -2.963385e-20, 
    2.004393e-20, 3.257456e-20, 6.419682e-21, 5.012246e-21, -2.399168e-20, 
    6.943587e-21, -2.091753e-23, 2.360491e-20, -9.983508e-21, 7.478264e-22, 
    1.091086e-20, 2.200788e-21, 3.556461e-21, -2.192579e-20, 3.091551e-20, 
    -3.426415e-20, -3.747587e-21, -3.560033e-20, 1.120755e-21, -3.226976e-20, 
    2.186752e-20, -7.61225e-21, 1.635371e-20, 3.940023e-20, -4.089107e-20, 
    2.097071e-20, 3.348127e-20, 7.913568e-22, 1.188289e-20, -1.382808e-20, 
    4.774333e-20, -1.585781e-20, 2.521846e-20, -2.573144e-21, 1.764719e-20, 
    -2.356276e-21, 2.917556e-20, 7.310016e-21, -4.049976e-20, 1.533078e-20, 
    -8.878306e-21, -1.262676e-20, -1.048139e-20, 1.311729e-20, 3.102134e-21, 
    1.074435e-20, -5.726687e-21, 2.217117e-20, 1.790562e-20, 7.735684e-22, 
    -1.546424e-20, -2.568694e-20, 2.736976e-20, -1.85624e-20, -1.929061e-21, 
    4.635349e-21, -1.605915e-22, -2.233403e-20, 3.229437e-20, 4.149916e-21, 
    -1.67761e-20, -4.834133e-21, -9.182962e-22, -9.997664e-21, 4.954857e-20, 
    -2.172136e-20, 1.186763e-20, -1.323944e-20, -2.31042e-20, -5.910197e-21, 
    6.49886e-21, 2.950662e-20, -1.704021e-21, 2.236343e-20, 4.008527e-20, 
    -2.155286e-20, 1.74227e-20, -3.458137e-20, 1.62047e-20, 4.659883e-20, 
    -3.986475e-20, -5.844059e-21, 1.898821e-20, 2.829291e-21, -3.32435e-21, 
    -5.050422e-20, -1.620217e-20, -1.165813e-20, -2.429223e-21, 3.611208e-20, 
    -1.405729e-21, -7.848329e-21, -1.339182e-20, -3.162713e-20, -3.92939e-21, 
    -6.589328e-21, -4.010988e-20, -1.510489e-20, 2.144116e-20, 1.861586e-20, 
    3.331672e-20, 3.999513e-21, -4.324093e-21, 2.408783e-20, -3.038959e-20, 
    -2.410476e-20, 2.145445e-20, -2.323877e-20, -3.474181e-21, 2.518963e-20, 
    1.683104e-21, -4.497143e-20, -3.252054e-20, -3.359378e-20, 3.891788e-20, 
    -2.360858e-20, -3.548694e-20, -8.427375e-21, 6.066275e-21, 1.525909e-21, 
    3.398904e-20, 2.557638e-20, 2.137671e-20, 3.534249e-20, -2.803388e-20, 
    -6.117994e-21, 7.336037e-21, -3.808355e-20, 5.18667e-20, -1.476929e-20, 
    3.317958e-20, -4.709362e-20, -1.378453e-20, 6.909083e-21, -5.853937e-21, 
    4.12135e-21, 1.149216e-20, -1.078082e-20, -1.975704e-21, -6.104719e-21, 
    1.010765e-21, -2.367928e-20, 1.326742e-20, 5.519696e-20, -1.322501e-20, 
    -3.406226e-20, -1.527256e-20, 1.149583e-21, 4.045862e-21, -2.76847e-20, 
    -1.662118e-20, -4.974223e-20, -1.568533e-20, -7.235925e-21, 2.368433e-21, 
    6.991085e-21, 7.138092e-21, -1.253769e-20, 5.595245e-22, -3.068177e-21, 
    3.447618e-20, 2.392975e-20, 6.293577e-21, -3.03667e-20, -1.854288e-20, 
    -8.015403e-21, -3.321266e-20, -7.452803e-21 ;

 M_SOIL3C_TO_LEACHING =
  1.057696e-20, 5.467455e-21, 1.364263e-20, 6.535876e-21, 1.456261e-20, 
    -5.792617e-20, -1.260417e-20, 1.990877e-20, -4.24424e-20, 3.577689e-21, 
    1.334348e-20, -3.335363e-21, 1.769837e-20, -2.199081e-20, 1.386258e-20, 
    4.836958e-21, -1.717562e-20, 1.130159e-20, -5.923373e-22, 1.916574e-20, 
    -9.807363e-21, 4.392223e-20, 1.375401e-20, 2.423708e-20, 2.672668e-21, 
    1.184812e-20, -4.849393e-21, 2.174907e-20, 1.613518e-20, -3.145663e-20, 
    -5.215393e-20, 1.223772e-20, 1.373139e-20, -4.901138e-21, 1.696158e-20, 
    -2.003826e-20, -9.835929e-21, 4.607806e-20, -3.122988e-20, 2.483508e-20, 
    -8.535695e-22, 3.679063e-20, 1.049808e-20, 1.577272e-20, 2.349448e-22, 
    -1.243166e-20, -1.208504e-20, -5.719689e-25, 6.538155e-21, 2.498717e-20, 
    -4.921205e-21, -2.690237e-20, 5.774775e-21, -8.773114e-22, 2.165713e-21, 
    -1.243705e-20, 2.050337e-20, 3.613328e-20, -7.779323e-21, 9.981802e-21, 
    -1.991896e-20, -3.082924e-20, -2.424982e-20, -1.566781e-20, 
    -1.650326e-20, 3.798768e-20, -2.183983e-20, 2.774096e-20, -6.409493e-21, 
    -4.930277e-21, -7.091171e-21, -2.490292e-21, -2.135297e-20, 
    -2.864429e-20, 7.682652e-21, -6.061381e-20, 1.674079e-20, 1.156171e-20, 
    -2.705705e-20, 1.613178e-20, 1.220069e-20, 9.977009e-21, 1.410854e-20, 
    1.301664e-20, 2.667085e-20, 5.503128e-20, -3.109018e-20, -1.374809e-20, 
    2.157524e-21, 7.793482e-21, 1.800288e-20, 2.729822e-20, 2.955837e-20, 
    -2.216892e-20, 7.233329e-20, -3.062567e-20, 3.795937e-21, 8.372207e-21, 
    5.256236e-21, 1.291911e-20, 1.215462e-20, -1.12688e-20, -2.021612e-20, 
    -2.02783e-20, 1.907009e-21, 1.832153e-20, 8.038321e-21, -4.211953e-20, 
    2.571295e-20, -8.381833e-21, 2.598635e-20, -2.400674e-21, 7.127079e-21, 
    1.465111e-20, -6.649835e-21, -3.449852e-20, -2.183304e-20, 3.005966e-20, 
    3.870045e-21, -6.570951e-21, -4.806763e-20, -1.291572e-20, -3.978595e-21, 
    -2.93746e-20, 1.309186e-20, 3.082953e-20, 3.055272e-20, -5.766586e-21, 
    -3.037405e-20, 2.223028e-20, -2.061333e-20, -7.764636e-21, -6.78217e-21, 
    9.652992e-21, -1.548489e-20, 1.628867e-20, -1.897179e-20, -2.220282e-21, 
    -3.684577e-20, 1.071859e-20, 1.275228e-20, -4.003861e-20, 5.55456e-21, 
    -2.270338e-21, 4.277149e-20, 3.601153e-21, 3.896089e-20, -2.488397e-20, 
    -9.843865e-21, -2.11101e-20, 3.959417e-20, -5.100747e-21, -4.855874e-20, 
    -1.219503e-20, 1.606109e-20, 1.284985e-20, -1.63031e-20, 1.011665e-20, 
    -2.691045e-21, 1.118199e-20, -6.59581e-21, -1.21105e-20, -2.441184e-20, 
    -3.989049e-20, 2.903956e-20, -2.025399e-20, -2.350256e-20, 3.286181e-20, 
    1.766104e-20, 9.641056e-22, -2.209145e-20, -3.909574e-20, 4.829047e-21, 
    -4.144352e-20, -3.756843e-20, -4.222863e-21, -2.535021e-20, 
    -1.328919e-20, -4.149216e-20, 3.077299e-20, -1.997778e-20, -2.207269e-21, 
    -2.2567e-20, 2.644184e-20, -7.85709e-21, -9.176008e-21, -2.722527e-20, 
    -1.657362e-21, -1.724826e-20, 3.443747e-20, -2.082315e-21, 2.27652e-20, 
    4.66206e-20, 1.199117e-20, 8.09939e-21, -7.330908e-21, -2.993751e-20, 
    1.336043e-20, 6.859528e-20, 1.775834e-21, -1.229595e-20, -1.903768e-20, 
    1.156637e-21, -2.364929e-20, -2.16501e-20, 1.052691e-20, -2.261762e-20, 
    -1.119132e-20, -6.013133e-21, -1.349759e-20, 3.948534e-20, -5.358737e-20, 
    3.334782e-20, 2.157601e-20, 3.084642e-22, 2.187685e-20, 1.51849e-20, 
    8.254879e-21, 4.350009e-20, 8.280059e-21, 3.771008e-20, -1.982513e-21, 
    9.064094e-21, 4.045453e-20, 2.186497e-20, 2.619787e-21, -7.78895e-21, 
    1.176896e-20, 1.768452e-20, 2.270779e-20, -3.626927e-20, 1.125778e-20, 
    2.324359e-20, 2.186754e-20, -2.188675e-20, -1.659518e-20, 4.110621e-21, 
    1.314643e-20, -3.50954e-21, -5.167473e-21, 1.557566e-20, 1.115318e-20, 
    -1.120264e-20, -1.936364e-20, -1.732741e-20, 1.155719e-20, -4.130705e-21, 
    1.292023e-20, -4.574215e-20, -2.84676e-20, -2.797705e-20, -2.944726e-20, 
    -3.315273e-20, 4.396321e-20, 2.782043e-20, -2.496003e-20, 1.376898e-20, 
    4.781253e-21, -2.747324e-20, -1.022182e-20, -1.037904e-20, 2.570391e-20, 
    -2.875289e-20, 1.451426e-20, -9.837897e-21, 1.227843e-20, 1.428243e-20, 
    -3.743609e-20, -1.275086e-20, 5.54997e-21, -4.460086e-21, -1.144219e-21, 
    -4.895774e-21, 2.44476e-21, -2.094271e-20, 4.80022e-21, -3.320382e-21, 
    -1.843334e-22, -2.113245e-20, 5.412035e-21, 2.624957e-20, 3.197134e-21, 
    1.864074e-20, 1.927665e-21, -4.502778e-21, -2.420712e-20, -2.546302e-20, 
    -1.857202e-20, 5.340795e-21, 7.081554e-21, -8.961703e-21, -1.627482e-20, 
    -5.777054e-21, -3.458938e-21, -9.595914e-22, 1.884486e-20, -2.121903e-21, 
    -1.548998e-20, -2.992507e-20, -3.597665e-20, -2.08839e-20, 2.750547e-20, 
    -2.869886e-20, -1.074498e-22, 2.265635e-20, -1.73034e-20, -1.73806e-20, 
    -6.37722e-20, 1.582387e-20, 2.517862e-20, -1.394768e-20, 9.392599e-21, 
    -3.795997e-20, -2.324444e-20, -1.853809e-20, 3.432183e-20, -3.145972e-20, 
    -2.743307e-20, -4.589572e-21, -4.580465e-20, 2.295209e-20, 2.479296e-20, 
    5.302323e-21, 2.894427e-20, 2.283589e-20, -1.290091e-21, 1.646114e-20, 
    -3.865751e-20, -2.627021e-20, -1.974761e-20, 2.255455e-20, 4.705912e-20, 
    7.807607e-21, 2.513618e-20, -3.360876e-20, 1.962717e-20, 1.207175e-20, 
    -2.179823e-20 ;

 NBP =
  -6.195836e-08, -6.223155e-08, -6.217844e-08, -6.23988e-08, -6.227657e-08, 
    -6.242085e-08, -6.201375e-08, -6.224239e-08, -6.209643e-08, 
    -6.198296e-08, -6.282642e-08, -6.240863e-08, -6.326049e-08, -6.2994e-08, 
    -6.366348e-08, -6.321901e-08, -6.375311e-08, -6.365067e-08, 
    -6.395901e-08, -6.387068e-08, -6.426506e-08, -6.399979e-08, 
    -6.446953e-08, -6.420172e-08, -6.424361e-08, -6.399104e-08, 
    -6.249272e-08, -6.27744e-08, -6.247603e-08, -6.251619e-08, -6.249817e-08, 
    -6.227909e-08, -6.216867e-08, -6.193749e-08, -6.197946e-08, 
    -6.214927e-08, -6.253426e-08, -6.240357e-08, -6.273295e-08, 
    -6.272551e-08, -6.309222e-08, -6.292688e-08, -6.354328e-08, 
    -6.336808e-08, -6.387437e-08, -6.374704e-08, -6.386838e-08, 
    -6.383159e-08, -6.386886e-08, -6.368212e-08, -6.376213e-08, 
    -6.359781e-08, -6.295784e-08, -6.314591e-08, -6.2585e-08, -6.224774e-08, 
    -6.202378e-08, -6.186485e-08, -6.188731e-08, -6.193014e-08, 
    -6.215026e-08, -6.235724e-08, -6.251497e-08, -6.262048e-08, 
    -6.272445e-08, -6.303911e-08, -6.32057e-08, -6.357869e-08, -6.351139e-08, 
    -6.362541e-08, -6.373437e-08, -6.391728e-08, -6.388717e-08, 
    -6.396776e-08, -6.362242e-08, -6.385192e-08, -6.347305e-08, 
    -6.357667e-08, -6.275266e-08, -6.243883e-08, -6.23054e-08, -6.218865e-08, 
    -6.190459e-08, -6.210075e-08, -6.202342e-08, -6.220741e-08, 
    -6.232432e-08, -6.22665e-08, -6.262336e-08, -6.248462e-08, -6.321557e-08, 
    -6.290072e-08, -6.372166e-08, -6.352521e-08, -6.376875e-08, 
    -6.364448e-08, -6.385741e-08, -6.366577e-08, -6.399775e-08, 
    -6.407004e-08, -6.402064e-08, -6.421042e-08, -6.365515e-08, 
    -6.386838e-08, -6.226487e-08, -6.22743e-08, -6.231824e-08, -6.212511e-08, 
    -6.21133e-08, -6.193633e-08, -6.20938e-08, -6.216086e-08, -6.23311e-08, 
    -6.243179e-08, -6.252751e-08, -6.273797e-08, -6.297304e-08, 
    -6.330175e-08, -6.353794e-08, -6.369626e-08, -6.359918e-08, 
    -6.368489e-08, -6.358908e-08, -6.354417e-08, -6.404295e-08, 
    -6.376287e-08, -6.418312e-08, -6.415987e-08, -6.396967e-08, 
    -6.416249e-08, -6.228093e-08, -6.222666e-08, -6.203825e-08, -6.21857e-08, 
    -6.191706e-08, -6.206743e-08, -6.215388e-08, -6.248751e-08, 
    -6.256082e-08, -6.262879e-08, -6.276304e-08, -6.293534e-08, 
    -6.323759e-08, -6.35006e-08, -6.374071e-08, -6.372311e-08, -6.372931e-08, 
    -6.378295e-08, -6.365008e-08, -6.380476e-08, -6.383071e-08, 
    -6.376284e-08, -6.415675e-08, -6.404422e-08, -6.415937e-08, -6.40861e-08, 
    -6.22443e-08, -6.233561e-08, -6.228627e-08, -6.237905e-08, -6.231368e-08, 
    -6.260434e-08, -6.269149e-08, -6.309931e-08, -6.293195e-08, 
    -6.319831e-08, -6.2959e-08, -6.300141e-08, -6.320698e-08, -6.297194e-08, 
    -6.348608e-08, -6.313749e-08, -6.378503e-08, -6.343689e-08, 
    -6.380684e-08, -6.373967e-08, -6.38509e-08, -6.395051e-08, -6.407584e-08, 
    -6.430709e-08, -6.425354e-08, -6.444694e-08, -6.247174e-08, 
    -6.259017e-08, -6.257976e-08, -6.270371e-08, -6.279537e-08, 
    -6.299408e-08, -6.331277e-08, -6.319293e-08, -6.341295e-08, 
    -6.345712e-08, -6.312285e-08, -6.332808e-08, -6.266944e-08, 
    -6.277585e-08, -6.27125e-08, -6.248108e-08, -6.322053e-08, -6.284102e-08, 
    -6.354184e-08, -6.333624e-08, -6.393631e-08, -6.363786e-08, 
    -6.422406e-08, -6.447465e-08, -6.471054e-08, -6.498618e-08, 
    -6.265482e-08, -6.257435e-08, -6.271845e-08, -6.291781e-08, 
    -6.310282e-08, -6.334877e-08, -6.337395e-08, -6.342002e-08, 
    -6.353938e-08, -6.363974e-08, -6.343458e-08, -6.36649e-08, -6.28005e-08, 
    -6.325348e-08, -6.254392e-08, -6.275756e-08, -6.290607e-08, 
    -6.284093e-08, -6.317924e-08, -6.325897e-08, -6.358299e-08, 
    -6.341549e-08, -6.44128e-08, -6.397154e-08, -6.519609e-08, -6.485385e-08, 
    -6.254623e-08, -6.265455e-08, -6.303155e-08, -6.285217e-08, -6.33652e-08, 
    -6.349148e-08, -6.359415e-08, -6.372539e-08, -6.373956e-08, 
    -6.381732e-08, -6.36899e-08, -6.381229e-08, -6.33493e-08, -6.355619e-08, 
    -6.298847e-08, -6.312663e-08, -6.306308e-08, -6.299335e-08, 
    -6.320855e-08, -6.343781e-08, -6.344272e-08, -6.351623e-08, 
    -6.372337e-08, -6.336728e-08, -6.446972e-08, -6.378883e-08, 
    -6.277267e-08, -6.298131e-08, -6.301112e-08, -6.29303e-08, -6.347882e-08, 
    -6.328006e-08, -6.381542e-08, -6.367073e-08, -6.390781e-08, -6.379e-08, 
    -6.377267e-08, -6.362136e-08, -6.352716e-08, -6.328918e-08, 
    -6.309555e-08, -6.294202e-08, -6.297773e-08, -6.314637e-08, 
    -6.345184e-08, -6.374083e-08, -6.367753e-08, -6.388979e-08, -6.3328e-08, 
    -6.356355e-08, -6.347251e-08, -6.370992e-08, -6.318974e-08, 
    -6.363265e-08, -6.307653e-08, -6.312529e-08, -6.327612e-08, 
    -6.357952e-08, -6.364667e-08, -6.371835e-08, -6.367412e-08, 
    -6.345959e-08, -6.342446e-08, -6.327246e-08, -6.323049e-08, 
    -6.311468e-08, -6.301879e-08, -6.310639e-08, -6.319839e-08, 
    -6.345969e-08, -6.369518e-08, -6.395192e-08, -6.401477e-08, 
    -6.431474e-08, -6.407053e-08, -6.447351e-08, -6.413087e-08, 
    -6.472403e-08, -6.365835e-08, -6.412082e-08, -6.328299e-08, 
    -6.337325e-08, -6.353649e-08, -6.391095e-08, -6.37088e-08, -6.394522e-08, 
    -6.342308e-08, -6.315219e-08, -6.308211e-08, -6.295136e-08, -6.30851e-08, 
    -6.307422e-08, -6.320221e-08, -6.316108e-08, -6.346837e-08, -6.33033e-08, 
    -6.377223e-08, -6.394335e-08, -6.442666e-08, -6.472296e-08, 
    -6.502461e-08, -6.515778e-08, -6.519831e-08, -6.521526e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.195836e-08, -6.223155e-08, -6.217844e-08, -6.23988e-08, -6.227657e-08, 
    -6.242085e-08, -6.201375e-08, -6.224239e-08, -6.209643e-08, 
    -6.198296e-08, -6.282642e-08, -6.240863e-08, -6.326049e-08, -6.2994e-08, 
    -6.366348e-08, -6.321901e-08, -6.375311e-08, -6.365067e-08, 
    -6.395901e-08, -6.387068e-08, -6.426506e-08, -6.399979e-08, 
    -6.446953e-08, -6.420172e-08, -6.424361e-08, -6.399104e-08, 
    -6.249272e-08, -6.27744e-08, -6.247603e-08, -6.251619e-08, -6.249817e-08, 
    -6.227909e-08, -6.216867e-08, -6.193749e-08, -6.197946e-08, 
    -6.214927e-08, -6.253426e-08, -6.240357e-08, -6.273295e-08, 
    -6.272551e-08, -6.309222e-08, -6.292688e-08, -6.354328e-08, 
    -6.336808e-08, -6.387437e-08, -6.374704e-08, -6.386838e-08, 
    -6.383159e-08, -6.386886e-08, -6.368212e-08, -6.376213e-08, 
    -6.359781e-08, -6.295784e-08, -6.314591e-08, -6.2585e-08, -6.224774e-08, 
    -6.202378e-08, -6.186485e-08, -6.188731e-08, -6.193014e-08, 
    -6.215026e-08, -6.235724e-08, -6.251497e-08, -6.262048e-08, 
    -6.272445e-08, -6.303911e-08, -6.32057e-08, -6.357869e-08, -6.351139e-08, 
    -6.362541e-08, -6.373437e-08, -6.391728e-08, -6.388717e-08, 
    -6.396776e-08, -6.362242e-08, -6.385192e-08, -6.347305e-08, 
    -6.357667e-08, -6.275266e-08, -6.243883e-08, -6.23054e-08, -6.218865e-08, 
    -6.190459e-08, -6.210075e-08, -6.202342e-08, -6.220741e-08, 
    -6.232432e-08, -6.22665e-08, -6.262336e-08, -6.248462e-08, -6.321557e-08, 
    -6.290072e-08, -6.372166e-08, -6.352521e-08, -6.376875e-08, 
    -6.364448e-08, -6.385741e-08, -6.366577e-08, -6.399775e-08, 
    -6.407004e-08, -6.402064e-08, -6.421042e-08, -6.365515e-08, 
    -6.386838e-08, -6.226487e-08, -6.22743e-08, -6.231824e-08, -6.212511e-08, 
    -6.21133e-08, -6.193633e-08, -6.20938e-08, -6.216086e-08, -6.23311e-08, 
    -6.243179e-08, -6.252751e-08, -6.273797e-08, -6.297304e-08, 
    -6.330175e-08, -6.353794e-08, -6.369626e-08, -6.359918e-08, 
    -6.368489e-08, -6.358908e-08, -6.354417e-08, -6.404295e-08, 
    -6.376287e-08, -6.418312e-08, -6.415987e-08, -6.396967e-08, 
    -6.416249e-08, -6.228093e-08, -6.222666e-08, -6.203825e-08, -6.21857e-08, 
    -6.191706e-08, -6.206743e-08, -6.215388e-08, -6.248751e-08, 
    -6.256082e-08, -6.262879e-08, -6.276304e-08, -6.293534e-08, 
    -6.323759e-08, -6.35006e-08, -6.374071e-08, -6.372311e-08, -6.372931e-08, 
    -6.378295e-08, -6.365008e-08, -6.380476e-08, -6.383071e-08, 
    -6.376284e-08, -6.415675e-08, -6.404422e-08, -6.415937e-08, -6.40861e-08, 
    -6.22443e-08, -6.233561e-08, -6.228627e-08, -6.237905e-08, -6.231368e-08, 
    -6.260434e-08, -6.269149e-08, -6.309931e-08, -6.293195e-08, 
    -6.319831e-08, -6.2959e-08, -6.300141e-08, -6.320698e-08, -6.297194e-08, 
    -6.348608e-08, -6.313749e-08, -6.378503e-08, -6.343689e-08, 
    -6.380684e-08, -6.373967e-08, -6.38509e-08, -6.395051e-08, -6.407584e-08, 
    -6.430709e-08, -6.425354e-08, -6.444694e-08, -6.247174e-08, 
    -6.259017e-08, -6.257976e-08, -6.270371e-08, -6.279537e-08, 
    -6.299408e-08, -6.331277e-08, -6.319293e-08, -6.341295e-08, 
    -6.345712e-08, -6.312285e-08, -6.332808e-08, -6.266944e-08, 
    -6.277585e-08, -6.27125e-08, -6.248108e-08, -6.322053e-08, -6.284102e-08, 
    -6.354184e-08, -6.333624e-08, -6.393631e-08, -6.363786e-08, 
    -6.422406e-08, -6.447465e-08, -6.471054e-08, -6.498618e-08, 
    -6.265482e-08, -6.257435e-08, -6.271845e-08, -6.291781e-08, 
    -6.310282e-08, -6.334877e-08, -6.337395e-08, -6.342002e-08, 
    -6.353938e-08, -6.363974e-08, -6.343458e-08, -6.36649e-08, -6.28005e-08, 
    -6.325348e-08, -6.254392e-08, -6.275756e-08, -6.290607e-08, 
    -6.284093e-08, -6.317924e-08, -6.325897e-08, -6.358299e-08, 
    -6.341549e-08, -6.44128e-08, -6.397154e-08, -6.519609e-08, -6.485385e-08, 
    -6.254623e-08, -6.265455e-08, -6.303155e-08, -6.285217e-08, -6.33652e-08, 
    -6.349148e-08, -6.359415e-08, -6.372539e-08, -6.373956e-08, 
    -6.381732e-08, -6.36899e-08, -6.381229e-08, -6.33493e-08, -6.355619e-08, 
    -6.298847e-08, -6.312663e-08, -6.306308e-08, -6.299335e-08, 
    -6.320855e-08, -6.343781e-08, -6.344272e-08, -6.351623e-08, 
    -6.372337e-08, -6.336728e-08, -6.446972e-08, -6.378883e-08, 
    -6.277267e-08, -6.298131e-08, -6.301112e-08, -6.29303e-08, -6.347882e-08, 
    -6.328006e-08, -6.381542e-08, -6.367073e-08, -6.390781e-08, -6.379e-08, 
    -6.377267e-08, -6.362136e-08, -6.352716e-08, -6.328918e-08, 
    -6.309555e-08, -6.294202e-08, -6.297773e-08, -6.314637e-08, 
    -6.345184e-08, -6.374083e-08, -6.367753e-08, -6.388979e-08, -6.3328e-08, 
    -6.356355e-08, -6.347251e-08, -6.370992e-08, -6.318974e-08, 
    -6.363265e-08, -6.307653e-08, -6.312529e-08, -6.327612e-08, 
    -6.357952e-08, -6.364667e-08, -6.371835e-08, -6.367412e-08, 
    -6.345959e-08, -6.342446e-08, -6.327246e-08, -6.323049e-08, 
    -6.311468e-08, -6.301879e-08, -6.310639e-08, -6.319839e-08, 
    -6.345969e-08, -6.369518e-08, -6.395192e-08, -6.401477e-08, 
    -6.431474e-08, -6.407053e-08, -6.447351e-08, -6.413087e-08, 
    -6.472403e-08, -6.365835e-08, -6.412082e-08, -6.328299e-08, 
    -6.337325e-08, -6.353649e-08, -6.391095e-08, -6.37088e-08, -6.394522e-08, 
    -6.342308e-08, -6.315219e-08, -6.308211e-08, -6.295136e-08, -6.30851e-08, 
    -6.307422e-08, -6.320221e-08, -6.316108e-08, -6.346837e-08, -6.33033e-08, 
    -6.377223e-08, -6.394335e-08, -6.442666e-08, -6.472296e-08, 
    -6.502461e-08, -6.515778e-08, -6.519831e-08, -6.521526e-08 ;

 NET_NMIN =
  8.728431e-09, 8.766915e-09, 8.759435e-09, 8.790474e-09, 8.773257e-09, 
    8.793581e-09, 8.736235e-09, 8.768443e-09, 8.747882e-09, 8.731897e-09, 
    8.850712e-09, 8.79186e-09, 8.911858e-09, 8.874319e-09, 8.968625e-09, 
    8.906015e-09, 8.98125e-09, 8.966821e-09, 9.010256e-09, 8.997812e-09, 
    9.053367e-09, 9.016e-09, 9.08217e-09, 9.044444e-09, 9.050344e-09, 
    9.014766e-09, 8.803704e-09, 8.843384e-09, 8.801353e-09, 8.807011e-09, 
    8.804473e-09, 8.773611e-09, 8.758058e-09, 8.725491e-09, 8.731404e-09, 
    8.755324e-09, 8.809556e-09, 8.791147e-09, 8.837546e-09, 8.836498e-09, 
    8.888154e-09, 8.864864e-09, 8.951692e-09, 8.927014e-09, 8.998332e-09, 
    8.980395e-09, 8.997489e-09, 8.992306e-09, 8.997556e-09, 8.97125e-09, 
    8.982521e-09, 8.959375e-09, 8.869224e-09, 8.895717e-09, 8.816705e-09, 
    8.769196e-09, 8.737647e-09, 8.715258e-09, 8.718423e-09, 8.724457e-09, 
    8.755464e-09, 8.78462e-09, 8.80684e-09, 8.821702e-09, 8.836348e-09, 
    8.880673e-09, 8.90414e-09, 8.956682e-09, 8.947201e-09, 8.963263e-09, 
    8.978611e-09, 9.004377e-09, 9.000136e-09, 9.011488e-09, 8.962841e-09, 
    8.995171e-09, 8.9418e-09, 8.956397e-09, 8.840322e-09, 8.796114e-09, 
    8.777318e-09, 8.760872e-09, 8.720857e-09, 8.74849e-09, 8.737596e-09, 
    8.763514e-09, 8.779983e-09, 8.771838e-09, 8.822108e-09, 8.802564e-09, 
    8.905531e-09, 8.861178e-09, 8.976821e-09, 8.949147e-09, 8.983454e-09, 
    8.965948e-09, 8.995944e-09, 8.968948e-09, 9.015713e-09, 9.025895e-09, 
    9.018937e-09, 9.045669e-09, 8.967452e-09, 8.997488e-09, 8.771609e-09, 
    8.772938e-09, 8.779127e-09, 8.751922e-09, 8.750257e-09, 8.725329e-09, 
    8.747511e-09, 8.756957e-09, 8.780938e-09, 8.795122e-09, 8.808606e-09, 
    8.838254e-09, 8.871366e-09, 8.917671e-09, 8.95094e-09, 8.973243e-09, 
    8.959568e-09, 8.97164e-09, 8.958144e-09, 8.951819e-09, 9.022079e-09, 
    8.982626e-09, 9.041824e-09, 9.038549e-09, 9.011757e-09, 9.038918e-09, 
    8.773871e-09, 8.766227e-09, 8.739685e-09, 8.760456e-09, 8.722615e-09, 
    8.743796e-09, 8.755975e-09, 8.802971e-09, 8.813299e-09, 8.822873e-09, 
    8.841785e-09, 8.866055e-09, 8.908632e-09, 8.945681e-09, 8.979504e-09, 
    8.977026e-09, 8.977898e-09, 8.985453e-09, 8.966738e-09, 8.988526e-09, 
    8.992183e-09, 8.982622e-09, 9.03811e-09, 9.022258e-09, 9.038479e-09, 
    9.028158e-09, 8.768712e-09, 8.781574e-09, 8.774624e-09, 8.787693e-09, 
    8.778485e-09, 8.819429e-09, 8.831705e-09, 8.889153e-09, 8.865577e-09, 
    8.9031e-09, 8.869389e-09, 8.875362e-09, 8.904321e-09, 8.871211e-09, 
    8.943637e-09, 8.894531e-09, 8.985747e-09, 8.936706e-09, 8.98882e-09, 
    8.979358e-09, 8.995026e-09, 9.009058e-09, 9.026713e-09, 9.059287e-09, 
    9.051743e-09, 9.078986e-09, 8.80075e-09, 8.817433e-09, 8.815966e-09, 
    8.833426e-09, 8.846339e-09, 8.874329e-09, 8.919223e-09, 8.902341e-09, 
    8.933335e-09, 8.939557e-09, 8.89247e-09, 8.921379e-09, 8.8286e-09, 
    8.843588e-09, 8.834665e-09, 8.802066e-09, 8.90623e-09, 8.85277e-09, 
    8.95149e-09, 8.922528e-09, 9.007056e-09, 8.965017e-09, 9.047591e-09, 
    9.08289e-09, 9.116119e-09, 9.154946e-09, 8.82654e-09, 8.815204e-09, 
    8.835503e-09, 8.863586e-09, 8.889648e-09, 8.924294e-09, 8.92784e-09, 
    8.934331e-09, 8.951145e-09, 8.965281e-09, 8.936381e-09, 8.968825e-09, 
    8.847062e-09, 8.91087e-09, 8.810917e-09, 8.841012e-09, 8.861932e-09, 
    8.852756e-09, 8.900412e-09, 8.911644e-09, 8.957287e-09, 8.933693e-09, 
    9.074177e-09, 9.01202e-09, 9.184515e-09, 9.136306e-09, 8.811242e-09, 
    8.826501e-09, 8.879608e-09, 8.854339e-09, 8.926608e-09, 8.944397e-09, 
    8.958859e-09, 8.977345e-09, 8.979342e-09, 8.990296e-09, 8.972346e-09, 
    8.989587e-09, 8.924368e-09, 8.953513e-09, 8.873539e-09, 8.893003e-09, 
    8.884049e-09, 8.874227e-09, 8.904541e-09, 8.936836e-09, 8.937528e-09, 
    8.947883e-09, 8.977062e-09, 8.926901e-09, 9.082195e-09, 8.986284e-09, 
    8.84314e-09, 8.87253e-09, 8.87673e-09, 8.865346e-09, 8.942614e-09, 
    8.914616e-09, 8.990028e-09, 8.969647e-09, 9.003043e-09, 8.986447e-09, 
    8.984006e-09, 8.962692e-09, 8.949423e-09, 8.915899e-09, 8.888623e-09, 
    8.866997e-09, 8.872026e-09, 8.895783e-09, 8.938812e-09, 8.979522e-09, 
    8.970604e-09, 9.000504e-09, 8.921368e-09, 8.954549e-09, 8.941724e-09, 
    8.975166e-09, 8.901892e-09, 8.964284e-09, 8.885944e-09, 8.892813e-09, 
    8.91406e-09, 8.956799e-09, 8.966258e-09, 8.976354e-09, 8.970124e-09, 
    8.939905e-09, 8.934955e-09, 8.913544e-09, 8.907631e-09, 8.891318e-09, 
    8.87781e-09, 8.890151e-09, 8.90311e-09, 8.939918e-09, 8.97309e-09, 
    9.009257e-09, 9.018109e-09, 9.060365e-09, 9.025964e-09, 9.08273e-09, 
    9.034465e-09, 9.118018e-09, 8.967902e-09, 9.033048e-09, 8.915027e-09, 
    8.927741e-09, 8.950737e-09, 9.003484e-09, 8.97501e-09, 9.008311e-09, 
    8.934761e-09, 8.896602e-09, 8.88673e-09, 8.868311e-09, 8.887151e-09, 
    8.885619e-09, 8.903648e-09, 8.897855e-09, 8.94114e-09, 8.91789e-09, 
    8.983944e-09, 9.008049e-09, 9.076131e-09, 9.117868e-09, 9.16036e-09, 
    9.179119e-09, 9.184828e-09, 9.187215e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.044949e-14, 5.058576e-14, 5.055929e-14, 5.066909e-14, 5.060821e-14, 
    5.068008e-14, 5.047715e-14, 5.059115e-14, 5.051839e-14, 5.046179e-14, 
    5.088186e-14, 5.067399e-14, 5.109757e-14, 5.096525e-14, 5.129742e-14, 
    5.107696e-14, 5.134183e-14, 5.129111e-14, 5.144381e-14, 5.140008e-14, 
    5.159509e-14, 5.146398e-14, 5.169611e-14, 5.156382e-14, 5.158451e-14, 
    5.145965e-14, 5.071589e-14, 5.085598e-14, 5.070758e-14, 5.072757e-14, 
    5.07186e-14, 5.060945e-14, 5.055439e-14, 5.04391e-14, 5.046004e-14, 
    5.054473e-14, 5.073656e-14, 5.06715e-14, 5.083547e-14, 5.083177e-14, 
    5.101405e-14, 5.093189e-14, 5.123788e-14, 5.1151e-14, 5.140191e-14, 
    5.133885e-14, 5.139894e-14, 5.138073e-14, 5.139918e-14, 5.130669e-14, 
    5.134632e-14, 5.126492e-14, 5.094728e-14, 5.10407e-14, 5.076183e-14, 
    5.059379e-14, 5.048214e-14, 5.040283e-14, 5.041405e-14, 5.043541e-14, 
    5.054522e-14, 5.064841e-14, 5.072698e-14, 5.07795e-14, 5.083124e-14, 
    5.09876e-14, 5.107037e-14, 5.125542e-14, 5.122208e-14, 5.127858e-14, 
    5.133258e-14, 5.142314e-14, 5.140825e-14, 5.144812e-14, 5.127711e-14, 
    5.139078e-14, 5.120307e-14, 5.125444e-14, 5.084517e-14, 5.068906e-14, 
    5.062253e-14, 5.056437e-14, 5.042267e-14, 5.052053e-14, 5.048196e-14, 
    5.057374e-14, 5.063201e-14, 5.06032e-14, 5.078094e-14, 5.071186e-14, 
    5.107527e-14, 5.091887e-14, 5.132628e-14, 5.122893e-14, 5.134961e-14, 
    5.128805e-14, 5.13935e-14, 5.12986e-14, 5.146297e-14, 5.149871e-14, 
    5.147428e-14, 5.156814e-14, 5.129333e-14, 5.139893e-14, 5.060239e-14, 
    5.060708e-14, 5.062899e-14, 5.053268e-14, 5.05268e-14, 5.043851e-14, 
    5.051708e-14, 5.055051e-14, 5.06354e-14, 5.068555e-14, 5.073322e-14, 
    5.083796e-14, 5.095482e-14, 5.111807e-14, 5.123524e-14, 5.131371e-14, 
    5.126561e-14, 5.130807e-14, 5.126059e-14, 5.123834e-14, 5.148531e-14, 
    5.134668e-14, 5.155464e-14, 5.154315e-14, 5.144906e-14, 5.154445e-14, 
    5.061038e-14, 5.058334e-14, 5.048937e-14, 5.056292e-14, 5.04289e-14, 
    5.050392e-14, 5.054702e-14, 5.071328e-14, 5.074981e-14, 5.078363e-14, 
    5.085044e-14, 5.09361e-14, 5.108622e-14, 5.121671e-14, 5.133573e-14, 
    5.132702e-14, 5.133008e-14, 5.135664e-14, 5.129082e-14, 5.136744e-14, 
    5.138028e-14, 5.134668e-14, 5.154161e-14, 5.148596e-14, 5.154291e-14, 
    5.150668e-14, 5.059214e-14, 5.063764e-14, 5.061305e-14, 5.065928e-14, 
    5.06267e-14, 5.077144e-14, 5.08148e-14, 5.101754e-14, 5.093441e-14, 
    5.106672e-14, 5.094787e-14, 5.096893e-14, 5.107098e-14, 5.09543e-14, 
    5.120949e-14, 5.103649e-14, 5.135767e-14, 5.118507e-14, 5.136848e-14, 
    5.133521e-14, 5.139029e-14, 5.143959e-14, 5.15016e-14, 5.161589e-14, 
    5.158944e-14, 5.168497e-14, 5.070545e-14, 5.07644e-14, 5.075924e-14, 
    5.082092e-14, 5.086651e-14, 5.09653e-14, 5.112355e-14, 5.106407e-14, 
    5.117327e-14, 5.119517e-14, 5.102928e-14, 5.113113e-14, 5.080386e-14, 
    5.085677e-14, 5.082528e-14, 5.071009e-14, 5.107774e-14, 5.088918e-14, 
    5.123717e-14, 5.11352e-14, 5.143256e-14, 5.128474e-14, 5.157487e-14, 
    5.169861e-14, 5.181506e-14, 5.195085e-14, 5.079659e-14, 5.075655e-14, 
    5.082826e-14, 5.092736e-14, 5.101932e-14, 5.114141e-14, 5.115391e-14, 
    5.117676e-14, 5.123596e-14, 5.12857e-14, 5.118396e-14, 5.129817e-14, 
    5.086898e-14, 5.109411e-14, 5.074138e-14, 5.084767e-14, 5.092153e-14, 
    5.088916e-14, 5.105728e-14, 5.109686e-14, 5.125756e-14, 5.117453e-14, 
    5.166806e-14, 5.144996e-14, 5.205423e-14, 5.188567e-14, 5.074255e-14, 
    5.079646e-14, 5.09839e-14, 5.089475e-14, 5.114957e-14, 5.12122e-14, 
    5.126311e-14, 5.132812e-14, 5.133515e-14, 5.137365e-14, 5.131056e-14, 
    5.137117e-14, 5.114167e-14, 5.124429e-14, 5.096252e-14, 5.103114e-14, 
    5.099959e-14, 5.096494e-14, 5.107183e-14, 5.118556e-14, 5.118803e-14, 
    5.122447e-14, 5.132701e-14, 5.115061e-14, 5.16961e-14, 5.135945e-14, 
    5.085523e-14, 5.095891e-14, 5.097376e-14, 5.093361e-14, 5.120592e-14, 
    5.110732e-14, 5.137272e-14, 5.130106e-14, 5.141846e-14, 5.136013e-14, 
    5.135155e-14, 5.12766e-14, 5.122989e-14, 5.111183e-14, 5.10157e-14, 
    5.093944e-14, 5.095718e-14, 5.104094e-14, 5.119252e-14, 5.133577e-14, 
    5.13044e-14, 5.140955e-14, 5.113111e-14, 5.124792e-14, 5.120278e-14, 
    5.132047e-14, 5.106248e-14, 5.128208e-14, 5.100627e-14, 5.103049e-14, 
    5.110536e-14, 5.125581e-14, 5.128914e-14, 5.132463e-14, 5.130274e-14, 
    5.119638e-14, 5.117896e-14, 5.110355e-14, 5.10827e-14, 5.102522e-14, 
    5.097758e-14, 5.102109e-14, 5.106677e-14, 5.119644e-14, 5.131315e-14, 
    5.144028e-14, 5.147139e-14, 5.161961e-14, 5.149891e-14, 5.169796e-14, 
    5.152867e-14, 5.182161e-14, 5.129486e-14, 5.152377e-14, 5.110878e-14, 
    5.115357e-14, 5.123449e-14, 5.141997e-14, 5.131992e-14, 5.143694e-14, 
    5.117828e-14, 5.104381e-14, 5.100904e-14, 5.094406e-14, 5.101053e-14, 
    5.100512e-14, 5.106868e-14, 5.104827e-14, 5.120074e-14, 5.111886e-14, 
    5.135132e-14, 5.143602e-14, 5.167495e-14, 5.182114e-14, 5.196983e-14, 
    5.203539e-14, 5.205534e-14, 5.206367e-14 ;

 POT_F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.100726e-43, 5.605194e-45, 
    3.498145e-40, 2.53635e-43, 1.405053e-39, 2.860358e-40, 3.155876e-38, 
    8.419162e-39, 2.624818e-36, 5.766906e-38, 4.399989e-35, 1.071883e-36, 
    1.939966e-36, 5.068994e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.942727e-44, 1.401298e-45, 5.228945e-41, 3.049225e-42, 8.900133e-39, 
    1.278835e-39, 8.133579e-39, 4.660608e-39, 8.192598e-39, 4.676525e-40, 
    1.613396e-39, 1.244143e-40, 2.802597e-45, 7.286752e-44, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.121039e-44, 2.031883e-43, 9.19462e-41, 3.137227e-41, 
    1.924305e-40, 1.051815e-39, 1.695091e-38, 1.079296e-38, 3.593701e-38, 
    1.834622e-40, 6.345298e-39, 1.690947e-41, 8.899506e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.39622e-43, 1.401298e-45, 8.642228e-40, 3.915788e-41, 
    1.785855e-39, 2.594924e-40, 6.893387e-39, 3.6223e-40, 5.59756e-38, 
    1.61379e-37, 7.839023e-38, 1.212262e-36, 3.067653e-40, 8.134899e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.203895e-45, 1.017343e-42, 
    4.801269e-41, 5.826459e-40, 1.27116e-40, 4.881381e-40, 1.083344e-40, 
    5.302794e-41, 1.08715e-37, 1.632183e-39, 8.222793e-37, 5.898124e-37, 
    3.697471e-38, 6.123528e-37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.401298e-45, 3.47522e-43, 2.638505e-41, 1.15981e-39, 8.837471e-40, 
    9.726132e-40, 2.220196e-39, 2.83372e-40, 3.098589e-39, 4.600644e-39, 
    1.630998e-39, 5.640851e-37, 1.106896e-37, 5.856523e-37, 2.036912e-37, 0, 
    0, 0, 0, 0, 0, 0, 3.222986e-44, 1.401298e-45, 1.793662e-43, 2.802597e-45, 
    5.605194e-45, 2.073922e-43, 4.203895e-45, 2.089476e-41, 6.305843e-44, 
    2.292201e-39, 9.419528e-42, 3.198822e-39, 1.14138e-39, 6.244441e-39, 
    2.781966e-38, 1.755172e-37, 4.722894e-36, 2.230228e-36, 3.237457e-35, 0, 
    0, 0, 0, 0, 5.605194e-45, 1.221932e-42, 1.625506e-43, 6.366099e-42, 
    1.306851e-41, 4.904545e-44, 1.575059e-42, 0, 0, 0, 0, 2.606415e-43, 0, 
    5.110676e-41, 1.80207e-42, 2.251942e-38, 2.340813e-40, 1.471128e-36, 
    4.718157e-35, 1.069506e-33, 3.474821e-32, 0, 0, 0, 1.401298e-45, 
    3.503246e-44, 2.218255e-42, 3.358912e-42, 7.146622e-42, 4.912392e-41, 
    2.409084e-40, 9.066401e-42, 3.573101e-40, 0, 4.540207e-43, 0, 0, 
    1.401298e-45, 0, 1.289195e-43, 4.97461e-43, 9.84216e-41, 6.63655e-42, 
    2.034721e-35, 3.803153e-38, 4.371386e-31, 6.681893e-33, 0, 0, 
    9.809089e-45, 0, 2.907694e-42, 2.277671e-41, 1.173952e-40, 9.156785e-40, 
    1.139511e-39, 3.752387e-39, 5.277444e-40, 3.475073e-39, 2.237874e-42, 
    6.425234e-41, 4.203895e-45, 5.324934e-44, 1.821688e-44, 5.605194e-45, 
    2.129974e-43, 9.555454e-42, 1.034298e-41, 3.392263e-41, 8.898455e-40, 
    3.009989e-42, 4.420301e-35, 2.435304e-39, 0, 4.203895e-45, 7.006492e-45, 
    1.401298e-45, 1.856861e-41, 7.076557e-43, 3.645385e-39, 3.914247e-40, 
    1.470874e-38, 2.473112e-39, 1.896537e-39, 1.804298e-40, 4.040644e-41, 
    8.239635e-43, 3.082857e-44, 1.401298e-45, 4.203895e-45, 7.426882e-44, 
    1.200072e-41, 1.162563e-39, 4.354619e-40, 1.122507e-38, 1.572257e-42, 
    7.226917e-41, 1.677214e-41, 7.204426e-40, 1.541428e-43, 2.160732e-40, 
    2.242078e-44, 5.184804e-44, 6.628142e-43, 9.319896e-41, 2.685967e-40, 
    8.211385e-40, 4.12688e-40, 1.360801e-41, 7.683319e-42, 6.235778e-43, 
    3.082857e-43, 4.344025e-44, 8.407791e-45, 3.643376e-44, 1.793662e-43, 
    1.362482e-41, 5.731339e-40, 2.841443e-38, 7.189204e-38, 5.260623e-36, 
    1.626792e-37, 4.653514e-35, 3.901921e-37, 1.275646e-33, 3.229811e-40, 
    3.37117e-37, 7.426882e-43, 3.319676e-42, 4.69449e-41, 1.543183e-38, 
    7.080719e-40, 2.572929e-38, 7.512361e-42, 8.127531e-44, 2.382207e-44, 
    2.802597e-45, 2.522337e-44, 2.101948e-44, 1.905766e-43, 9.52883e-44, 
    1.568053e-41, 1.042566e-42, 1.884194e-39, 2.502087e-38, 2.457097e-35, 
    1.256787e-33, 5.56119e-32, 2.773154e-31, 4.486484e-31, 5.4801e-31 ;

 POT_F_NIT =
  3.837638e-11, 3.870687e-11, 3.864251e-11, 3.890991e-11, 3.876146e-11, 
    3.893671e-11, 3.844325e-11, 3.871999e-11, 3.85432e-11, 3.840604e-11, 
    3.943156e-11, 3.892183e-11, 3.996478e-11, 3.963697e-11, 4.046314e-11, 
    3.991366e-11, 4.057441e-11, 4.044724e-11, 4.083065e-11, 4.072061e-11, 
    4.121304e-11, 4.088148e-11, 4.146955e-11, 4.113373e-11, 4.118616e-11, 
    4.087053e-11, 3.902418e-11, 3.936794e-11, 3.900385e-11, 3.905276e-11, 
    3.903081e-11, 3.87645e-11, 3.863064e-11, 3.835115e-11, 3.84018e-11, 
    3.860712e-11, 3.907473e-11, 3.891567e-11, 3.93172e-11, 3.930811e-11, 
    3.97576e-11, 3.95546e-11, 4.031413e-11, 4.009748e-11, 4.072519e-11, 
    4.056684e-11, 4.071773e-11, 4.067194e-11, 4.071832e-11, 4.048622e-11, 
    4.058556e-11, 4.038165e-11, 3.959263e-11, 3.982369e-11, 3.913661e-11, 
    3.872647e-11, 3.845534e-11, 3.826354e-11, 3.829061e-11, 3.834227e-11, 
    3.860832e-11, 3.885935e-11, 3.905122e-11, 3.917984e-11, 3.930679e-11, 
    3.969234e-11, 3.989723e-11, 4.035799e-11, 4.027464e-11, 4.041589e-11, 
    4.05511e-11, 4.077861e-11, 4.074111e-11, 4.08415e-11, 4.041215e-11, 
    4.069722e-11, 4.022717e-11, 4.035544e-11, 3.934133e-11, 3.895857e-11, 
    3.879643e-11, 3.865483e-11, 3.831144e-11, 3.85484e-11, 3.845489e-11, 
    3.867754e-11, 3.881936e-11, 3.874918e-11, 3.918335e-11, 3.901425e-11, 
    3.990938e-11, 3.952251e-11, 4.053532e-11, 4.029174e-11, 4.059381e-11, 
    4.043952e-11, 4.070406e-11, 4.046593e-11, 4.087889e-11, 4.096911e-11, 
    4.090744e-11, 4.114458e-11, 4.045272e-11, 4.071768e-11, 3.874724e-11, 
    3.875868e-11, 3.8812e-11, 3.857787e-11, 3.856357e-11, 3.834973e-11, 
    3.853997e-11, 3.862113e-11, 3.882758e-11, 3.894995e-11, 3.906647e-11, 
    3.932332e-11, 3.96112e-11, 4.001561e-11, 4.030749e-11, 4.050376e-11, 
    4.038335e-11, 4.048964e-11, 4.037082e-11, 4.031519e-11, 4.093528e-11, 
    4.058647e-11, 4.111041e-11, 4.108133e-11, 4.084385e-11, 4.108459e-11, 
    3.87667e-11, 3.870088e-11, 3.847281e-11, 3.865122e-11, 3.832647e-11, 
    3.850806e-11, 3.861268e-11, 3.901776e-11, 3.910706e-11, 3.918996e-11, 
    3.935395e-11, 3.956494e-11, 3.99365e-11, 4.026126e-11, 4.055896e-11, 
    4.053709e-11, 4.054479e-11, 4.061142e-11, 4.044644e-11, 4.063853e-11, 
    4.06708e-11, 4.058642e-11, 4.107742e-11, 4.093683e-11, 4.108069e-11, 
    4.098911e-11, 3.872226e-11, 3.883307e-11, 3.877316e-11, 3.888584e-11, 
    3.880643e-11, 3.916014e-11, 3.926651e-11, 3.976628e-11, 3.956078e-11, 
    3.988811e-11, 3.959396e-11, 3.964599e-11, 3.989878e-11, 3.960982e-11, 
    4.024329e-11, 3.981321e-11, 4.061401e-11, 4.018243e-11, 4.064112e-11, 
    4.055763e-11, 4.06959e-11, 4.081996e-11, 4.09763e-11, 4.126561e-11, 
    4.119851e-11, 4.144108e-11, 3.899858e-11, 3.914286e-11, 3.913015e-11, 
    3.928143e-11, 3.93935e-11, 3.963701e-11, 4.00292e-11, 3.988147e-11, 
    4.015288e-11, 4.020748e-11, 3.979522e-11, 4.004806e-11, 3.923955e-11, 
    3.936957e-11, 3.929213e-11, 3.900987e-11, 3.991543e-11, 3.944932e-11, 
    4.031227e-11, 4.005809e-11, 4.080224e-11, 4.043125e-11, 4.11616e-11, 
    4.147589e-11, 4.177288e-11, 4.212129e-11, 3.922173e-11, 3.912355e-11, 
    3.929944e-11, 3.954346e-11, 3.97706e-11, 4.007362e-11, 4.010469e-11, 
    4.016161e-11, 4.030926e-11, 4.043362e-11, 4.017959e-11, 4.046481e-11, 
    3.939973e-11, 3.995603e-11, 3.908639e-11, 3.934719e-11, 3.952899e-11, 
    3.944919e-11, 3.986455e-11, 3.996277e-11, 4.036321e-11, 4.015595e-11, 
    4.139818e-11, 4.084614e-11, 4.238762e-11, 4.195382e-11, 3.908927e-11, 
    3.922138e-11, 3.968301e-11, 3.946301e-11, 4.009388e-11, 4.024997e-11, 
    4.03771e-11, 4.05399e-11, 4.05575e-11, 4.065415e-11, 4.049583e-11, 
    4.064788e-11, 4.007421e-11, 4.033004e-11, 3.963006e-11, 3.979982e-11, 
    3.972167e-11, 3.963604e-11, 3.990063e-11, 4.018353e-11, 4.018959e-11, 
    4.028053e-11, 4.053733e-11, 4.009636e-11, 4.146967e-11, 4.061865e-11, 
    3.936571e-11, 3.962132e-11, 3.965791e-11, 3.955874e-11, 4.02343e-11, 
    3.998882e-11, 4.065179e-11, 4.047205e-11, 4.076676e-11, 4.062017e-11, 
    4.059861e-11, 4.04108e-11, 4.029408e-11, 4.000002e-11, 3.976158e-11, 
    3.957306e-11, 3.961685e-11, 3.982409e-11, 4.020086e-11, 4.055902e-11, 
    4.048042e-11, 4.074426e-11, 4.004787e-11, 4.03391e-11, 4.02264e-11, 
    4.05206e-11, 3.987753e-11, 4.042483e-11, 3.973825e-11, 3.97982e-11, 
    3.998394e-11, 4.035896e-11, 4.044219e-11, 4.053113e-11, 4.047623e-11, 
    4.021049e-11, 4.016704e-11, 3.997939e-11, 3.992765e-11, 3.97851e-11, 
    3.966726e-11, 3.97749e-11, 3.98881e-11, 4.021057e-11, 4.050232e-11, 
    4.082166e-11, 4.090002e-11, 4.127515e-11, 4.096961e-11, 4.147441e-11, 
    4.104499e-11, 4.178983e-11, 4.045668e-11, 4.103252e-11, 3.999241e-11, 
    4.010379e-11, 4.030565e-11, 4.077065e-11, 4.051928e-11, 4.081335e-11, 
    4.016533e-11, 3.983125e-11, 3.974506e-11, 3.95845e-11, 3.974873e-11, 
    3.973535e-11, 3.989281e-11, 3.984217e-11, 4.022128e-11, 4.00174e-11, 
    4.0598e-11, 4.081097e-11, 4.141557e-11, 4.178849e-11, 4.216993e-11, 
    4.23389e-11, 4.23904e-11, 4.241194e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005857514, 0.0005857557, 0.0005857549, 0.0005857582, 0.0005857564, 
    0.0005857585, 0.0005857524, 0.0005857558, 0.0005857536, 0.0005857519, 
    0.0005857646, 0.0005857584, 0.0005857715, 0.0005857674, 0.0005857777, 
    0.0005857708, 0.0005857791, 0.0005857776, 0.0005857825, 0.0005857811, 
    0.0005857871, 0.0005857831, 0.0005857904, 0.0005857862, 0.0005857868, 
    0.0005857829, 0.0005857597, 0.0005857638, 0.0005857594, 0.00058576, 
    0.0005857598, 0.0005857564, 0.0005857546, 0.0005857512, 0.0005857518, 
    0.0005857544, 0.0005857603, 0.0005857584, 0.0005857634, 0.0005857633, 
    0.0005857689, 0.0005857664, 0.0005857759, 0.0005857732, 0.0005857811, 
    0.0005857791, 0.000585781, 0.0005857804, 0.000585781, 0.0005857781, 
    0.0005857793, 0.0005857768, 0.0005857669, 0.0005857697, 0.0005857611, 
    0.0005857558, 0.0005857525, 0.0005857501, 0.0005857504, 0.000585751, 
    0.0005857544, 0.0005857576, 0.00058576, 0.0005857617, 0.0005857633, 
    0.000585768, 0.0005857706, 0.0005857764, 0.0005857755, 0.0005857772, 
    0.0005857789, 0.0005857818, 0.0005857813, 0.0005857825, 0.0005857772, 
    0.0005857807, 0.0005857749, 0.0005857765, 0.0005857634, 0.0005857589, 
    0.0005857567, 0.000585755, 0.0005857507, 0.0005857536, 0.0005857525, 
    0.0005857553, 0.0005857571, 0.0005857563, 0.0005857617, 0.0005857596, 
    0.0005857708, 0.0005857659, 0.0005857787, 0.0005857756, 0.0005857794, 
    0.0005857775, 0.0005857808, 0.0005857779, 0.000585783, 0.0005857841, 
    0.0005857834, 0.0005857864, 0.0005857777, 0.000585781, 0.0005857562, 
    0.0005857563, 0.000585757, 0.000585754, 0.0005857538, 0.0005857511, 
    0.0005857536, 0.0005857546, 0.0005857573, 0.0005857588, 0.0005857602, 
    0.0005857635, 0.000585767, 0.0005857722, 0.0005857758, 0.0005857783, 
    0.0005857768, 0.0005857782, 0.0005857766, 0.000585776, 0.0005857837, 
    0.0005857793, 0.000585786, 0.0005857855, 0.0005857826, 0.0005857856, 
    0.0005857564, 0.0005857556, 0.0005857527, 0.000585755, 0.0005857509, 
    0.0005857532, 0.0005857545, 0.0005857596, 0.0005857607, 0.0005857618, 
    0.0005857639, 0.0005857665, 0.0005857712, 0.0005857752, 0.000585779, 
    0.0005857787, 0.0005857788, 0.0005857797, 0.0005857776, 0.00058578, 
    0.0005857804, 0.0005857794, 0.0005857855, 0.0005857837, 0.0005857855, 
    0.0005857844, 0.0005857559, 0.0005857573, 0.0005857566, 0.000585758, 
    0.0005857569, 0.0005857613, 0.0005857627, 0.000585769, 0.0005857665, 
    0.0005857705, 0.0005857669, 0.0005857675, 0.0005857705, 0.0005857671, 
    0.0005857749, 0.0005857695, 0.0005857797, 0.0005857741, 0.0005857801, 
    0.000585779, 0.0005857808, 0.0005857823, 0.0005857843, 0.0005857878, 
    0.000585787, 0.00058579, 0.0005857594, 0.0005857612, 0.000585761, 
    0.000585763, 0.0005857644, 0.0005857674, 0.0005857723, 0.0005857705, 
    0.0005857739, 0.0005857746, 0.0005857694, 0.0005857726, 0.0005857624, 
    0.0005857639, 0.0005857631, 0.0005857595, 0.0005857709, 0.000585765, 
    0.0005857759, 0.0005857727, 0.0005857821, 0.0005857773, 0.0005857865, 
    0.0005857904, 0.0005857942, 0.0005857984, 0.0005857622, 0.000585761, 
    0.0005857632, 0.0005857662, 0.0005857691, 0.0005857729, 0.0005857733, 
    0.000585774, 0.0005857759, 0.0005857775, 0.0005857742, 0.0005857779, 
    0.0005857642, 0.0005857714, 0.0005857605, 0.0005857637, 0.000585766, 
    0.0005857651, 0.0005857703, 0.0005857715, 0.0005857765, 0.000585774, 
    0.0005857894, 0.0005857825, 0.0005858018, 0.0005857964, 0.0005857605, 
    0.0005857622, 0.000585768, 0.0005857652, 0.0005857732, 0.0005857751, 
    0.0005857768, 0.0005857787, 0.000585779, 0.0005857802, 0.0005857782, 
    0.0005857801, 0.0005857729, 0.0005857761, 0.0005857674, 0.0005857695, 
    0.0005857685, 0.0005857674, 0.0005857708, 0.0005857743, 0.0005857744, 
    0.0005857755, 0.0005857784, 0.0005857732, 0.0005857901, 0.0005857795, 
    0.000585764, 0.0005857671, 0.0005857677, 0.0005857665, 0.0005857749, 
    0.0005857719, 0.0005857802, 0.0005857779, 0.0005857816, 0.0005857798, 
    0.0005857795, 0.0005857772, 0.0005857757, 0.000585772, 0.000585769, 
    0.0005857666, 0.0005857672, 0.0005857698, 0.0005857745, 0.000585779, 
    0.000585778, 0.0005857814, 0.0005857726, 0.0005857762, 0.0005857748, 
    0.0005857786, 0.0005857705, 0.000585777, 0.0005857687, 0.0005857695, 
    0.0005857718, 0.0005857764, 0.0005857776, 0.0005857786, 0.000585778, 
    0.0005857746, 0.0005857741, 0.0005857717, 0.000585771, 0.0005857693, 
    0.0005857678, 0.0005857692, 0.0005857705, 0.0005857747, 0.0005857783, 
    0.0005857823, 0.0005857833, 0.0005857878, 0.000585784, 0.0005857901, 
    0.0005857847, 0.0005857942, 0.0005857776, 0.0005857848, 0.0005857719, 
    0.0005857733, 0.0005857758, 0.0005857816, 0.0005857785, 0.0005857821, 
    0.0005857741, 0.0005857698, 0.0005857688, 0.0005857667, 0.0005857688, 
    0.0005857687, 0.0005857706, 0.0005857701, 0.0005857748, 0.0005857722, 
    0.0005857795, 0.0005857821, 0.0005857897, 0.0005857943, 0.0005857992, 
    0.0005858013, 0.0005858019, 0.0005858022 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  8.869452e-06, 8.895217e-06, 8.890214e-06, 8.910991e-06, 8.899478e-06, 
    8.913074e-06, 8.874689e-06, 8.896227e-06, 8.882485e-06, 8.871792e-06, 
    8.951301e-06, 8.911921e-06, 8.992404e-06, 8.967228e-06, 9.030551e-06, 
    8.988463e-06, 9.03905e-06, 9.029372e-06, 9.058596e-06, 9.050224e-06, 
    9.087552e-06, 9.062462e-06, 9.106976e-06, 9.081577e-06, 9.085536e-06, 
    9.061628e-06, 8.919877e-06, 8.946384e-06, 8.918299e-06, 8.922079e-06, 
    8.92039e-06, 8.899702e-06, 8.889259e-06, 8.867508e-06, 8.871462e-06, 
    8.887451e-06, 8.92378e-06, 8.911466e-06, 8.942577e-06, 8.941875e-06, 
    8.976519e-06, 8.960894e-06, 9.019202e-06, 9.002628e-06, 9.050574e-06, 
    9.038505e-06, 9.050001e-06, 9.046519e-06, 9.050046e-06, 9.032348e-06, 
    9.039928e-06, 9.024371e-06, 8.963812e-06, 8.981588e-06, 8.928582e-06, 
    8.896698e-06, 8.875627e-06, 8.860659e-06, 8.862775e-06, 8.8668e-06, 
    8.887544e-06, 8.907093e-06, 8.921988e-06, 8.93195e-06, 8.941774e-06, 
    8.971433e-06, 8.98722e-06, 9.022537e-06, 9.016191e-06, 9.026966e-06, 
    9.037306e-06, 9.054631e-06, 9.051783e-06, 9.05941e-06, 9.026704e-06, 
    9.048426e-06, 9.01257e-06, 9.022369e-06, 8.944324e-06, 8.914793e-06, 
    8.902147e-06, 8.891172e-06, 8.864398e-06, 8.882877e-06, 8.875588e-06, 
    8.892959e-06, 8.903985e-06, 8.898536e-06, 8.932223e-06, 8.919117e-06, 
    8.988156e-06, 8.958403e-06, 9.0361e-06, 9.017496e-06, 9.040565e-06, 
    9.028798e-06, 9.048952e-06, 9.030813e-06, 9.06226e-06, 9.069096e-06, 
    9.064422e-06, 9.082425e-06, 9.029804e-06, 9.049989e-06, 8.898378e-06, 
    8.899266e-06, 8.903417e-06, 8.885173e-06, 8.884063e-06, 8.867394e-06, 
    8.882237e-06, 8.888551e-06, 8.904633e-06, 8.914128e-06, 8.923163e-06, 
    8.94304e-06, 8.965233e-06, 8.996326e-06, 9.0187e-06, 9.033701e-06, 
    9.02451e-06, 9.032623e-06, 9.023549e-06, 9.019303e-06, 9.066527e-06, 
    9.039992e-06, 9.079835e-06, 9.077633e-06, 9.059588e-06, 9.077881e-06, 
    8.899891e-06, 8.894778e-06, 8.876995e-06, 8.890912e-06, 8.865581e-06, 
    8.879741e-06, 8.887878e-06, 8.919365e-06, 8.926316e-06, 8.932725e-06, 
    8.945415e-06, 8.961692e-06, 8.99026e-06, 9.015153e-06, 9.037913e-06, 
    9.036246e-06, 9.036832e-06, 9.041905e-06, 9.029322e-06, 9.043973e-06, 
    9.04642e-06, 9.040003e-06, 9.077337e-06, 9.066669e-06, 9.077587e-06, 
    9.070643e-06, 8.896443e-06, 8.905053e-06, 8.900398e-06, 8.909145e-06, 
    8.902973e-06, 8.93039e-06, 8.938614e-06, 8.977159e-06, 8.961365e-06, 
    8.986539e-06, 8.963932e-06, 8.967929e-06, 8.987309e-06, 8.96516e-06, 
    9.013757e-06, 8.980756e-06, 9.042103e-06, 9.009073e-06, 9.044171e-06, 
    9.037813e-06, 9.048352e-06, 9.057779e-06, 9.069665e-06, 9.091571e-06, 
    9.086502e-06, 9.10485e-06, 8.917903e-06, 8.929067e-06, 8.928107e-06, 
    8.939809e-06, 8.948461e-06, 8.967251e-06, 8.997382e-06, 8.986056e-06, 
    9.006878e-06, 9.011051e-06, 8.979433e-06, 8.998821e-06, 8.936558e-06, 
    8.946586e-06, 8.940631e-06, 8.918771e-06, 8.988634e-06, 8.952748e-06, 
    9.019066e-06, 8.999608e-06, 9.056432e-06, 9.028136e-06, 9.083707e-06, 
    9.107428e-06, 9.129874e-06, 9.155996e-06, 8.935186e-06, 8.927596e-06, 
    8.941208e-06, 8.960007e-06, 8.977524e-06, 9.000791e-06, 9.003184e-06, 
    9.007538e-06, 9.018847e-06, 9.028347e-06, 9.008892e-06, 9.030731e-06, 
    8.948866e-06, 8.991761e-06, 8.924706e-06, 8.944853e-06, 8.958908e-06, 
    8.952765e-06, 8.984767e-06, 8.992306e-06, 9.022951e-06, 9.007119e-06, 
    9.101552e-06, 9.059738e-06, 9.175975e-06, 9.143441e-06, 8.924939e-06, 
    8.935171e-06, 8.970771e-06, 8.953831e-06, 9.002356e-06, 9.014301e-06, 
    9.024035e-06, 9.036443e-06, 9.0378e-06, 9.045157e-06, 9.033099e-06, 
    9.044689e-06, 9.00084e-06, 9.020432e-06, 8.966726e-06, 8.979777e-06, 
    8.97378e-06, 8.967188e-06, 8.987538e-06, 9.009193e-06, 9.009693e-06, 
    9.016633e-06, 9.036133e-06, 9.002553e-06, 9.106883e-06, 9.042352e-06, 
    8.946328e-06, 8.966001e-06, 8.968856e-06, 8.961226e-06, 9.013102e-06, 
    8.994291e-06, 9.044983e-06, 9.031283e-06, 9.053742e-06, 9.042576e-06, 
    9.040933e-06, 9.026607e-06, 9.017681e-06, 8.995146e-06, 8.976834e-06, 
    8.962337e-06, 8.965711e-06, 8.981637e-06, 9.010527e-06, 9.037905e-06, 
    9.031902e-06, 9.052035e-06, 8.998834e-06, 9.021113e-06, 9.012489e-06, 
    9.034989e-06, 8.985747e-06, 9.027563e-06, 8.975054e-06, 8.979661e-06, 
    8.993919e-06, 9.022599e-06, 9.029004e-06, 9.035775e-06, 9.031604e-06, 
    9.011267e-06, 9.007953e-06, 8.993581e-06, 8.989596e-06, 8.978661e-06, 
    8.969593e-06, 8.977869e-06, 8.986554e-06, 9.011292e-06, 9.033579e-06, 
    9.057908e-06, 9.063878e-06, 9.092236e-06, 9.069099e-06, 9.107235e-06, 
    9.074733e-06, 9.131053e-06, 9.030042e-06, 9.073852e-06, 8.99458e-06, 
    9.003121e-06, 9.018534e-06, 9.053991e-06, 9.034883e-06, 9.057248e-06, 
    9.007827e-06, 8.982168e-06, 8.975579e-06, 8.963211e-06, 8.975861e-06, 
    8.974834e-06, 8.98694e-06, 8.983051e-06, 9.012114e-06, 8.996501e-06, 
    9.040881e-06, 9.05708e-06, 9.102913e-06, 9.131013e-06, 9.159698e-06, 
    9.172349e-06, 9.176203e-06, 9.177813e-06 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.68618, 81.68539, 81.68554, 81.6849, 81.68525, 81.68484, 81.68601, 
    81.68536, 81.68578, 81.6861, 81.68369, 81.68487, 81.6824, 81.68316, 
    81.68121, 81.68252, 81.68095, 81.68124, 81.68033, 81.68059, 81.67946, 
    81.68021, 81.67885, 81.67963, 81.67951, 81.68024, 81.68462, 81.68384, 
    81.68467, 81.68456, 81.6846, 81.68524, 81.68558, 81.68623, 81.68611, 
    81.68562, 81.6845, 81.68488, 81.68391, 81.68393, 81.68287, 81.68335, 
    81.68155, 81.68206, 81.68057, 81.68095, 81.6806, 81.6807, 81.6806, 
    81.68114, 81.68091, 81.68139, 81.68327, 81.68272, 81.68435, 81.68536, 
    81.68599, 81.68645, 81.68638, 81.68626, 81.68562, 81.68501, 81.68455, 
    81.68424, 81.68394, 81.68305, 81.68256, 81.68146, 81.68164, 81.68132, 
    81.68098, 81.68046, 81.68054, 81.68031, 81.68131, 81.68065, 81.68175, 
    81.68145, 81.68391, 81.68478, 81.68519, 81.68551, 81.68633, 81.68577, 
    81.68599, 81.68545, 81.6851, 81.68527, 81.68423, 81.68464, 81.68253, 
    81.68343, 81.68103, 81.6816, 81.68089, 81.68125, 81.68063, 81.68119, 
    81.68022, 81.68002, 81.68015, 81.6796, 81.68122, 81.6806, 81.68528, 
    81.68525, 81.68512, 81.6857, 81.68573, 81.68624, 81.68578, 81.68559, 
    81.68508, 81.68479, 81.68452, 81.6839, 81.68323, 81.68227, 81.68156, 
    81.6811, 81.68138, 81.68113, 81.68141, 81.68154, 81.68009, 81.68091, 
    81.67967, 81.67974, 81.68031, 81.67973, 81.68523, 81.68539, 81.68594, 
    81.68551, 81.68629, 81.68586, 81.68562, 81.68464, 81.68442, 81.68422, 
    81.68383, 81.68333, 81.68245, 81.68168, 81.68097, 81.68102, 81.681, 
    81.68085, 81.68124, 81.68079, 81.68071, 81.68091, 81.67975, 81.68008, 
    81.67974, 81.67995, 81.68533, 81.68507, 81.68522, 81.68495, 81.68514, 
    81.6843, 81.68405, 81.68286, 81.68334, 81.68256, 81.68326, 81.68314, 
    81.68256, 81.68321, 81.68173, 81.68275, 81.68084, 81.68188, 81.68078, 
    81.68097, 81.68064, 81.68036, 81.67999, 81.67932, 81.67947, 81.6789, 
    81.68468, 81.68434, 81.68436, 81.684, 81.68374, 81.68315, 81.68223, 
    81.68257, 81.68192, 81.6818, 81.68278, 81.68218, 81.6841, 81.68381, 
    81.68398, 81.68465, 81.6825, 81.68362, 81.68156, 81.68215, 81.6804, 
    81.68128, 81.67956, 81.67885, 81.67813, 81.67735, 81.68414, 81.68437, 
    81.68395, 81.68339, 81.68284, 81.68212, 81.68204, 81.68191, 81.68156, 
    81.68127, 81.68188, 81.68119, 81.68375, 81.6824, 81.68447, 81.68386, 
    81.68342, 81.6836, 81.68261, 81.68237, 81.68144, 81.68192, 81.67903, 
    81.68031, 81.67671, 81.67773, 81.68446, 81.68414, 81.68305, 81.68357, 
    81.68207, 81.6817, 81.6814, 81.68102, 81.68097, 81.68075, 81.68111, 
    81.68076, 81.68212, 81.68151, 81.68317, 81.68277, 81.68295, 81.68315, 
    81.68253, 81.68187, 81.68184, 81.68163, 81.68108, 81.68206, 81.67889, 
    81.68088, 81.6838, 81.6832, 81.68311, 81.68333, 81.68174, 81.68232, 
    81.68075, 81.68118, 81.68048, 81.68082, 81.68088, 81.68132, 81.68159, 
    81.6823, 81.68286, 81.6833, 81.6832, 81.68272, 81.68182, 81.68098, 
    81.68117, 81.68053, 81.68217, 81.6815, 81.68176, 81.68106, 81.68259, 
    81.68134, 81.68291, 81.68277, 81.68233, 81.68146, 81.68124, 81.68104, 
    81.68116, 81.6818, 81.6819, 81.68233, 81.68246, 81.6828, 81.68307, 
    81.68282, 81.68256, 81.68179, 81.68111, 81.68036, 81.68017, 81.67932, 
    81.68003, 81.67889, 81.67989, 81.67813, 81.68124, 81.67989, 81.6823, 
    81.68204, 81.68158, 81.68049, 81.68106, 81.68039, 81.6819, 81.68271, 
    81.68289, 81.68327, 81.68288, 81.68291, 81.68254, 81.68266, 81.68177, 
    81.68224, 81.68089, 81.68039, 81.67897, 81.67811, 81.67721, 81.67682, 
    81.6767, 81.67664 ;

 RH2M_R =
  81.68618, 81.68539, 81.68554, 81.6849, 81.68525, 81.68484, 81.68601, 
    81.68536, 81.68578, 81.6861, 81.68369, 81.68487, 81.6824, 81.68316, 
    81.68121, 81.68252, 81.68095, 81.68124, 81.68033, 81.68059, 81.67946, 
    81.68021, 81.67885, 81.67963, 81.67951, 81.68024, 81.68462, 81.68384, 
    81.68467, 81.68456, 81.6846, 81.68524, 81.68558, 81.68623, 81.68611, 
    81.68562, 81.6845, 81.68488, 81.68391, 81.68393, 81.68287, 81.68335, 
    81.68155, 81.68206, 81.68057, 81.68095, 81.6806, 81.6807, 81.6806, 
    81.68114, 81.68091, 81.68139, 81.68327, 81.68272, 81.68435, 81.68536, 
    81.68599, 81.68645, 81.68638, 81.68626, 81.68562, 81.68501, 81.68455, 
    81.68424, 81.68394, 81.68305, 81.68256, 81.68146, 81.68164, 81.68132, 
    81.68098, 81.68046, 81.68054, 81.68031, 81.68131, 81.68065, 81.68175, 
    81.68145, 81.68391, 81.68478, 81.68519, 81.68551, 81.68633, 81.68577, 
    81.68599, 81.68545, 81.6851, 81.68527, 81.68423, 81.68464, 81.68253, 
    81.68343, 81.68103, 81.6816, 81.68089, 81.68125, 81.68063, 81.68119, 
    81.68022, 81.68002, 81.68015, 81.6796, 81.68122, 81.6806, 81.68528, 
    81.68525, 81.68512, 81.6857, 81.68573, 81.68624, 81.68578, 81.68559, 
    81.68508, 81.68479, 81.68452, 81.6839, 81.68323, 81.68227, 81.68156, 
    81.6811, 81.68138, 81.68113, 81.68141, 81.68154, 81.68009, 81.68091, 
    81.67967, 81.67974, 81.68031, 81.67973, 81.68523, 81.68539, 81.68594, 
    81.68551, 81.68629, 81.68586, 81.68562, 81.68464, 81.68442, 81.68422, 
    81.68383, 81.68333, 81.68245, 81.68168, 81.68097, 81.68102, 81.681, 
    81.68085, 81.68124, 81.68079, 81.68071, 81.68091, 81.67975, 81.68008, 
    81.67974, 81.67995, 81.68533, 81.68507, 81.68522, 81.68495, 81.68514, 
    81.6843, 81.68405, 81.68286, 81.68334, 81.68256, 81.68326, 81.68314, 
    81.68256, 81.68321, 81.68173, 81.68275, 81.68084, 81.68188, 81.68078, 
    81.68097, 81.68064, 81.68036, 81.67999, 81.67932, 81.67947, 81.6789, 
    81.68468, 81.68434, 81.68436, 81.684, 81.68374, 81.68315, 81.68223, 
    81.68257, 81.68192, 81.6818, 81.68278, 81.68218, 81.6841, 81.68381, 
    81.68398, 81.68465, 81.6825, 81.68362, 81.68156, 81.68215, 81.6804, 
    81.68128, 81.67956, 81.67885, 81.67813, 81.67735, 81.68414, 81.68437, 
    81.68395, 81.68339, 81.68284, 81.68212, 81.68204, 81.68191, 81.68156, 
    81.68127, 81.68188, 81.68119, 81.68375, 81.6824, 81.68447, 81.68386, 
    81.68342, 81.6836, 81.68261, 81.68237, 81.68144, 81.68192, 81.67903, 
    81.68031, 81.67671, 81.67773, 81.68446, 81.68414, 81.68305, 81.68357, 
    81.68207, 81.6817, 81.6814, 81.68102, 81.68097, 81.68075, 81.68111, 
    81.68076, 81.68212, 81.68151, 81.68317, 81.68277, 81.68295, 81.68315, 
    81.68253, 81.68187, 81.68184, 81.68163, 81.68108, 81.68206, 81.67889, 
    81.68088, 81.6838, 81.6832, 81.68311, 81.68333, 81.68174, 81.68232, 
    81.68075, 81.68118, 81.68048, 81.68082, 81.68088, 81.68132, 81.68159, 
    81.6823, 81.68286, 81.6833, 81.6832, 81.68272, 81.68182, 81.68098, 
    81.68117, 81.68053, 81.68217, 81.6815, 81.68176, 81.68106, 81.68259, 
    81.68134, 81.68291, 81.68277, 81.68233, 81.68146, 81.68124, 81.68104, 
    81.68116, 81.6818, 81.6819, 81.68233, 81.68246, 81.6828, 81.68307, 
    81.68282, 81.68256, 81.68179, 81.68111, 81.68036, 81.68017, 81.67932, 
    81.68003, 81.67889, 81.67989, 81.67813, 81.68124, 81.67989, 81.6823, 
    81.68204, 81.68158, 81.68049, 81.68106, 81.68039, 81.6819, 81.68271, 
    81.68289, 81.68327, 81.68288, 81.68291, 81.68254, 81.68266, 81.68177, 
    81.68224, 81.68089, 81.68039, 81.67897, 81.67811, 81.67721, 81.67682, 
    81.6767, 81.67664 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004365606, 0.0004384049, 0.0004380463, 0.0004395339, 0.0004387087, 
    0.0004396826, 0.0004369343, 0.0004384778, 0.0004374924, 0.0004367262, 
    0.0004424202, 0.0004395998, 0.0004453503, 0.0004435513, 0.0004480703, 
    0.0004450702, 0.0004486752, 0.0004479837, 0.0004500649, 0.0004494686, 
    0.0004521304, 0.00045034, 0.0004535103, 0.0004517028, 0.0004519854, 
    0.0004502806, 0.0004401679, 0.0004420695, 0.0004400551, 0.0004403263, 
    0.0004402045, 0.0004387254, 0.0004379801, 0.0004364192, 0.0004367025, 
    0.0004378489, 0.0004404478, 0.0004395655, 0.000441789, 0.0004417388, 
    0.0004442141, 0.000443098, 0.0004472587, 0.0004460761, 0.0004494934, 
    0.0004486339, 0.0004494529, 0.0004492045, 0.000449456, 0.0004481956, 
    0.0004487355, 0.0004476264, 0.0004433077, 0.0004445771, 0.0004407907, 
    0.0004385138, 0.0004370017, 0.0004359287, 0.0004360803, 0.0004363695, 
    0.0004378555, 0.0004392526, 0.0004403175, 0.0004410296, 0.0004417314, 
    0.0004438556, 0.00044498, 0.0004474977, 0.0004470434, 0.000447813, 
    0.0004485483, 0.0004497828, 0.0004495796, 0.0004501234, 0.0004477924, 
    0.0004493415, 0.0004467841, 0.0004474835, 0.0004419225, 0.0004398038, 
    0.000438903, 0.0004381147, 0.0004361969, 0.0004375213, 0.0004369991, 
    0.0004382411, 0.0004390304, 0.00043864, 0.0004410491, 0.0004401123, 
    0.0004450466, 0.0004429212, 0.0004484626, 0.0004471365, 0.0004487803, 
    0.0004479415, 0.0004493786, 0.0004480851, 0.0004503258, 0.0004508137, 
    0.0004504801, 0.000451761, 0.0004480131, 0.0004494523, 0.0004386293, 
    0.000438693, 0.0004389895, 0.0004376856, 0.0004376059, 0.000436411, 
    0.0004374741, 0.0004379268, 0.000439076, 0.0004397556, 0.0004404018, 
    0.0004418226, 0.0004434093, 0.0004456282, 0.0004472224, 0.0004482909, 
    0.0004476357, 0.0004482141, 0.0004475673, 0.0004472641, 0.0004506307, 
    0.0004487403, 0.0004515766, 0.0004514197, 0.0004501359, 0.0004514372, 
    0.0004387376, 0.0004383711, 0.0004370991, 0.0004380945, 0.0004362808, 
    0.000437296, 0.0004378796, 0.0004401318, 0.0004406266, 0.0004410855, 
    0.0004419917, 0.0004431547, 0.000445195, 0.0004469702, 0.0004485909, 
    0.0004484721, 0.0004485138, 0.0004488758, 0.000447979, 0.0004490229, 
    0.000449198, 0.0004487399, 0.0004513985, 0.000450639, 0.0004514162, 
    0.0004509215, 0.0004384902, 0.0004391065, 0.0004387734, 0.0004393997, 
    0.0004389583, 0.0004409205, 0.0004415087, 0.0004442616, 0.0004431318, 
    0.0004449299, 0.0004433143, 0.0004436006, 0.0004449883, 0.0004434015, 
    0.0004468721, 0.000444519, 0.0004488898, 0.0004465398, 0.0004490369, 
    0.0004485834, 0.0004493341, 0.0004500065, 0.0004508523, 0.000452413, 
    0.0004520515, 0.0004533568, 0.0004400255, 0.0004408249, 0.0004407545, 
    0.0004415912, 0.0004422099, 0.0004435513, 0.0004457025, 0.0004448934, 
    0.0004463785, 0.0004466767, 0.0004444203, 0.0004458056, 0.0004413595, 
    0.0004420776, 0.00044165, 0.0004400877, 0.0004450793, 0.0004425174, 
    0.0004472481, 0.0004458601, 0.0004499104, 0.0004478961, 0.0004518525, 
    0.0004535438, 0.0004551358, 0.0004569959, 0.0004412612, 0.0004407179, 
    0.0004416906, 0.0004430364, 0.0004442852, 0.0004459455, 0.0004461153, 
    0.0004464262, 0.0004472318, 0.0004479092, 0.0004465244, 0.0004480789, 
    0.0004422441, 0.0004453017, 0.0004405117, 0.000441954, 0.0004429564, 
    0.0004425167, 0.0004448003, 0.0004453384, 0.0004475255, 0.0004463949, 
    0.0004531262, 0.000450148, 0.0004584124, 0.0004561027, 0.000440528, 
    0.0004412592, 0.000443804, 0.0004425932, 0.0004460561, 0.0004469086, 
    0.0004476015, 0.0004484873, 0.0004485828, 0.0004491077, 0.0004482475, 
    0.0004490736, 0.0004459484, 0.0004473449, 0.0004435126, 0.0004444452, 
    0.0004440162, 0.0004435454, 0.000444998, 0.0004465455, 0.0004465786, 
    0.0004470747, 0.0004484729, 0.0004460692, 0.0004535102, 0.0004489145, 
    0.0004420565, 0.0004434648, 0.000443666, 0.0004431204, 0.000446823, 
    0.0004454813, 0.0004490949, 0.0004481182, 0.0004497183, 0.0004489232, 
    0.000448806, 0.0004477848, 0.0004471488, 0.0004455424, 0.0004442353, 
    0.0004431989, 0.0004434398, 0.0004445782, 0.0004466401, 0.0004485908, 
    0.0004481634, 0.000449596, 0.0004458039, 0.0004473939, 0.0004467792, 
    0.0004483818, 0.0004448717, 0.0004478614, 0.0004441074, 0.0004444365, 
    0.0004454546, 0.0004475026, 0.0004479557, 0.0004484394, 0.0004481408, 
    0.0004466928, 0.0004464556, 0.0004454295, 0.0004451461, 0.0004443643, 
    0.000443717, 0.0004443083, 0.0004449292, 0.000446693, 0.0004482825, 
    0.0004500154, 0.0004504395, 0.000452464, 0.0004508157, 0.0004535355, 
    0.000451223, 0.0004552261, 0.0004480347, 0.0004511562, 0.0004455009, 
    0.0004461101, 0.000447212, 0.0004497394, 0.0004483749, 0.0004499706, 
    0.0004464462, 0.0004446176, 0.0004441445, 0.0004432618, 0.0004441646, 
    0.0004440912, 0.000444955, 0.0004446773, 0.0004467515, 0.0004456373, 
    0.0004488023, 0.0004499574, 0.0004532194, 0.000455219, 0.0004572547, 
    0.0004581533, 0.0004584268, 0.0004585411 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.502156e-14, 3.511612e-14, 3.509775e-14, 3.517395e-14, 3.51317e-14, 
    3.518158e-14, 3.504075e-14, 3.511986e-14, 3.506937e-14, 3.503009e-14, 
    3.532161e-14, 3.517735e-14, 3.54713e-14, 3.537948e-14, 3.561e-14, 
    3.545701e-14, 3.564082e-14, 3.560561e-14, 3.571158e-14, 3.568124e-14, 
    3.581657e-14, 3.572558e-14, 3.588667e-14, 3.579486e-14, 3.580922e-14, 
    3.572257e-14, 3.520643e-14, 3.530365e-14, 3.520066e-14, 3.521453e-14, 
    3.520831e-14, 3.513257e-14, 3.509435e-14, 3.501434e-14, 3.502888e-14, 
    3.508765e-14, 3.522077e-14, 3.517562e-14, 3.528942e-14, 3.528685e-14, 
    3.541334e-14, 3.535633e-14, 3.556868e-14, 3.550838e-14, 3.568251e-14, 
    3.563875e-14, 3.568045e-14, 3.566781e-14, 3.568061e-14, 3.561643e-14, 
    3.564393e-14, 3.558744e-14, 3.536701e-14, 3.543184e-14, 3.523831e-14, 
    3.512169e-14, 3.504422e-14, 3.498917e-14, 3.499696e-14, 3.501179e-14, 
    3.508799e-14, 3.51596e-14, 3.521413e-14, 3.525058e-14, 3.528648e-14, 
    3.539499e-14, 3.545243e-14, 3.558085e-14, 3.555771e-14, 3.559692e-14, 
    3.563439e-14, 3.569724e-14, 3.56869e-14, 3.571458e-14, 3.55959e-14, 
    3.567478e-14, 3.554452e-14, 3.558017e-14, 3.529614e-14, 3.518781e-14, 
    3.514164e-14, 3.510128e-14, 3.500294e-14, 3.507086e-14, 3.504409e-14, 
    3.510778e-14, 3.514822e-14, 3.512822e-14, 3.525157e-14, 3.520363e-14, 
    3.545583e-14, 3.534729e-14, 3.563002e-14, 3.556246e-14, 3.564621e-14, 
    3.560349e-14, 3.567667e-14, 3.561081e-14, 3.572488e-14, 3.574968e-14, 
    3.573273e-14, 3.579786e-14, 3.560716e-14, 3.568044e-14, 3.512766e-14, 
    3.513092e-14, 3.514612e-14, 3.507929e-14, 3.50752e-14, 3.501394e-14, 
    3.506846e-14, 3.509166e-14, 3.515057e-14, 3.518537e-14, 3.521845e-14, 
    3.529114e-14, 3.537223e-14, 3.548553e-14, 3.556684e-14, 3.56213e-14, 
    3.558792e-14, 3.561739e-14, 3.558444e-14, 3.556899e-14, 3.574038e-14, 
    3.564418e-14, 3.57885e-14, 3.578052e-14, 3.571523e-14, 3.578142e-14, 
    3.513321e-14, 3.511445e-14, 3.504923e-14, 3.510027e-14, 3.500727e-14, 
    3.505933e-14, 3.508924e-14, 3.520462e-14, 3.522997e-14, 3.525344e-14, 
    3.52998e-14, 3.535925e-14, 3.546343e-14, 3.555398e-14, 3.563658e-14, 
    3.563053e-14, 3.563266e-14, 3.565109e-14, 3.560542e-14, 3.565859e-14, 
    3.56675e-14, 3.564418e-14, 3.577945e-14, 3.574083e-14, 3.578035e-14, 
    3.575521e-14, 3.512055e-14, 3.515212e-14, 3.513506e-14, 3.516714e-14, 
    3.514454e-14, 3.524498e-14, 3.527507e-14, 3.541577e-14, 3.535808e-14, 
    3.544989e-14, 3.536741e-14, 3.538203e-14, 3.545285e-14, 3.537188e-14, 
    3.554898e-14, 3.542891e-14, 3.565181e-14, 3.553202e-14, 3.56593e-14, 
    3.563622e-14, 3.567445e-14, 3.570865e-14, 3.575169e-14, 3.5831e-14, 
    3.581264e-14, 3.587894e-14, 3.519919e-14, 3.524009e-14, 3.523651e-14, 
    3.527932e-14, 3.531095e-14, 3.537951e-14, 3.548933e-14, 3.544806e-14, 
    3.552383e-14, 3.553903e-14, 3.542391e-14, 3.54946e-14, 3.526748e-14, 
    3.530419e-14, 3.528235e-14, 3.52024e-14, 3.545754e-14, 3.532669e-14, 
    3.556818e-14, 3.549742e-14, 3.570377e-14, 3.560119e-14, 3.580253e-14, 
    3.58884e-14, 3.596922e-14, 3.606345e-14, 3.526243e-14, 3.523464e-14, 
    3.528441e-14, 3.535318e-14, 3.5417e-14, 3.550173e-14, 3.55104e-14, 
    3.552626e-14, 3.556734e-14, 3.560186e-14, 3.553126e-14, 3.561052e-14, 
    3.531267e-14, 3.54689e-14, 3.522412e-14, 3.529788e-14, 3.534914e-14, 
    3.532667e-14, 3.544334e-14, 3.547081e-14, 3.558233e-14, 3.552471e-14, 
    3.58672e-14, 3.571585e-14, 3.613519e-14, 3.601822e-14, 3.522493e-14, 
    3.526234e-14, 3.539242e-14, 3.533056e-14, 3.550739e-14, 3.555086e-14, 
    3.558619e-14, 3.56313e-14, 3.563618e-14, 3.56629e-14, 3.561911e-14, 
    3.566117e-14, 3.550191e-14, 3.557312e-14, 3.537758e-14, 3.542521e-14, 
    3.540331e-14, 3.537927e-14, 3.545344e-14, 3.553236e-14, 3.553408e-14, 
    3.555936e-14, 3.563053e-14, 3.550811e-14, 3.588667e-14, 3.565304e-14, 
    3.530313e-14, 3.537508e-14, 3.538539e-14, 3.535752e-14, 3.55465e-14, 
    3.547807e-14, 3.566225e-14, 3.561252e-14, 3.5694e-14, 3.565352e-14, 
    3.564756e-14, 3.559554e-14, 3.556313e-14, 3.54812e-14, 3.541449e-14, 
    3.536157e-14, 3.537387e-14, 3.5432e-14, 3.55372e-14, 3.563661e-14, 
    3.561484e-14, 3.568781e-14, 3.549458e-14, 3.557564e-14, 3.554431e-14, 
    3.562599e-14, 3.544695e-14, 3.559935e-14, 3.540795e-14, 3.542475e-14, 
    3.547671e-14, 3.558112e-14, 3.560425e-14, 3.562888e-14, 3.561369e-14, 
    3.553987e-14, 3.552778e-14, 3.547545e-14, 3.546099e-14, 3.54211e-14, 
    3.538804e-14, 3.541823e-14, 3.544992e-14, 3.553991e-14, 3.562091e-14, 
    3.570914e-14, 3.573072e-14, 3.583358e-14, 3.574982e-14, 3.588796e-14, 
    3.577047e-14, 3.597376e-14, 3.560821e-14, 3.576707e-14, 3.547908e-14, 
    3.551017e-14, 3.556632e-14, 3.569504e-14, 3.562561e-14, 3.570682e-14, 
    3.552731e-14, 3.543399e-14, 3.540987e-14, 3.536478e-14, 3.54109e-14, 
    3.540715e-14, 3.545126e-14, 3.543709e-14, 3.55429e-14, 3.548608e-14, 
    3.56474e-14, 3.570618e-14, 3.587199e-14, 3.597344e-14, 3.607662e-14, 
    3.612212e-14, 3.613596e-14, 3.614175e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.164501e-14, 1.167648e-14, 1.167037e-14, 1.169573e-14, 1.168167e-14, 
    1.169827e-14, 1.16514e-14, 1.167773e-14, 1.166092e-14, 1.164785e-14, 
    1.174488e-14, 1.169687e-14, 1.179471e-14, 1.176414e-14, 1.184087e-14, 
    1.178995e-14, 1.185113e-14, 1.183941e-14, 1.187469e-14, 1.186459e-14, 
    1.190963e-14, 1.187935e-14, 1.193297e-14, 1.190241e-14, 1.190719e-14, 
    1.187835e-14, 1.170654e-14, 1.17389e-14, 1.170462e-14, 1.170924e-14, 
    1.170717e-14, 1.168196e-14, 1.166924e-14, 1.164261e-14, 1.164745e-14, 
    1.166701e-14, 1.171132e-14, 1.169629e-14, 1.173417e-14, 1.173331e-14, 
    1.177541e-14, 1.175644e-14, 1.182712e-14, 1.180705e-14, 1.186501e-14, 
    1.185044e-14, 1.186432e-14, 1.186012e-14, 1.186438e-14, 1.184301e-14, 
    1.185217e-14, 1.183336e-14, 1.175999e-14, 1.178157e-14, 1.171715e-14, 
    1.167834e-14, 1.165255e-14, 1.163423e-14, 1.163682e-14, 1.164176e-14, 
    1.166712e-14, 1.169096e-14, 1.17091e-14, 1.172124e-14, 1.173319e-14, 
    1.176931e-14, 1.178842e-14, 1.183117e-14, 1.182347e-14, 1.183652e-14, 
    1.184899e-14, 1.186991e-14, 1.186647e-14, 1.187568e-14, 1.183618e-14, 
    1.186244e-14, 1.181908e-14, 1.183094e-14, 1.17364e-14, 1.170035e-14, 
    1.168498e-14, 1.167154e-14, 1.163881e-14, 1.166142e-14, 1.165251e-14, 
    1.167371e-14, 1.168717e-14, 1.168051e-14, 1.172157e-14, 1.170561e-14, 
    1.178956e-14, 1.175343e-14, 1.184754e-14, 1.182505e-14, 1.185293e-14, 
    1.183871e-14, 1.186307e-14, 1.184114e-14, 1.187911e-14, 1.188737e-14, 
    1.188173e-14, 1.190341e-14, 1.183993e-14, 1.186432e-14, 1.168033e-14, 
    1.168141e-14, 1.168647e-14, 1.166422e-14, 1.166286e-14, 1.164247e-14, 
    1.166062e-14, 1.166834e-14, 1.168795e-14, 1.169954e-14, 1.171055e-14, 
    1.173474e-14, 1.176173e-14, 1.179944e-14, 1.182651e-14, 1.184463e-14, 
    1.183352e-14, 1.184333e-14, 1.183237e-14, 1.182722e-14, 1.188427e-14, 
    1.185225e-14, 1.190029e-14, 1.189763e-14, 1.18759e-14, 1.189793e-14, 
    1.168217e-14, 1.167593e-14, 1.165422e-14, 1.167121e-14, 1.164025e-14, 
    1.165758e-14, 1.166754e-14, 1.170594e-14, 1.171438e-14, 1.172219e-14, 
    1.173762e-14, 1.175741e-14, 1.179209e-14, 1.182223e-14, 1.184972e-14, 
    1.184771e-14, 1.184842e-14, 1.185455e-14, 1.183935e-14, 1.185705e-14, 
    1.186001e-14, 1.185225e-14, 1.189728e-14, 1.188442e-14, 1.189758e-14, 
    1.188921e-14, 1.167796e-14, 1.168847e-14, 1.168279e-14, 1.169347e-14, 
    1.168594e-14, 1.171937e-14, 1.172939e-14, 1.177622e-14, 1.175702e-14, 
    1.178758e-14, 1.176013e-14, 1.176499e-14, 1.178856e-14, 1.176161e-14, 
    1.182056e-14, 1.17806e-14, 1.185479e-14, 1.181492e-14, 1.185729e-14, 
    1.18496e-14, 1.186233e-14, 1.187371e-14, 1.188804e-14, 1.191444e-14, 
    1.190833e-14, 1.193039e-14, 1.170413e-14, 1.171775e-14, 1.171656e-14, 
    1.17308e-14, 1.174133e-14, 1.176415e-14, 1.180071e-14, 1.178697e-14, 
    1.181219e-14, 1.181725e-14, 1.177893e-14, 1.180246e-14, 1.172686e-14, 
    1.173908e-14, 1.173181e-14, 1.17052e-14, 1.179013e-14, 1.174657e-14, 
    1.182695e-14, 1.18034e-14, 1.187209e-14, 1.183794e-14, 1.190496e-14, 
    1.193354e-14, 1.196044e-14, 1.199181e-14, 1.172518e-14, 1.171593e-14, 
    1.17325e-14, 1.175539e-14, 1.177663e-14, 1.180484e-14, 1.180772e-14, 
    1.1813e-14, 1.182668e-14, 1.183816e-14, 1.181466e-14, 1.184104e-14, 
    1.174191e-14, 1.179391e-14, 1.171243e-14, 1.173698e-14, 1.175404e-14, 
    1.174657e-14, 1.17854e-14, 1.179454e-14, 1.183166e-14, 1.181248e-14, 
    1.192649e-14, 1.187611e-14, 1.201569e-14, 1.197676e-14, 1.17127e-14, 
    1.172515e-14, 1.176845e-14, 1.174786e-14, 1.180672e-14, 1.182119e-14, 
    1.183295e-14, 1.184796e-14, 1.184959e-14, 1.185848e-14, 1.184391e-14, 
    1.185791e-14, 1.180489e-14, 1.18286e-14, 1.176351e-14, 1.177936e-14, 
    1.177207e-14, 1.176407e-14, 1.178876e-14, 1.181503e-14, 1.18156e-14, 
    1.182402e-14, 1.184771e-14, 1.180696e-14, 1.193296e-14, 1.18552e-14, 
    1.173873e-14, 1.176268e-14, 1.176611e-14, 1.175683e-14, 1.181974e-14, 
    1.179696e-14, 1.185827e-14, 1.184171e-14, 1.186883e-14, 1.185536e-14, 
    1.185337e-14, 1.183606e-14, 1.182527e-14, 1.1798e-14, 1.17758e-14, 
    1.175818e-14, 1.176228e-14, 1.178163e-14, 1.181664e-14, 1.184973e-14, 
    1.184248e-14, 1.186677e-14, 1.180246e-14, 1.182944e-14, 1.181901e-14, 
    1.18462e-14, 1.17866e-14, 1.183733e-14, 1.177362e-14, 1.177921e-14, 
    1.179651e-14, 1.183126e-14, 1.183896e-14, 1.184716e-14, 1.18421e-14, 
    1.181753e-14, 1.181351e-14, 1.179609e-14, 1.179127e-14, 1.177799e-14, 
    1.176699e-14, 1.177704e-14, 1.178759e-14, 1.181755e-14, 1.184451e-14, 
    1.187387e-14, 1.188106e-14, 1.19153e-14, 1.188741e-14, 1.193339e-14, 
    1.189429e-14, 1.196196e-14, 1.184028e-14, 1.189316e-14, 1.17973e-14, 
    1.180764e-14, 1.182634e-14, 1.186918e-14, 1.184607e-14, 1.18731e-14, 
    1.181335e-14, 1.178229e-14, 1.177426e-14, 1.175925e-14, 1.17746e-14, 
    1.177335e-14, 1.178804e-14, 1.178332e-14, 1.181854e-14, 1.179963e-14, 
    1.185332e-14, 1.187289e-14, 1.192808e-14, 1.196185e-14, 1.19962e-14, 
    1.201134e-14, 1.201595e-14, 1.201787e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.152213e-11, -8.188185e-11, -8.181192e-11, -8.210205e-11, -8.194111e-11, 
    -8.213109e-11, -8.159506e-11, -8.189612e-11, -8.170394e-11, 
    -8.155453e-11, -8.266511e-11, -8.2115e-11, -8.323666e-11, -8.288577e-11, 
    -8.376728e-11, -8.318205e-11, -8.388529e-11, -8.375042e-11, 
    -8.415642e-11, -8.404011e-11, -8.45594e-11, -8.421011e-11, -8.482864e-11, 
    -8.4476e-11, -8.453115e-11, -8.419859e-11, -8.222572e-11, -8.259662e-11, 
    -8.220374e-11, -8.225663e-11, -8.22329e-11, -8.194444e-11, -8.179905e-11, 
    -8.149465e-11, -8.154992e-11, -8.17735e-11, -8.228041e-11, -8.210835e-11, 
    -8.254204e-11, -8.253224e-11, -8.301509e-11, -8.279739e-11, 
    -8.360901e-11, -8.337833e-11, -8.404497e-11, -8.387731e-11, 
    -8.403709e-11, -8.398864e-11, -8.403772e-11, -8.379183e-11, 
    -8.389717e-11, -8.368082e-11, -8.283815e-11, -8.308579e-11, 
    -8.234723e-11, -8.190316e-11, -8.160827e-11, -8.1399e-11, -8.142858e-11, 
    -8.148498e-11, -8.177481e-11, -8.204733e-11, -8.225502e-11, 
    -8.239395e-11, -8.253084e-11, -8.294516e-11, -8.316452e-11, 
    -8.365564e-11, -8.356703e-11, -8.371717e-11, -8.386063e-11, 
    -8.410147e-11, -8.406183e-11, -8.416794e-11, -8.371322e-11, 
    -8.401541e-11, -8.351654e-11, -8.365298e-11, -8.256799e-11, 
    -8.215477e-11, -8.197908e-11, -8.182536e-11, -8.145132e-11, 
    -8.170962e-11, -8.16078e-11, -8.185005e-11, -8.200399e-11, -8.192786e-11, 
    -8.239775e-11, -8.221506e-11, -8.317751e-11, -8.276294e-11, 
    -8.384389e-11, -8.358522e-11, -8.39059e-11, -8.374226e-11, -8.402264e-11, 
    -8.37703e-11, -8.420743e-11, -8.430261e-11, -8.423757e-11, -8.448745e-11, 
    -8.375631e-11, -8.403708e-11, -8.192572e-11, -8.193814e-11, 
    -8.199599e-11, -8.17417e-11, -8.172614e-11, -8.149313e-11, -8.170047e-11, 
    -8.178876e-11, -8.201292e-11, -8.21455e-11, -8.227154e-11, -8.254866e-11, 
    -8.285816e-11, -8.3291e-11, -8.360198e-11, -8.381044e-11, -8.368262e-11, 
    -8.379547e-11, -8.366931e-11, -8.36102e-11, -8.426694e-11, -8.389816e-11, 
    -8.445151e-11, -8.442089e-11, -8.417046e-11, -8.442434e-11, 
    -8.194686e-11, -8.187541e-11, -8.162732e-11, -8.182147e-11, 
    -8.146776e-11, -8.166574e-11, -8.177958e-11, -8.221886e-11, -8.23154e-11, 
    -8.24049e-11, -8.258166e-11, -8.280852e-11, -8.320651e-11, -8.355282e-11, 
    -8.386897e-11, -8.384581e-11, -8.385397e-11, -8.392459e-11, 
    -8.374965e-11, -8.395331e-11, -8.398748e-11, -8.389812e-11, 
    -8.441679e-11, -8.426861e-11, -8.442024e-11, -8.432376e-11, 
    -8.189863e-11, -8.201886e-11, -8.19539e-11, -8.207606e-11, -8.198999e-11, 
    -8.23727e-11, -8.248745e-11, -8.302442e-11, -8.280406e-11, -8.31548e-11, 
    -8.283969e-11, -8.289552e-11, -8.316621e-11, -8.285672e-11, 
    -8.353371e-11, -8.307471e-11, -8.392733e-11, -8.346892e-11, 
    -8.395606e-11, -8.386761e-11, -8.401406e-11, -8.414523e-11, 
    -8.431025e-11, -8.461474e-11, -8.454423e-11, -8.479888e-11, -8.21981e-11, 
    -8.235405e-11, -8.234033e-11, -8.250353e-11, -8.262423e-11, 
    -8.288587e-11, -8.33055e-11, -8.31477e-11, -8.343741e-11, -8.349556e-11, 
    -8.305544e-11, -8.332566e-11, -8.245842e-11, -8.259852e-11, 
    -8.251511e-11, -8.221041e-11, -8.318405e-11, -8.268435e-11, 
    -8.360712e-11, -8.33364e-11, -8.412652e-11, -8.373355e-11, -8.450542e-11, 
    -8.483537e-11, -8.514598e-11, -8.550892e-11, -8.243917e-11, 
    -8.233321e-11, -8.252295e-11, -8.278545e-11, -8.302906e-11, 
    -8.335291e-11, -8.338605e-11, -8.344672e-11, -8.360389e-11, 
    -8.373603e-11, -8.346589e-11, -8.376915e-11, -8.263099e-11, 
    -8.322742e-11, -8.229314e-11, -8.257444e-11, -8.276999e-11, 
    -8.268421e-11, -8.312967e-11, -8.323466e-11, -8.366131e-11, 
    -8.344075e-11, -8.475393e-11, -8.417292e-11, -8.578532e-11, 
    -8.533468e-11, -8.229618e-11, -8.243881e-11, -8.293521e-11, 
    -8.269902e-11, -8.337454e-11, -8.354081e-11, -8.3676e-11, -8.38488e-11, 
    -8.386746e-11, -8.396984e-11, -8.380207e-11, -8.396322e-11, 
    -8.335359e-11, -8.362602e-11, -8.287848e-11, -8.306041e-11, 
    -8.297672e-11, -8.288491e-11, -8.316827e-11, -8.347014e-11, 
    -8.347661e-11, -8.357341e-11, -8.384615e-11, -8.337727e-11, 
    -8.482888e-11, -8.393234e-11, -8.259434e-11, -8.286905e-11, 
    -8.290831e-11, -8.280189e-11, -8.352415e-11, -8.326244e-11, 
    -8.396735e-11, -8.377683e-11, -8.4089e-11, -8.393387e-11, -8.391105e-11, 
    -8.371183e-11, -8.358779e-11, -8.327443e-11, -8.301948e-11, 
    -8.281733e-11, -8.286434e-11, -8.30864e-11, -8.348861e-11, -8.386914e-11, 
    -8.378578e-11, -8.406528e-11, -8.332555e-11, -8.363572e-11, 
    -8.351583e-11, -8.382843e-11, -8.314351e-11, -8.37267e-11, -8.299444e-11, 
    -8.305864e-11, -8.325724e-11, -8.365674e-11, -8.374516e-11, 
    -8.383953e-11, -8.378129e-11, -8.349883e-11, -8.345256e-11, 
    -8.325242e-11, -8.319715e-11, -8.304466e-11, -8.291841e-11, 
    -8.303376e-11, -8.315489e-11, -8.349895e-11, -8.380902e-11, 
    -8.414709e-11, -8.422983e-11, -8.462481e-11, -8.430326e-11, 
    -8.483387e-11, -8.438272e-11, -8.516374e-11, -8.376053e-11, 
    -8.436948e-11, -8.326628e-11, -8.338513e-11, -8.360008e-11, 
    -8.409313e-11, -8.382697e-11, -8.413825e-11, -8.345075e-11, 
    -8.309405e-11, -8.300179e-11, -8.282962e-11, -8.300573e-11, 
    -8.299141e-11, -8.315992e-11, -8.310577e-11, -8.351038e-11, 
    -8.329304e-11, -8.391048e-11, -8.41358e-11, -8.477219e-11, -8.516234e-11, 
    -8.555952e-11, -8.573487e-11, -8.578824e-11, -8.581056e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -1.964839e-12, -1.973507e-12, -1.971822e-12, -1.978813e-12, -1.974935e-12, 
    -1.979513e-12, -1.966597e-12, -1.973851e-12, -1.96922e-12, -1.96562e-12, 
    -1.992381e-12, -1.979125e-12, -2.006153e-12, -1.997698e-12, -2.01894e-12, 
    -2.004838e-12, -2.021783e-12, -2.018533e-12, -2.028317e-12, 
    -2.025514e-12, -2.038027e-12, -2.02961e-12, -2.044515e-12, -2.036017e-12, 
    -2.037346e-12, -2.029333e-12, -1.981793e-12, -1.99073e-12, -1.981264e-12, 
    -1.982538e-12, -1.981966e-12, -1.975015e-12, -1.971512e-12, 
    -1.964177e-12, -1.965509e-12, -1.970896e-12, -1.983111e-12, 
    -1.978965e-12, -1.989416e-12, -1.98918e-12, -2.000814e-12, -1.995568e-12, 
    -2.015126e-12, -2.009567e-12, -2.025631e-12, -2.021591e-12, 
    -2.025441e-12, -2.024274e-12, -2.025456e-12, -2.019531e-12, -2.02207e-12, 
    -2.016856e-12, -1.996551e-12, -2.002518e-12, -1.984721e-12, 
    -1.974021e-12, -1.966915e-12, -1.961872e-12, -1.962585e-12, 
    -1.963944e-12, -1.970928e-12, -1.977495e-12, -1.982499e-12, 
    -1.985847e-12, -1.989146e-12, -1.99913e-12, -2.004415e-12, -2.01625e-12, 
    -2.014114e-12, -2.017732e-12, -2.021189e-12, -2.026992e-12, 
    -2.026037e-12, -2.028594e-12, -2.017637e-12, -2.024919e-12, 
    -2.012898e-12, -2.016185e-12, -1.990041e-12, -1.980084e-12, -1.97585e-12, 
    -1.972146e-12, -1.963133e-12, -1.969357e-12, -1.966903e-12, 
    -1.972741e-12, -1.97645e-12, -1.974616e-12, -1.985939e-12, -1.981536e-12, 
    -2.004728e-12, -1.994738e-12, -2.020786e-12, -2.014553e-12, -2.02228e-12, 
    -2.018337e-12, -2.025093e-12, -2.019013e-12, -2.029546e-12, 
    -2.031839e-12, -2.030272e-12, -2.036293e-12, -2.018675e-12, 
    -2.025441e-12, -1.974564e-12, -1.974863e-12, -1.976257e-12, -1.97013e-12, 
    -1.969755e-12, -1.96414e-12, -1.969136e-12, -1.971264e-12, -1.976665e-12, 
    -1.97986e-12, -1.982897e-12, -1.989575e-12, -1.997033e-12, -2.007463e-12, 
    -2.014957e-12, -2.01998e-12, -2.0169e-12, -2.019619e-12, -2.016579e-12, 
    -2.015154e-12, -2.03098e-12, -2.022093e-12, -2.035427e-12, -2.034689e-12, 
    -2.028655e-12, -2.034773e-12, -1.975074e-12, -1.973352e-12, 
    -1.967374e-12, -1.972052e-12, -1.963529e-12, -1.9683e-12, -1.971043e-12, 
    -1.981628e-12, -1.983954e-12, -1.986111e-12, -1.99037e-12, -1.995837e-12, 
    -2.005427e-12, -2.013772e-12, -2.02139e-12, -2.020832e-12, -2.021029e-12, 
    -2.02273e-12, -2.018515e-12, -2.023422e-12, -2.024246e-12, -2.022092e-12, 
    -2.034591e-12, -2.03102e-12, -2.034674e-12, -2.032349e-12, -1.973911e-12, 
    -1.976809e-12, -1.975243e-12, -1.978187e-12, -1.976113e-12, 
    -1.985335e-12, -1.9881e-12, -2.001039e-12, -1.995729e-12, -2.004181e-12, 
    -1.996588e-12, -1.997933e-12, -2.004456e-12, -1.996998e-12, 
    -2.013311e-12, -2.002251e-12, -2.022796e-12, -2.01175e-12, -2.023489e-12, 
    -2.021357e-12, -2.024886e-12, -2.028047e-12, -2.032023e-12, -2.03936e-12, 
    -2.037661e-12, -2.043798e-12, -1.981128e-12, -1.984886e-12, 
    -1.984555e-12, -1.988488e-12, -1.991396e-12, -1.997701e-12, 
    -2.007812e-12, -2.00401e-12, -2.010991e-12, -2.012392e-12, -2.001787e-12, 
    -2.008298e-12, -1.987401e-12, -1.990776e-12, -1.988767e-12, 
    -1.981424e-12, -2.004886e-12, -1.992845e-12, -2.01508e-12, -2.008557e-12, 
    -2.027596e-12, -2.018127e-12, -2.036726e-12, -2.044677e-12, 
    -2.052161e-12, -2.060907e-12, -1.986937e-12, -1.984383e-12, 
    -1.988955e-12, -1.995281e-12, -2.001151e-12, -2.008955e-12, 
    -2.009753e-12, -2.011215e-12, -2.015002e-12, -2.018187e-12, 
    -2.011677e-12, -2.018985e-12, -1.991559e-12, -2.005931e-12, 
    -1.983418e-12, -1.990196e-12, -1.994908e-12, -1.992841e-12, 
    -2.003575e-12, -2.006105e-12, -2.016386e-12, -2.011072e-12, 
    -2.042714e-12, -2.028714e-12, -2.067567e-12, -2.056708e-12, 
    -1.983491e-12, -1.986928e-12, -1.99889e-12, -1.993198e-12, -2.009476e-12, 
    -2.013482e-12, -2.01674e-12, -2.020904e-12, -2.021354e-12, -2.023821e-12, 
    -2.019778e-12, -2.023661e-12, -2.008971e-12, -2.015536e-12, 
    -1.997523e-12, -2.001907e-12, -1.99989e-12, -1.997678e-12, -2.004506e-12, 
    -2.01178e-12, -2.011936e-12, -2.014268e-12, -2.02084e-12, -2.009542e-12, 
    -2.04452e-12, -2.022917e-12, -1.990676e-12, -1.997295e-12, -1.998241e-12, 
    -1.995677e-12, -2.013081e-12, -2.006775e-12, -2.023761e-12, -2.01917e-12, 
    -2.026692e-12, -2.022954e-12, -2.022404e-12, -2.017604e-12, 
    -2.014615e-12, -2.007064e-12, -2.00092e-12, -1.996049e-12, -1.997182e-12, 
    -2.002533e-12, -2.012225e-12, -2.021394e-12, -2.019386e-12, -2.02612e-12, 
    -2.008295e-12, -2.015769e-12, -2.012881e-12, -2.020413e-12, 
    -2.003909e-12, -2.017962e-12, -2.000317e-12, -2.001864e-12, 
    -2.006649e-12, -2.016276e-12, -2.018406e-12, -2.02068e-12, -2.019277e-12, 
    -2.012471e-12, -2.011356e-12, -2.006533e-12, -2.005202e-12, 
    -2.001527e-12, -1.998485e-12, -2.001264e-12, -2.004183e-12, 
    -2.012474e-12, -2.019945e-12, -2.028092e-12, -2.030086e-12, 
    -2.039603e-12, -2.031855e-12, -2.044641e-12, -2.033769e-12, 
    -2.052589e-12, -2.018777e-12, -2.03345e-12, -2.006867e-12, -2.009731e-12, 
    -2.014911e-12, -2.026791e-12, -2.020378e-12, -2.027879e-12, 
    -2.011312e-12, -2.002717e-12, -2.000494e-12, -1.996345e-12, 
    -2.000589e-12, -2.000244e-12, -2.004304e-12, -2.003e-12, -2.012749e-12, 
    -2.007512e-12, -2.02239e-12, -2.02782e-12, -2.043154e-12, -2.052555e-12, 
    -2.062126e-12, -2.066351e-12, -2.067638e-12, -2.068175e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.782927e-15, 3.793152e-15, 3.791166e-15, 3.799406e-15, 3.794837e-15, 
    3.80023e-15, 3.785003e-15, 3.793557e-15, 3.788098e-15, 3.78385e-15, 
    3.815371e-15, 3.799773e-15, 3.831558e-15, 3.821628e-15, 3.846554e-15, 
    3.830012e-15, 3.849887e-15, 3.846081e-15, 3.857539e-15, 3.854258e-15, 
    3.868892e-15, 3.859053e-15, 3.876472e-15, 3.866544e-15, 3.868097e-15, 
    3.858728e-15, 3.802917e-15, 3.81343e-15, 3.802294e-15, 3.803793e-15, 
    3.803121e-15, 3.79493e-15, 3.790798e-15, 3.782147e-15, 3.783719e-15, 
    3.790073e-15, 3.804468e-15, 3.799586e-15, 3.811891e-15, 3.811613e-15, 
    3.825291e-15, 3.819126e-15, 3.842086e-15, 3.835567e-15, 3.854395e-15, 
    3.849664e-15, 3.854173e-15, 3.852806e-15, 3.85419e-15, 3.84725e-15, 
    3.850224e-15, 3.844115e-15, 3.82028e-15, 3.827291e-15, 3.806364e-15, 
    3.793755e-15, 3.785378e-15, 3.779426e-15, 3.780267e-15, 3.781871e-15, 
    3.790111e-15, 3.797854e-15, 3.80375e-15, 3.807691e-15, 3.811573e-15, 
    3.823306e-15, 3.829517e-15, 3.843403e-15, 3.840901e-15, 3.845141e-15, 
    3.849193e-15, 3.855988e-15, 3.854871e-15, 3.857863e-15, 3.845031e-15, 
    3.85356e-15, 3.839475e-15, 3.843329e-15, 3.812618e-15, 3.800904e-15, 
    3.795912e-15, 3.791548e-15, 3.780915e-15, 3.788258e-15, 3.785364e-15, 
    3.792251e-15, 3.796623e-15, 3.794461e-15, 3.807798e-15, 3.802615e-15, 
    3.829885e-15, 3.818149e-15, 3.84872e-15, 3.841415e-15, 3.850471e-15, 
    3.845851e-15, 3.853764e-15, 3.846643e-15, 3.858977e-15, 3.861659e-15, 
    3.859826e-15, 3.866869e-15, 3.846248e-15, 3.854171e-15, 3.7944e-15, 
    3.794752e-15, 3.796396e-15, 3.78917e-15, 3.788728e-15, 3.782104e-15, 
    3.787999e-15, 3.790508e-15, 3.796877e-15, 3.800641e-15, 3.804218e-15, 
    3.812077e-15, 3.820846e-15, 3.833096e-15, 3.841888e-15, 3.847777e-15, 
    3.844167e-15, 3.847354e-15, 3.843791e-15, 3.842121e-15, 3.860654e-15, 
    3.850251e-15, 3.865856e-15, 3.864994e-15, 3.857934e-15, 3.865091e-15, 
    3.795e-15, 3.792971e-15, 3.78592e-15, 3.791438e-15, 3.781382e-15, 
    3.787011e-15, 3.790246e-15, 3.802721e-15, 3.805462e-15, 3.808001e-15, 
    3.813013e-15, 3.819441e-15, 3.830707e-15, 3.840498e-15, 3.849429e-15, 
    3.848775e-15, 3.849005e-15, 3.850998e-15, 3.846059e-15, 3.851809e-15, 
    3.852773e-15, 3.850251e-15, 3.864878e-15, 3.860702e-15, 3.864975e-15, 
    3.862257e-15, 3.793631e-15, 3.797045e-15, 3.795201e-15, 3.798669e-15, 
    3.796225e-15, 3.807085e-15, 3.810339e-15, 3.825552e-15, 3.819314e-15, 
    3.829243e-15, 3.820324e-15, 3.821905e-15, 3.829562e-15, 3.820807e-15, 
    3.839957e-15, 3.826974e-15, 3.851076e-15, 3.838124e-15, 3.851887e-15, 
    3.84939e-15, 3.853523e-15, 3.857222e-15, 3.861876e-15, 3.870452e-15, 
    3.868467e-15, 3.875637e-15, 3.802134e-15, 3.806558e-15, 3.80617e-15, 
    3.810798e-15, 3.814219e-15, 3.821632e-15, 3.833507e-15, 3.829044e-15, 
    3.837238e-15, 3.838881e-15, 3.826434e-15, 3.834076e-15, 3.809518e-15, 
    3.813488e-15, 3.811126e-15, 3.802482e-15, 3.83007e-15, 3.815921e-15, 
    3.842033e-15, 3.834381e-15, 3.856695e-15, 3.845603e-15, 3.867374e-15, 
    3.876659e-15, 3.885398e-15, 3.895588e-15, 3.808973e-15, 3.805968e-15, 
    3.811349e-15, 3.818786e-15, 3.825686e-15, 3.834848e-15, 3.835786e-15, 
    3.837501e-15, 3.841943e-15, 3.845675e-15, 3.838041e-15, 3.846611e-15, 
    3.814405e-15, 3.831298e-15, 3.80483e-15, 3.812805e-15, 3.818348e-15, 
    3.815919e-15, 3.828534e-15, 3.831504e-15, 3.843563e-15, 3.837332e-15, 
    3.874367e-15, 3.858001e-15, 3.903345e-15, 3.890697e-15, 3.804917e-15, 
    3.808963e-15, 3.823028e-15, 3.816339e-15, 3.83546e-15, 3.84016e-15, 
    3.84398e-15, 3.848858e-15, 3.849386e-15, 3.852275e-15, 3.84754e-15, 
    3.852089e-15, 3.834867e-15, 3.842568e-15, 3.821424e-15, 3.826573e-15, 
    3.824206e-15, 3.821606e-15, 3.829627e-15, 3.83816e-15, 3.838346e-15, 
    3.84108e-15, 3.848775e-15, 3.835538e-15, 3.876471e-15, 3.851209e-15, 
    3.813373e-15, 3.821153e-15, 3.822268e-15, 3.819254e-15, 3.839688e-15, 
    3.83229e-15, 3.852205e-15, 3.846828e-15, 3.855638e-15, 3.851261e-15, 
    3.850616e-15, 3.844992e-15, 3.841488e-15, 3.832628e-15, 3.825415e-15, 
    3.819692e-15, 3.821023e-15, 3.827308e-15, 3.838683e-15, 3.849432e-15, 
    3.847078e-15, 3.854968e-15, 3.834075e-15, 3.84284e-15, 3.839453e-15, 
    3.848284e-15, 3.828925e-15, 3.845403e-15, 3.824707e-15, 3.826524e-15, 
    3.832143e-15, 3.843432e-15, 3.845933e-15, 3.848596e-15, 3.846953e-15, 
    3.838972e-15, 3.837665e-15, 3.832007e-15, 3.830442e-15, 3.826129e-15, 
    3.822554e-15, 3.82582e-15, 3.829246e-15, 3.838977e-15, 3.847735e-15, 
    3.857275e-15, 3.859609e-15, 3.870731e-15, 3.861674e-15, 3.876611e-15, 
    3.863907e-15, 3.88589e-15, 3.846362e-15, 3.86354e-15, 3.832399e-15, 
    3.83576e-15, 3.841832e-15, 3.85575e-15, 3.848243e-15, 3.857024e-15, 
    3.837614e-15, 3.827524e-15, 3.824915e-15, 3.820039e-15, 3.825026e-15, 
    3.824621e-15, 3.82939e-15, 3.827858e-15, 3.8393e-15, 3.833156e-15, 
    3.850599e-15, 3.856955e-15, 3.874884e-15, 3.885855e-15, 3.897012e-15, 
    3.901931e-15, 3.903429e-15, 3.904054e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.535308e-09, -8.572939e-09, -8.565624e-09, -8.595976e-09, -8.579139e-09, 
    -8.599014e-09, -8.542937e-09, -8.574432e-09, -8.554327e-09, 
    -8.538696e-09, -8.65488e-09, -8.597331e-09, -8.714673e-09, -8.677964e-09, 
    -8.770182e-09, -8.708959e-09, -8.782528e-09, -8.768418e-09, 
    -8.810892e-09, -8.798724e-09, -8.853048e-09, -8.816508e-09, 
    -8.881213e-09, -8.844323e-09, -8.850092e-09, -8.815302e-09, 
    -8.608914e-09, -8.647715e-09, -8.606614e-09, -8.612147e-09, 
    -8.609665e-09, -8.579486e-09, -8.564277e-09, -8.532433e-09, 
    -8.538214e-09, -8.561604e-09, -8.614635e-09, -8.596635e-09, 
    -8.642005e-09, -8.64098e-09, -8.691494e-09, -8.668718e-09, -8.753624e-09, 
    -8.729493e-09, -8.799232e-09, -8.781692e-09, -8.798407e-09, 
    -8.793339e-09, -8.798473e-09, -8.772751e-09, -8.783771e-09, 
    -8.761137e-09, -8.672983e-09, -8.698889e-09, -8.621626e-09, 
    -8.575169e-09, -8.544318e-09, -8.522425e-09, -8.525521e-09, -8.53142e-09, 
    -8.561742e-09, -8.590251e-09, -8.611979e-09, -8.626513e-09, 
    -8.640834e-09, -8.684178e-09, -8.707125e-09, -8.758503e-09, 
    -8.749232e-09, -8.76494e-09, -8.779947e-09, -8.805142e-09, -8.800995e-09, 
    -8.812096e-09, -8.764526e-09, -8.79614e-09, -8.743951e-09, -8.758225e-09, 
    -8.64472e-09, -8.601491e-09, -8.583112e-09, -8.56703e-09, -8.5279e-09, 
    -8.554921e-09, -8.544269e-09, -8.569613e-09, -8.585717e-09, 
    -8.577753e-09, -8.62691e-09, -8.607798e-09, -8.708485e-09, -8.665114e-09, 
    -8.778197e-09, -8.751136e-09, -8.784683e-09, -8.767565e-09, 
    -8.796896e-09, -8.770498e-09, -8.816228e-09, -8.826184e-09, -8.81938e-09, 
    -8.845521e-09, -8.769035e-09, -8.798406e-09, -8.577529e-09, 
    -8.578828e-09, -8.584879e-09, -8.558277e-09, -8.55665e-09, -8.532274e-09, 
    -8.553964e-09, -8.563201e-09, -8.586651e-09, -8.600521e-09, 
    -8.613706e-09, -8.642698e-09, -8.675077e-09, -8.720356e-09, -8.75289e-09, 
    -8.774697e-09, -8.761326e-09, -8.773132e-09, -8.759934e-09, 
    -8.753749e-09, -8.822453e-09, -8.783873e-09, -8.841761e-09, 
    -8.838558e-09, -8.81236e-09, -8.838919e-09, -8.57974e-09, -8.572266e-09, 
    -8.546312e-09, -8.566623e-09, -8.529619e-09, -8.550331e-09, -8.56224e-09, 
    -8.608196e-09, -8.618295e-09, -8.627658e-09, -8.64615e-09, -8.669883e-09, 
    -8.711518e-09, -8.747747e-09, -8.780821e-09, -8.778398e-09, -8.77925e-09, 
    -8.786638e-09, -8.768337e-09, -8.789643e-09, -8.793219e-09, -8.78387e-09, 
    -8.838128e-09, -8.822627e-09, -8.83849e-09, -8.828397e-09, -8.574696e-09, 
    -8.587273e-09, -8.580477e-09, -8.593257e-09, -8.584252e-09, -8.62429e-09, 
    -8.636294e-09, -8.692469e-09, -8.669416e-09, -8.706108e-09, 
    -8.673144e-09, -8.678984e-09, -8.707302e-09, -8.674926e-09, 
    -8.745747e-09, -8.69773e-09, -8.786926e-09, -8.73897e-09, -8.789931e-09, 
    -8.780678e-09, -8.795999e-09, -8.80972e-09, -8.826984e-09, -8.858836e-09, 
    -8.851461e-09, -8.878101e-09, -8.606024e-09, -8.622338e-09, 
    -8.620903e-09, -8.637977e-09, -8.650604e-09, -8.677975e-09, 
    -8.721874e-09, -8.705366e-09, -8.735674e-09, -8.741758e-09, 
    -8.695713e-09, -8.723982e-09, -8.633258e-09, -8.647913e-09, 
    -8.639188e-09, -8.607311e-09, -8.709168e-09, -8.656892e-09, 
    -8.753427e-09, -8.725106e-09, -8.807763e-09, -8.766654e-09, -8.8474e-09, 
    -8.881917e-09, -8.914411e-09, -8.952378e-09, -8.631243e-09, 
    -8.620158e-09, -8.640008e-09, -8.667469e-09, -8.692954e-09, 
    -8.726833e-09, -8.7303e-09, -8.736647e-09, -8.753089e-09, -8.766913e-09, 
    -8.738653e-09, -8.770378e-09, -8.651311e-09, -8.713706e-09, 
    -8.615967e-09, -8.645395e-09, -8.665851e-09, -8.656879e-09, -8.70348e-09, 
    -8.714463e-09, -8.759096e-09, -8.736023e-09, -8.873397e-09, 
    -8.812616e-09, -8.981292e-09, -8.93415e-09, -8.616285e-09, -8.631206e-09, 
    -8.683136e-09, -8.658428e-09, -8.729096e-09, -8.746491e-09, 
    -8.760633e-09, -8.778709e-09, -8.780662e-09, -8.791373e-09, 
    -8.773822e-09, -8.79068e-09, -8.726905e-09, -8.755404e-09, -8.677202e-09, 
    -8.696235e-09, -8.687479e-09, -8.677874e-09, -8.707517e-09, 
    -8.739097e-09, -8.739774e-09, -8.7499e-09, -8.778432e-09, -8.729383e-09, 
    -8.881239e-09, -8.78745e-09, -8.647477e-09, -8.676215e-09, -8.680323e-09, 
    -8.66919e-09, -8.744746e-09, -8.717369e-09, -8.791112e-09, -8.771182e-09, 
    -8.803838e-09, -8.787611e-09, -8.785222e-09, -8.764381e-09, 
    -8.751405e-09, -8.718624e-09, -8.691952e-09, -8.670805e-09, 
    -8.675722e-09, -8.698953e-09, -8.74103e-09, -8.780838e-09, -8.772117e-09, 
    -8.801356e-09, -8.723972e-09, -8.756419e-09, -8.743877e-09, 
    -8.776579e-09, -8.704927e-09, -8.765936e-09, -8.689332e-09, 
    -8.696049e-09, -8.716825e-09, -8.758618e-09, -8.767867e-09, -8.77774e-09, 
    -8.771648e-09, -8.742099e-09, -8.737258e-09, -8.716321e-09, 
    -8.710539e-09, -8.694586e-09, -8.681379e-09, -8.693446e-09, 
    -8.706118e-09, -8.742111e-09, -8.774548e-09, -8.809915e-09, 
    -8.818571e-09, -8.859891e-09, -8.826252e-09, -8.881761e-09, 
    -8.834564e-09, -8.916268e-09, -8.769476e-09, -8.83318e-09, -8.717771e-09, 
    -8.730204e-09, -8.75269e-09, -8.80427e-09, -8.776426e-09, -8.808991e-09, 
    -8.737068e-09, -8.699754e-09, -8.690101e-09, -8.67209e-09, -8.690513e-09, 
    -8.689015e-09, -8.706644e-09, -8.700979e-09, -8.743307e-09, -8.72057e-09, 
    -8.785162e-09, -8.808734e-09, -8.875308e-09, -8.916121e-09, 
    -8.957672e-09, -8.976015e-09, -8.981599e-09, -8.983933e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.012876e-10, -1.017343e-10, -1.016474e-10, -1.020078e-10, -1.018079e-10, 
    -1.020438e-10, -1.013781e-10, -1.01752e-10, -1.015133e-10, -1.013278e-10, 
    -1.02707e-10, -1.020238e-10, -1.034169e-10, -1.029811e-10, -1.040759e-10, 
    -1.033491e-10, -1.042225e-10, -1.040549e-10, -1.045592e-10, 
    -1.044147e-10, -1.050597e-10, -1.046259e-10, -1.053941e-10, 
    -1.049561e-10, -1.050246e-10, -1.046115e-10, -1.021614e-10, -1.02622e-10, 
    -1.021341e-10, -1.021997e-10, -1.021703e-10, -1.01812e-10, -1.016315e-10, 
    -1.012534e-10, -1.013221e-10, -1.015997e-10, -1.022293e-10, 
    -1.020156e-10, -1.025542e-10, -1.02542e-10, -1.031417e-10, -1.028713e-10, 
    -1.038793e-10, -1.035928e-10, -1.044207e-10, -1.042125e-10, -1.04411e-10, 
    -1.043508e-10, -1.044118e-10, -1.041064e-10, -1.042372e-10, 
    -1.039685e-10, -1.02922e-10, -1.032295e-10, -1.023123e-10, -1.017608e-10, 
    -1.013945e-10, -1.011346e-10, -1.011714e-10, -1.012414e-10, 
    -1.016014e-10, -1.019398e-10, -1.021977e-10, -1.023703e-10, 
    -1.025403e-10, -1.030549e-10, -1.033273e-10, -1.039372e-10, 
    -1.038272e-10, -1.040136e-10, -1.041918e-10, -1.044909e-10, 
    -1.044417e-10, -1.045735e-10, -1.040087e-10, -1.043841e-10, 
    -1.037645e-10, -1.039339e-10, -1.025864e-10, -1.020732e-10, 
    -1.018551e-10, -1.016641e-10, -1.011996e-10, -1.015204e-10, 
    -1.013939e-10, -1.016948e-10, -1.01886e-10, -1.017914e-10, -1.02375e-10, 
    -1.021481e-10, -1.033434e-10, -1.028285e-10, -1.04171e-10, -1.038498e-10, 
    -1.04248e-10, -1.040448e-10, -1.04393e-10, -1.040796e-10, -1.046225e-10, 
    -1.047407e-10, -1.0466e-10, -1.049703e-10, -1.040623e-10, -1.04411e-10, 
    -1.017888e-10, -1.018042e-10, -1.01876e-10, -1.015602e-10, -1.015409e-10, 
    -1.012515e-10, -1.01509e-10, -1.016187e-10, -1.018971e-10, -1.020617e-10, 
    -1.022182e-10, -1.025624e-10, -1.029468e-10, -1.034844e-10, 
    -1.038706e-10, -1.041295e-10, -1.039707e-10, -1.041109e-10, 
    -1.039542e-10, -1.038808e-10, -1.046964e-10, -1.042384e-10, 
    -1.049257e-10, -1.048876e-10, -1.045766e-10, -1.048919e-10, -1.01815e-10, 
    -1.017263e-10, -1.014182e-10, -1.016593e-10, -1.0122e-10, -1.014659e-10, 
    -1.016073e-10, -1.021528e-10, -1.022727e-10, -1.023839e-10, 
    -1.026034e-10, -1.028852e-10, -1.033794e-10, -1.038095e-10, 
    -1.042022e-10, -1.041734e-10, -1.041835e-10, -1.042712e-10, -1.04054e-10, 
    -1.043069e-10, -1.043494e-10, -1.042384e-10, -1.048825e-10, 
    -1.046985e-10, -1.048868e-10, -1.04767e-10, -1.017551e-10, -1.019045e-10, 
    -1.018238e-10, -1.019755e-10, -1.018686e-10, -1.023439e-10, 
    -1.024864e-10, -1.031533e-10, -1.028796e-10, -1.033152e-10, 
    -1.029239e-10, -1.029932e-10, -1.033294e-10, -1.02945e-10, -1.037858e-10, 
    -1.032157e-10, -1.042747e-10, -1.037053e-10, -1.043103e-10, 
    -1.042005e-10, -1.043824e-10, -1.045453e-10, -1.047502e-10, 
    -1.051284e-10, -1.050408e-10, -1.053571e-10, -1.021271e-10, 
    -1.023207e-10, -1.023037e-10, -1.025064e-10, -1.026563e-10, 
    -1.029812e-10, -1.035024e-10, -1.033064e-10, -1.036662e-10, 
    -1.037384e-10, -1.031918e-10, -1.035274e-10, -1.024504e-10, 
    -1.026243e-10, -1.025208e-10, -1.021423e-10, -1.033515e-10, 
    -1.027309e-10, -1.03877e-10, -1.035407e-10, -1.04522e-10, -1.04034e-10, 
    -1.049926e-10, -1.054024e-10, -1.057882e-10, -1.06239e-10, -1.024264e-10, 
    -1.022948e-10, -1.025305e-10, -1.028565e-10, -1.03159e-10, -1.035612e-10, 
    -1.036024e-10, -1.036778e-10, -1.038729e-10, -1.040371e-10, 
    -1.037016e-10, -1.040782e-10, -1.026647e-10, -1.034054e-10, 
    -1.022451e-10, -1.025944e-10, -1.028373e-10, -1.027308e-10, -1.03284e-10, 
    -1.034144e-10, -1.039443e-10, -1.036704e-10, -1.053013e-10, 
    -1.045797e-10, -1.065822e-10, -1.060226e-10, -1.022489e-10, -1.02426e-10, 
    -1.030425e-10, -1.027492e-10, -1.035881e-10, -1.037946e-10, 
    -1.039625e-10, -1.041771e-10, -1.042003e-10, -1.043275e-10, 
    -1.041191e-10, -1.043192e-10, -1.035621e-10, -1.039004e-10, -1.02972e-10, 
    -1.03198e-10, -1.03094e-10, -1.0298e-10, -1.033319e-10, -1.037068e-10, 
    -1.037149e-10, -1.038351e-10, -1.041738e-10, -1.035915e-10, 
    -1.053944e-10, -1.042809e-10, -1.026191e-10, -1.029603e-10, 
    -1.030091e-10, -1.028769e-10, -1.037739e-10, -1.034489e-10, 
    -1.043244e-10, -1.040877e-10, -1.044754e-10, -1.042828e-10, 
    -1.042544e-10, -1.04007e-10, -1.03853e-10, -1.034638e-10, -1.031472e-10, 
    -1.028961e-10, -1.029545e-10, -1.032303e-10, -1.037298e-10, 
    -1.042024e-10, -1.040989e-10, -1.04446e-10, -1.035273e-10, -1.039125e-10, 
    -1.037636e-10, -1.041518e-10, -1.033012e-10, -1.040255e-10, -1.03116e-10, 
    -1.031958e-10, -1.034424e-10, -1.039386e-10, -1.040484e-10, 
    -1.041656e-10, -1.040933e-10, -1.037425e-10, -1.03685e-10, -1.034364e-10, 
    -1.033678e-10, -1.031784e-10, -1.030216e-10, -1.031649e-10, 
    -1.033153e-10, -1.037426e-10, -1.041277e-10, -1.045476e-10, 
    -1.046504e-10, -1.051409e-10, -1.047415e-10, -1.054006e-10, 
    -1.048402e-10, -1.058102e-10, -1.040675e-10, -1.048238e-10, 
    -1.034537e-10, -1.036013e-10, -1.038682e-10, -1.044806e-10, -1.0415e-10, 
    -1.045366e-10, -1.036828e-10, -1.032398e-10, -1.031252e-10, 
    -1.029114e-10, -1.031301e-10, -1.031123e-10, -1.033216e-10, 
    -1.032543e-10, -1.037568e-10, -1.034869e-10, -1.042537e-10, 
    -1.045336e-10, -1.053239e-10, -1.058085e-10, -1.063018e-10, 
    -1.065196e-10, -1.065859e-10, -1.066136e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.400407e-12, -8.437474e-12, -8.430269e-12, -8.460165e-12, -8.443581e-12, 
    -8.463157e-12, -8.407923e-12, -8.438944e-12, -8.419141e-12, 
    -8.403745e-12, -8.518184e-12, -8.461499e-12, -8.57708e-12, -8.540922e-12, 
    -8.631758e-12, -8.571453e-12, -8.643918e-12, -8.630019e-12, 
    -8.671857e-12, -8.659871e-12, -8.713382e-12, -8.677389e-12, 
    -8.741124e-12, -8.704787e-12, -8.71047e-12, -8.676201e-12, -8.472908e-12, 
    -8.511127e-12, -8.470643e-12, -8.476093e-12, -8.473648e-12, 
    -8.443923e-12, -8.428942e-12, -8.397575e-12, -8.40327e-12, -8.426309e-12, 
    -8.478544e-12, -8.460814e-12, -8.505503e-12, -8.504494e-12, 
    -8.554248e-12, -8.531815e-12, -8.615448e-12, -8.591678e-12, 
    -8.660371e-12, -8.643095e-12, -8.659559e-12, -8.654567e-12, 
    -8.659624e-12, -8.634287e-12, -8.645142e-12, -8.622847e-12, 
    -8.536016e-12, -8.561533e-12, -8.485429e-12, -8.43967e-12, -8.409283e-12, 
    -8.387718e-12, -8.390767e-12, -8.396579e-12, -8.426444e-12, 
    -8.454526e-12, -8.475927e-12, -8.490243e-12, -8.504349e-12, 
    -8.547043e-12, -8.569646e-12, -8.620254e-12, -8.611122e-12, 
    -8.626593e-12, -8.641376e-12, -8.666194e-12, -8.662109e-12, 
    -8.673042e-12, -8.626187e-12, -8.657326e-12, -8.60592e-12, -8.61998e-12, 
    -8.508178e-12, -8.465597e-12, -8.447494e-12, -8.431653e-12, 
    -8.393111e-12, -8.419727e-12, -8.409234e-12, -8.434198e-12, -8.45006e-12, 
    -8.442215e-12, -8.490634e-12, -8.471809e-12, -8.570985e-12, 
    -8.528266e-12, -8.639651e-12, -8.612997e-12, -8.646041e-12, 
    -8.629179e-12, -8.658071e-12, -8.632069e-12, -8.677112e-12, -8.68692e-12, 
    -8.680218e-12, -8.705967e-12, -8.630627e-12, -8.659558e-12, 
    -8.441994e-12, -8.443274e-12, -8.449235e-12, -8.423032e-12, 
    -8.421429e-12, -8.397419e-12, -8.418784e-12, -8.427882e-12, 
    -8.450979e-12, -8.464641e-12, -8.477629e-12, -8.506185e-12, 
    -8.538078e-12, -8.582679e-12, -8.614724e-12, -8.636205e-12, 
    -8.623034e-12, -8.634662e-12, -8.621662e-12, -8.61557e-12, -8.683245e-12, 
    -8.645243e-12, -8.702263e-12, -8.699108e-12, -8.673303e-12, 
    -8.699464e-12, -8.444172e-12, -8.43681e-12, -8.411247e-12, -8.431252e-12, 
    -8.394804e-12, -8.415205e-12, -8.426935e-12, -8.472201e-12, 
    -8.482149e-12, -8.491371e-12, -8.509586e-12, -8.532963e-12, 
    -8.573973e-12, -8.609657e-12, -8.642236e-12, -8.639849e-12, -8.64069e-12, 
    -8.647967e-12, -8.62994e-12, -8.650926e-12, -8.654449e-12, -8.64524e-12, 
    -8.698686e-12, -8.683416e-12, -8.699041e-12, -8.689099e-12, 
    -8.439203e-12, -8.451593e-12, -8.444898e-12, -8.457486e-12, 
    -8.448617e-12, -8.488053e-12, -8.499878e-12, -8.55521e-12, -8.532503e-12, 
    -8.568644e-12, -8.536174e-12, -8.541927e-12, -8.56982e-12, -8.537929e-12, 
    -8.607689e-12, -8.560391e-12, -8.64825e-12, -8.601013e-12, -8.65121e-12, 
    -8.642096e-12, -8.657187e-12, -8.670702e-12, -8.687708e-12, 
    -8.719083e-12, -8.711818e-12, -8.738059e-12, -8.470062e-12, 
    -8.486131e-12, -8.484718e-12, -8.501535e-12, -8.513973e-12, 
    -8.540933e-12, -8.584173e-12, -8.567913e-12, -8.597766e-12, 
    -8.603758e-12, -8.558406e-12, -8.586251e-12, -8.496887e-12, 
    -8.511323e-12, -8.502728e-12, -8.47133e-12, -8.571658e-12, -8.520167e-12, 
    -8.615253e-12, -8.587357e-12, -8.668775e-12, -8.628282e-12, 
    -8.707818e-12, -8.741818e-12, -8.773825e-12, -8.811223e-12, 
    -8.494903e-12, -8.483984e-12, -8.503536e-12, -8.530585e-12, 
    -8.555687e-12, -8.589058e-12, -8.592474e-12, -8.598725e-12, -8.61492e-12, 
    -8.628536e-12, -8.600701e-12, -8.63195e-12, -8.514669e-12, -8.576129e-12, 
    -8.479855e-12, -8.508842e-12, -8.528991e-12, -8.520153e-12, 
    -8.566055e-12, -8.576874e-12, -8.620837e-12, -8.598111e-12, 
    -8.733425e-12, -8.673556e-12, -8.839705e-12, -8.793269e-12, 
    -8.480169e-12, -8.494865e-12, -8.546017e-12, -8.521679e-12, 
    -8.591287e-12, -8.608421e-12, -8.622351e-12, -8.640157e-12, -8.64208e-12, 
    -8.652631e-12, -8.635342e-12, -8.651948e-12, -8.589129e-12, 
    -8.617202e-12, -8.540171e-12, -8.558918e-12, -8.550294e-12, 
    -8.540834e-12, -8.570033e-12, -8.601139e-12, -8.601805e-12, -8.61178e-12, 
    -8.639884e-12, -8.591569e-12, -8.741149e-12, -8.648766e-12, 
    -8.510893e-12, -8.5392e-12, -8.543246e-12, -8.532279e-12, -8.606703e-12, 
    -8.579736e-12, -8.652373e-12, -8.632742e-12, -8.664908e-12, 
    -8.648924e-12, -8.646572e-12, -8.626043e-12, -8.613262e-12, 
    -8.580972e-12, -8.5547e-12, -8.53387e-12, -8.538714e-12, -8.561596e-12, 
    -8.603042e-12, -8.642254e-12, -8.633664e-12, -8.662464e-12, 
    -8.586239e-12, -8.6182e-12, -8.605847e-12, -8.638058e-12, -8.567481e-12, 
    -8.627575e-12, -8.55212e-12, -8.558735e-12, -8.579201e-12, -8.620367e-12, 
    -8.629477e-12, -8.639201e-12, -8.633202e-12, -8.604095e-12, 
    -8.599327e-12, -8.578704e-12, -8.573009e-12, -8.557295e-12, 
    -8.544286e-12, -8.556171e-12, -8.568654e-12, -8.604107e-12, 
    -8.636058e-12, -8.670894e-12, -8.679421e-12, -8.720121e-12, 
    -8.686987e-12, -8.741664e-12, -8.695174e-12, -8.775655e-12, 
    -8.631061e-12, -8.69381e-12, -8.580132e-12, -8.592379e-12, -8.614527e-12, 
    -8.665334e-12, -8.637907e-12, -8.669984e-12, -8.59914e-12, -8.562385e-12, 
    -8.552877e-12, -8.535136e-12, -8.553283e-12, -8.551808e-12, 
    -8.569172e-12, -8.563592e-12, -8.605285e-12, -8.582889e-12, 
    -8.646512e-12, -8.669732e-12, -8.735308e-12, -8.77551e-12, -8.816438e-12, 
    -8.834507e-12, -8.840007e-12, -8.842306e-12 ;

 SMIN_NH4 =
  0.0004353462, 0.00043718, 0.0004368234, 0.0004383026, 0.000437482, 
    0.0004384504, 0.0004357177, 0.0004372525, 0.0004362726, 0.0004355108, 
    0.0004411724, 0.0004383681, 0.0004440855, 0.0004422969, 0.0004467897, 
    0.000443807, 0.0004473911, 0.0004467036, 0.0004487727, 0.0004481798, 
    0.000450826, 0.0004490461, 0.0004521978, 0.0004504009, 0.0004506819, 
    0.0004489871, 0.0004389329, 0.0004408236, 0.0004388208, 0.0004390904, 
    0.0004389693, 0.0004374987, 0.0004367575, 0.0004352055, 0.0004354872, 
    0.0004366271, 0.0004392112, 0.000438334, 0.0004405447, 0.0004404948, 
    0.0004429559, 0.0004418462, 0.0004459828, 0.0004448071, 0.0004482045, 
    0.00044735, 0.0004481643, 0.0004479173, 0.0004481673, 0.0004469142, 
    0.000447451, 0.0004463484, 0.0004420547, 0.0004433168, 0.0004395522, 
    0.0004372883, 0.0004357848, 0.0004347179, 0.0004348686, 0.0004351561, 
    0.0004366337, 0.0004380229, 0.0004390816, 0.0004397898, 0.0004404875, 
    0.0004425995, 0.0004437174, 0.0004462204, 0.0004457688, 0.0004465339, 
    0.000447265, 0.0004484922, 0.0004482902, 0.0004488309, 0.0004465134, 
    0.0004480535, 0.000445511, 0.0004462064, 0.0004406775, 0.0004385709, 
    0.0004376753, 0.0004368915, 0.0004349845, 0.0004363014, 0.0004357822, 
    0.0004370172, 0.0004378019, 0.0004374137, 0.0004398091, 0.0004388777, 
    0.0004437836, 0.0004416704, 0.0004471797, 0.0004458613, 0.0004474956, 
    0.0004466617, 0.0004480904, 0.0004468044, 0.000449032, 0.000449517, 
    0.0004491855, 0.0004504588, 0.0004467328, 0.0004481637, 0.0004374031, 
    0.0004374664, 0.0004377613, 0.0004364648, 0.0004363855, 0.0004351975, 
    0.0004362545, 0.0004367046, 0.0004378473, 0.000438523, 0.0004391655, 
    0.0004405782, 0.0004421557, 0.0004443618, 0.0004459467, 0.000447009, 
    0.0004463576, 0.0004469326, 0.0004462897, 0.0004459883, 0.0004493351, 
    0.0004474558, 0.0004502755, 0.0004501195, 0.0004488433, 0.000450137, 
    0.0004375108, 0.0004371464, 0.0004358817, 0.0004368714, 0.000435068, 
    0.0004360774, 0.0004366577, 0.000438897, 0.0004393891, 0.0004398453, 
    0.0004407463, 0.0004419026, 0.0004439311, 0.000445696, 0.0004473073, 
    0.0004471891, 0.0004472307, 0.0004475905, 0.0004466989, 0.0004477368, 
    0.0004479109, 0.0004474554, 0.0004500985, 0.0004493434, 0.000450116, 
    0.0004496243, 0.0004372648, 0.0004378776, 0.0004375463, 0.0004381691, 
    0.0004377303, 0.0004396812, 0.0004402661, 0.0004430031, 0.0004418798, 
    0.0004436676, 0.0004420613, 0.0004423459, 0.0004437256, 0.000442148, 
    0.0004455985, 0.000443259, 0.0004476044, 0.0004452681, 0.0004477507, 
    0.0004472999, 0.0004480461, 0.0004487146, 0.0004495554, 0.000451107, 
    0.0004507476, 0.0004520452, 0.0004387913, 0.0004395862, 0.0004395162, 
    0.0004403481, 0.0004409633, 0.0004422969, 0.0004444357, 0.0004436313, 
    0.0004451078, 0.0004454042, 0.0004431609, 0.0004445381, 0.0004401177, 
    0.0004408317, 0.0004404065, 0.0004388531, 0.0004438161, 0.000441269, 
    0.0004459723, 0.0004445924, 0.0004486191, 0.0004466165, 0.0004505498, 
    0.0004522311, 0.0004538137, 0.0004556628, 0.00044002, 0.0004394798, 
    0.0004404469, 0.000441785, 0.0004430266, 0.0004446772, 0.0004448461, 
    0.0004451552, 0.0004459561, 0.0004466296, 0.0004452528, 0.0004467983, 
    0.0004409972, 0.0004440372, 0.0004392748, 0.0004407088, 0.0004417054, 
    0.0004412682, 0.0004435387, 0.0004440737, 0.0004462481, 0.0004451241, 
    0.000451816, 0.0004488553, 0.0004570708, 0.0004547749, 0.000439291, 
    0.000440018, 0.0004425482, 0.0004413443, 0.0004447873, 0.0004456348, 
    0.0004463236, 0.0004472042, 0.0004472992, 0.000447821, 0.0004469659, 
    0.0004477872, 0.0004446801, 0.0004460686, 0.0004422584, 0.0004431857, 
    0.0004427591, 0.000442291, 0.0004437352, 0.0004452738, 0.0004453067, 
    0.0004458, 0.00044719, 0.0004448002, 0.0004521977, 0.000447629, 
    0.0004408107, 0.0004422109, 0.000442411, 0.0004418685, 0.0004455496, 
    0.0004442158, 0.0004478083, 0.0004468373, 0.0004484281, 0.0004476376, 
    0.0004475212, 0.0004465058, 0.0004458736, 0.0004442765, 0.0004429769, 
    0.0004419466, 0.000442186, 0.0004433179, 0.0004453678, 0.0004473072, 
    0.0004468822, 0.0004483065, 0.0004445365, 0.0004461173, 0.0004455062, 
    0.0004470994, 0.0004436097, 0.0004465821, 0.0004428498, 0.000443177, 
    0.0004441892, 0.0004462253, 0.0004466758, 0.0004471567, 0.0004468598, 
    0.0004454202, 0.0004451844, 0.0004441642, 0.0004438825, 0.0004431053, 
    0.0004424616, 0.0004430496, 0.0004436669, 0.0004454204, 0.0004470006, 
    0.0004487234, 0.000449145, 0.0004511577, 0.0004495191, 0.0004522229, 
    0.0004499239, 0.0004539035, 0.0004467543, 0.0004498576, 0.0004442353, 
    0.0004448409, 0.0004459364, 0.000448449, 0.0004470925, 0.0004486789, 
    0.0004451751, 0.000443357, 0.0004428867, 0.0004420091, 0.0004429066, 
    0.0004428336, 0.0004436925, 0.0004434164, 0.0004454785, 0.0004443708, 
    0.0004475175, 0.0004486658, 0.0004519086, 0.0004538964, 0.00045592, 
    0.0004568133, 0.0004570851, 0.0004571987 ;

 SMIN_NH4_vr =
  0.002856641, 0.002861575, 0.002860609, 0.002864585, 0.002862377, 
    0.002864974, 0.002857627, 0.002861748, 0.002859114, 0.00285706, 
    0.00287226, 0.002864738, 0.002880068, 0.002875273, 0.002887296, 
    0.002879313, 0.0028889, 0.002887059, 0.002892588, 0.002891, 0.002898056, 
    0.00289331, 0.002901709, 0.002896918, 0.002897663, 0.002893138, 
    0.002866277, 0.002871347, 0.002865969, 0.002866693, 0.002866365, 
    0.002862409, 0.002860413, 0.002856236, 0.00285699, 0.002860056, 
    0.002866996, 0.002864637, 0.002870569, 0.002870436, 0.002877027, 
    0.002874054, 0.002885129, 0.002881978, 0.002891062, 0.002888774, 
    0.002890948, 0.002890284, 0.002890948, 0.002887599, 0.002889028, 
    0.002886081, 0.002874648, 0.002878025, 0.002867928, 0.002861838, 
    0.002857794, 0.002854924, 0.002855323, 0.002856097, 0.002860068, 
    0.002863799, 0.002866642, 0.002868538, 0.002870407, 0.002876067, 
    0.002879061, 0.002885756, 0.002884548, 0.002886589, 0.002888543, 
    0.002891818, 0.002891277, 0.002892716, 0.00288652, 0.002890636, 
    0.002883833, 0.002885693, 0.00287094, 0.002865287, 0.002862876, 
    0.002860766, 0.002855633, 0.002859176, 0.002857776, 0.002861093, 
    0.002863201, 0.002862154, 0.002868587, 0.002866081, 0.002879233, 
    0.002873572, 0.002888319, 0.002884789, 0.002889155, 0.002886927, 
    0.002890738, 0.002887303, 0.002893247, 0.002894542, 0.002893651, 
    0.00289705, 0.002887093, 0.002890917, 0.002862143, 0.002862313, 
    0.002863102, 0.002859611, 0.002859396, 0.002856196, 0.002859036, 
    0.002860247, 0.002863316, 0.002865126, 0.002866848, 0.00287064, 
    0.002874867, 0.002880773, 0.002885014, 0.002887851, 0.002886108, 
    0.002887641, 0.00288592, 0.00288511, 0.002894048, 0.002889029, 
    0.002896553, 0.002896137, 0.002892726, 0.002896175, 0.002862427, 
    0.002861443, 0.002858039, 0.002860697, 0.002855842, 0.002858558, 
    0.002860114, 0.002866128, 0.002867447, 0.002868671, 0.002871086, 
    0.002874183, 0.002879616, 0.002884336, 0.002888645, 0.002888324, 
    0.002888434, 0.002889391, 0.002887006, 0.002889776, 0.002890236, 
    0.002889021, 0.002896072, 0.002894058, 0.002896116, 0.002894799, 
    0.002861758, 0.0028634, 0.002862506, 0.00286418, 0.002862994, 
    0.002868233, 0.002869799, 0.002877134, 0.002874121, 0.002878912, 
    0.002874602, 0.002875365, 0.002879055, 0.002874827, 0.002884065, 
    0.002877795, 0.002889425, 0.002883168, 0.00288981, 0.002888601, 
    0.002890591, 0.002892376, 0.002894615, 0.002898754, 0.00289779, 
    0.00290125, 0.002865851, 0.00286798, 0.002867793, 0.00287002, 
    0.002871667, 0.002875244, 0.00288097, 0.002878811, 0.002882761, 
    0.002883554, 0.002877542, 0.00288123, 0.002869376, 0.002871287, 
    0.002870146, 0.002865971, 0.00287928, 0.002872448, 0.002885047, 
    0.00288135, 0.002892113, 0.002886761, 0.00289726, 0.002901741, 
    0.002905955, 0.002910867, 0.002869142, 0.002867688, 0.00287028, 
    0.002873868, 0.002877191, 0.002881612, 0.002882061, 0.002882883, 
    0.002885023, 0.002886825, 0.002883136, 0.002887267, 0.002871724, 
    0.002879872, 0.002867098, 0.002870945, 0.002873613, 0.002872442, 
    0.002878525, 0.002879953, 0.002885767, 0.002882762, 0.002900625, 
    0.002892728, 0.002914606, 0.002908501, 0.002867178, 0.002869125, 
    0.002875906, 0.00287268, 0.002881899, 0.002884167, 0.002886004, 
    0.002888358, 0.002888606, 0.002890001, 0.002887709, 0.002889905, 
    0.002881588, 0.002885304, 0.002875098, 0.002877578, 0.002876434, 
    0.002875175, 0.002879041, 0.002883159, 0.002883245, 0.002884559, 
    0.002888268, 0.002881879, 0.002901627, 0.002889432, 0.002871249, 
    0.002874997, 0.002875531, 0.002874078, 0.002883931, 0.002880361, 
    0.002889967, 0.002887368, 0.002891615, 0.002889503, 0.002889185, 
    0.002886472, 0.002884774, 0.0028805, 0.002877012, 0.002874252, 
    0.002874888, 0.002877921, 0.002883402, 0.00288859, 0.00288745, 
    0.002891253, 0.002881167, 0.002885396, 0.002883755, 0.002888017, 
    0.002878741, 0.002886691, 0.002876703, 0.002877575, 0.002880281, 
    0.002885729, 0.002886929, 0.002888215, 0.002887416, 0.002883565, 
    0.00288293, 0.002880195, 0.002879436, 0.002877356, 0.002875624, 
    0.0028772, 0.002878847, 0.002883543, 0.002887764, 0.002892363, 
    0.002893489, 0.002898849, 0.002894477, 0.002901679, 0.002895547, 
    0.002906152, 0.002887145, 0.002895435, 0.002880406, 0.002882023, 
    0.00288495, 0.002891662, 0.002888035, 0.002892273, 0.002882903, 
    0.002878029, 0.002876767, 0.002874415, 0.002876815, 0.00287662, 
    0.002878917, 0.002878173, 0.002883689, 0.002880726, 0.002889135, 
    0.002892203, 0.002900851, 0.00290614, 0.002911525, 0.002913895, 
    0.002914616, 0.002914914,
  0.001594047, 0.001600114, 0.001598935, 0.001603825, 0.001601113, 
    0.001604314, 0.001595278, 0.001600354, 0.001597114, 0.001594594, 
    0.001613302, 0.001604043, 0.001622913, 0.001617017, 0.00163182, 
    0.001621995, 0.0016338, 0.001631538, 0.001638346, 0.001636396, 
    0.001645092, 0.001639245, 0.001649598, 0.001643697, 0.00164462, 
    0.001639052, 0.001605909, 0.00161215, 0.001605538, 0.001606429, 
    0.00160603, 0.001601169, 0.001598717, 0.001593584, 0.001594516, 
    0.001598287, 0.001606829, 0.001603932, 0.001611235, 0.00161107, 
    0.001619191, 0.00161553, 0.001629166, 0.001625293, 0.001636478, 
    0.001633667, 0.001636345, 0.001635533, 0.001636356, 0.001632233, 
    0.001634, 0.001630371, 0.001616216, 0.001620379, 0.001607955, 
    0.001600472, 0.0015955, 0.001591969, 0.001592468, 0.00159342, 
    0.001598309, 0.001602904, 0.001606403, 0.001608742, 0.001611046, 
    0.001618013, 0.001621701, 0.001629948, 0.001628461, 0.00163098, 
    0.001633387, 0.001637424, 0.00163676, 0.001638538, 0.001630914, 
    0.001635982, 0.001627614, 0.001629904, 0.001611668, 0.001604714, 
    0.001601752, 0.001599161, 0.001592852, 0.00159721, 0.001595492, 
    0.001599578, 0.001602173, 0.00160089, 0.001608806, 0.001605729, 
    0.001621919, 0.00161495, 0.001633106, 0.001628766, 0.001634146, 
    0.001631402, 0.001636103, 0.001631872, 0.0016392, 0.001640794, 
    0.001639705, 0.00164389, 0.001631637, 0.001636345, 0.001600854, 
    0.001601063, 0.001602038, 0.00159775, 0.001597488, 0.001593558, 
    0.001597056, 0.001598544, 0.001602324, 0.001604557, 0.00160668, 
    0.001611346, 0.001616552, 0.001623826, 0.001629048, 0.001632545, 
    0.001630401, 0.001632294, 0.001630178, 0.001629186, 0.001640196, 
    0.001634016, 0.001643288, 0.001642775, 0.00163858, 0.001642833, 
    0.00160121, 0.001600006, 0.001595822, 0.001599096, 0.00159313, 
    0.00159647, 0.001598389, 0.001605793, 0.001607419, 0.001608926, 
    0.001611902, 0.001615718, 0.001622407, 0.001628222, 0.001633527, 
    0.001633139, 0.001633275, 0.001634459, 0.001631525, 0.001634941, 
    0.001635514, 0.001634016, 0.001642707, 0.001640225, 0.001642764, 
    0.001641149, 0.001600398, 0.001602424, 0.001601329, 0.001603387, 
    0.001601937, 0.001608383, 0.001610314, 0.001619347, 0.001615642, 
    0.001621538, 0.001616242, 0.00161718, 0.001621728, 0.001616528, 
    0.001627901, 0.001620191, 0.001634505, 0.001626812, 0.001634987, 
    0.001633504, 0.00163596, 0.001638158, 0.001640922, 0.001646019, 
    0.00164484, 0.001649101, 0.001605444, 0.001608069, 0.001607839, 
    0.001610587, 0.001612618, 0.001617019, 0.00162407, 0.00162142, 
    0.001626286, 0.001627262, 0.001619869, 0.001624408, 0.001609827, 
    0.001612184, 0.001610781, 0.00160565, 0.001622029, 0.001613628, 
    0.001629134, 0.001624589, 0.001637844, 0.001631255, 0.00164419, 
    0.001649709, 0.001654903, 0.001660963, 0.001609503, 0.001607719, 
    0.001610914, 0.001615329, 0.001619425, 0.001624866, 0.001625423, 
    0.001626442, 0.00162908, 0.001631297, 0.001626763, 0.001631853, 
    0.001612729, 0.001622758, 0.001607044, 0.001611779, 0.001615069, 
    0.001613627, 0.001621117, 0.001622881, 0.001630043, 0.001626342, 
    0.001648347, 0.00163862, 0.001665575, 0.001658054, 0.001607096, 
    0.001609497, 0.001617847, 0.001613876, 0.00162523, 0.001628021, 
    0.00163029, 0.001633188, 0.001633502, 0.001635218, 0.001632405, 
    0.001635107, 0.001624878, 0.001629451, 0.001616895, 0.001619952, 
    0.001618546, 0.001617003, 0.001621765, 0.001626834, 0.001626944, 
    0.001628568, 0.00163314, 0.001625276, 0.001649598, 0.001634586, 
    0.001612115, 0.001616734, 0.001617396, 0.001615607, 0.001627741, 
    0.001623347, 0.001635176, 0.001631982, 0.001637216, 0.001634615, 
    0.001634232, 0.001630891, 0.00162881, 0.001623548, 0.001619264, 
    0.001615866, 0.001616657, 0.001620389, 0.001627144, 0.001633529, 
    0.001632131, 0.001636818, 0.001624407, 0.001629613, 0.001627601, 
    0.001632847, 0.001621349, 0.001631137, 0.001618844, 0.001619923, 
    0.00162326, 0.001629965, 0.00163145, 0.001633033, 0.001632057, 
    0.001627316, 0.00162654, 0.001623179, 0.00162225, 0.001619688, 
    0.001617566, 0.001619505, 0.00162154, 0.001627318, 0.001632521, 
    0.001638189, 0.001639575, 0.001646186, 0.001640803, 0.001649681, 
    0.001642131, 0.001655197, 0.001631706, 0.001641912, 0.001623412, 
    0.001625408, 0.001629015, 0.001637283, 0.001632822, 0.00163804, 
    0.001626509, 0.001620517, 0.001618968, 0.001616073, 0.001619034, 
    0.001618793, 0.001621625, 0.001620715, 0.00162751, 0.001623861, 
    0.001634222, 0.001637999, 0.001648654, 0.001655175, 0.001661809, 
    0.001664735, 0.001665625, 0.001665997,
  0.001500661, 0.001507298, 0.001506009, 0.00151136, 0.001508392, 
    0.001511895, 0.001502007, 0.001507562, 0.001504016, 0.001501259, 
    0.001521736, 0.001511598, 0.001532258, 0.0015258, 0.001542016, 
    0.001531253, 0.001544185, 0.001541706, 0.001549166, 0.001547029, 
    0.001556563, 0.001550152, 0.001561502, 0.001555033, 0.001556045, 
    0.00154994, 0.00151364, 0.001520474, 0.001513235, 0.00151421, 
    0.001513772, 0.001508453, 0.001505771, 0.001500154, 0.001501174, 
    0.0015053, 0.001514648, 0.001511476, 0.00151947, 0.001519289, 
    0.001528181, 0.001524173, 0.001539107, 0.001534865, 0.001547119, 
    0.001544038, 0.001546974, 0.001546084, 0.001546985, 0.001542467, 
    0.001544403, 0.001540427, 0.001524923, 0.001529482, 0.00151588, 
    0.001507691, 0.001502251, 0.001498388, 0.001498934, 0.001499975, 
    0.001505324, 0.001510351, 0.00151418, 0.001516741, 0.001519263, 
    0.001526893, 0.001530931, 0.001539964, 0.001538335, 0.001541095, 
    0.001543732, 0.001548156, 0.001547428, 0.001549377, 0.001541023, 
    0.001546576, 0.001537407, 0.001539915, 0.001519946, 0.001512332, 
    0.001509092, 0.001506256, 0.001499354, 0.001504121, 0.001502242, 
    0.001506712, 0.001509552, 0.001508147, 0.001516811, 0.001513444, 
    0.00153117, 0.001523538, 0.001543424, 0.001538669, 0.001544564, 
    0.001541557, 0.001546708, 0.001542072, 0.001550102, 0.00155185, 
    0.001550656, 0.001555243, 0.001541815, 0.001546974, 0.001508108, 
    0.001508337, 0.001509404, 0.001504713, 0.001504426, 0.001500126, 
    0.001503952, 0.001505581, 0.001509716, 0.001512161, 0.001514485, 
    0.001519592, 0.001525292, 0.001533258, 0.001538978, 0.00154281, 
    0.00154046, 0.001542534, 0.001540216, 0.001539129, 0.001551195, 
    0.001544421, 0.001554583, 0.001554021, 0.001549423, 0.001554085, 
    0.001508498, 0.00150718, 0.001502602, 0.001506185, 0.001499657, 
    0.001503311, 0.001505412, 0.001513513, 0.001515293, 0.001516943, 
    0.0015202, 0.001524378, 0.001531704, 0.001538074, 0.001543885, 
    0.00154346, 0.001543609, 0.001544907, 0.001541692, 0.001545435, 
    0.001546063, 0.001544421, 0.001553946, 0.001551226, 0.00155401, 
    0.001552238, 0.001507608, 0.001509826, 0.001508628, 0.001510881, 
    0.001509293, 0.001516349, 0.001518463, 0.001528352, 0.001524296, 
    0.001530752, 0.001524952, 0.00152598, 0.001530961, 0.001525266, 
    0.001537722, 0.001529278, 0.001544958, 0.00153653, 0.001545485, 
    0.00154386, 0.001546551, 0.00154896, 0.00155199, 0.001557578, 
    0.001556285, 0.001560957, 0.001513131, 0.001516005, 0.001515753, 
    0.00151876, 0.001520984, 0.001525802, 0.001533525, 0.001530622, 
    0.001535952, 0.001537021, 0.001528924, 0.001533896, 0.001517929, 
    0.00152051, 0.001518973, 0.001513358, 0.00153129, 0.001522091, 
    0.001539072, 0.001534093, 0.001548616, 0.001541396, 0.001555573, 
    0.001561625, 0.00156732, 0.001573969, 0.001517574, 0.001515621, 
    0.001519118, 0.001523953, 0.001528438, 0.001534397, 0.001535007, 
    0.001536123, 0.001539013, 0.001541442, 0.001536475, 0.001542051, 
    0.001521107, 0.001532088, 0.001514883, 0.001520066, 0.001523668, 
    0.001522089, 0.00153029, 0.001532222, 0.001540068, 0.001536013, 
    0.001560131, 0.001549468, 0.001579029, 0.001570778, 0.001514939, 
    0.001517568, 0.00152671, 0.001522361, 0.001534795, 0.001537853, 
    0.001540339, 0.001543514, 0.001543857, 0.001545739, 0.001542656, 
    0.001545617, 0.00153441, 0.00153942, 0.001525666, 0.001529015, 
    0.001527475, 0.001525785, 0.001531, 0.001536553, 0.001536672, 
    0.001538452, 0.001543464, 0.001534845, 0.001561505, 0.001545048, 
    0.001520433, 0.001525492, 0.001526215, 0.001524256, 0.001537546, 
    0.001532733, 0.001545693, 0.001542192, 0.001547928, 0.001545078, 
    0.001544658, 0.001540997, 0.001538717, 0.001532953, 0.001528262, 
    0.00152454, 0.001525406, 0.001529493, 0.001536893, 0.001543888, 
    0.001542356, 0.001547492, 0.001533894, 0.001539598, 0.001537393, 
    0.00154314, 0.001530544, 0.001541269, 0.001527801, 0.001528983, 
    0.001532637, 0.001539984, 0.00154161, 0.001543344, 0.001542274, 
    0.001537081, 0.00153623, 0.001532549, 0.001531531, 0.001528725, 
    0.001526401, 0.001528525, 0.001530754, 0.001537083, 0.001542783, 
    0.001548994, 0.001550514, 0.001557763, 0.001551861, 0.001561597, 
    0.001553319, 0.001567645, 0.001541891, 0.001553077, 0.001532804, 
    0.00153499, 0.001538942, 0.001548003, 0.001543113, 0.001548832, 
    0.001536197, 0.001529634, 0.001527936, 0.001524766, 0.001528009, 
    0.001527745, 0.001530847, 0.00152985, 0.001537293, 0.001533296, 
    0.001544648, 0.001548787, 0.001560467, 0.00156762, 0.001574896, 
    0.001578106, 0.001579083, 0.001579492,
  0.00142892, 0.001435685, 0.00143437, 0.001439825, 0.001436799, 0.001440371, 
    0.001430292, 0.001435953, 0.001432339, 0.001429529, 0.00145041, 
    0.001440069, 0.001461149, 0.001454556, 0.001471115, 0.001460123, 
    0.001473331, 0.001470799, 0.001478422, 0.001476238, 0.001485987, 
    0.00147943, 0.001491039, 0.001484421, 0.001485456, 0.001479213, 
    0.00144215, 0.001449122, 0.001441737, 0.001442731, 0.001442285, 
    0.001436862, 0.001434128, 0.001428403, 0.001429443, 0.001433647, 
    0.001443178, 0.001439943, 0.001448096, 0.001447912, 0.001456986, 
    0.001452895, 0.001468143, 0.00146381, 0.001476329, 0.001473181, 
    0.001476181, 0.001475272, 0.001476193, 0.001471576, 0.001473554, 
    0.001469491, 0.001453661, 0.001458314, 0.001444434, 0.001436086, 
    0.00143054, 0.001426604, 0.00142716, 0.001428221, 0.001433672, 
    0.001438796, 0.001442701, 0.001445312, 0.001447885, 0.001455672, 
    0.001459793, 0.001469019, 0.001467354, 0.001470174, 0.001472868, 
    0.00147739, 0.001476646, 0.001478638, 0.0014701, 0.001475775, 
    0.001466406, 0.001468969, 0.001448584, 0.001440816, 0.001437513, 
    0.001434623, 0.001427588, 0.001432446, 0.001430531, 0.001435087, 
    0.001437981, 0.00143655, 0.001445384, 0.00144195, 0.001460038, 
    0.001452248, 0.001472554, 0.001467696, 0.001473718, 0.001470645, 
    0.00147591, 0.001471172, 0.00147938, 0.001481166, 0.001479945, 
    0.001484636, 0.001470909, 0.001476181, 0.00143651, 0.001436743, 
    0.001437831, 0.001433049, 0.001432757, 0.001428375, 0.001432274, 
    0.001433934, 0.001438149, 0.001440642, 0.001443011, 0.00144822, 
    0.001454037, 0.001462169, 0.001468011, 0.001471926, 0.001469525, 
    0.001471645, 0.001469275, 0.001468165, 0.001480497, 0.001473573, 
    0.001483961, 0.001483387, 0.001478686, 0.001483451, 0.001436907, 
    0.001435564, 0.001430898, 0.001434549, 0.001427897, 0.001431621, 
    0.001433762, 0.001442021, 0.001443836, 0.001445518, 0.001448841, 
    0.001453104, 0.001460582, 0.001467087, 0.001473025, 0.00147259, 
    0.001472743, 0.001474069, 0.001470784, 0.001474608, 0.00147525, 
    0.001473572, 0.00148331, 0.001480528, 0.001483374, 0.001481563, 0.001436, 
    0.001438261, 0.001437039, 0.001439336, 0.001437718, 0.001444913, 
    0.00144707, 0.001457161, 0.00145302, 0.001459611, 0.00145369, 
    0.001454739, 0.001459825, 0.00145401, 0.001466729, 0.001458106, 
    0.001474121, 0.001465512, 0.00147466, 0.001472999, 0.001475749, 
    0.001478212, 0.00148131, 0.001487025, 0.001485702, 0.001490481, 
    0.001441631, 0.001444562, 0.001444304, 0.001447372, 0.001449641, 
    0.001454558, 0.001462442, 0.001459477, 0.00146492, 0.001466012, 
    0.001457744, 0.001462821, 0.001446524, 0.001449158, 0.00144759, 
    0.001441862, 0.00146016, 0.001450771, 0.001468107, 0.001463022, 
    0.001477861, 0.001470482, 0.001484973, 0.001491166, 0.001496993, 
    0.001503802, 0.001446162, 0.001444171, 0.001447737, 0.001452671, 
    0.001457248, 0.001463332, 0.001463955, 0.001465095, 0.001468046, 
    0.001470528, 0.001465455, 0.00147115, 0.001449768, 0.001460975, 
    0.001443417, 0.001448705, 0.00145238, 0.001450768, 0.001459138, 
    0.001461111, 0.001469125, 0.001464983, 0.001489638, 0.001478732, 
    0.001508985, 0.001500533, 0.001443475, 0.001446156, 0.001455485, 
    0.001451046, 0.001463739, 0.001466862, 0.001469401, 0.001472646, 
    0.001472996, 0.001474919, 0.001471768, 0.001474794, 0.001463345, 
    0.001468462, 0.001454419, 0.001457837, 0.001456265, 0.00145454, 
    0.001459864, 0.001465535, 0.001465656, 0.001467474, 0.001472597, 
    0.00146379, 0.001491045, 0.001474215, 0.001449079, 0.001454242, 
    0.001454979, 0.00145298, 0.001466549, 0.001461633, 0.001474872, 
    0.001471295, 0.001477156, 0.001474243, 0.001473815, 0.001470074, 
    0.001467744, 0.001461858, 0.001457068, 0.00145327, 0.001454153, 
    0.001458326, 0.001465882, 0.001473028, 0.001471463, 0.001476711, 
    0.001462818, 0.001468644, 0.001466393, 0.001472263, 0.001459399, 
    0.001470354, 0.001456598, 0.001457804, 0.001461535, 0.001469039, 
    0.0014707, 0.001472472, 0.001471378, 0.001466073, 0.001465204, 
    0.001461445, 0.001460406, 0.001457541, 0.001455169, 0.001457336, 
    0.001459613, 0.001466076, 0.001471899, 0.001478247, 0.0014798, 
    0.001487215, 0.001481179, 0.001491138, 0.001482671, 0.001497327, 
    0.001470989, 0.001482422, 0.001461705, 0.001463938, 0.001467975, 
    0.001477234, 0.001472236, 0.001478081, 0.00146517, 0.00145847, 
    0.001456736, 0.001453501, 0.00145681, 0.001456541, 0.001459707, 
    0.001458689, 0.00146629, 0.001462208, 0.001473804, 0.001478035, 
    0.00148998, 0.0014973, 0.00150475, 0.001508039, 0.00150904, 0.001509458,
  0.001343027, 0.001349267, 0.001348053, 0.001353088, 0.001350295, 
    0.001353592, 0.001344292, 0.001349515, 0.00134618, 0.001343588, 
    0.001362868, 0.001353313, 0.001372802, 0.001366701, 0.001382034, 
    0.001371852, 0.001384088, 0.00138174, 0.001388809, 0.001386783, 
    0.001395833, 0.001389744, 0.001400527, 0.001394378, 0.00139534, 
    0.001389544, 0.001355235, 0.001361678, 0.001354853, 0.001355772, 
    0.001355359, 0.001350353, 0.001347831, 0.00134255, 0.001343508, 
    0.001347387, 0.001356185, 0.001353197, 0.001360728, 0.001360558, 
    0.001368948, 0.001365164, 0.001379278, 0.001375265, 0.001386868, 
    0.001383948, 0.001386731, 0.001385887, 0.001386742, 0.001382461, 
    0.001384295, 0.001380528, 0.001365873, 0.001370178, 0.001357345, 
    0.001349637, 0.001344521, 0.001340892, 0.001341405, 0.001342383, 
    0.00134741, 0.001352138, 0.001355743, 0.001358156, 0.001360533, 
    0.001367734, 0.001371547, 0.00138009, 0.001378548, 0.001381161, 
    0.001383658, 0.001387852, 0.001387162, 0.00138901, 0.001381092, 
    0.001386354, 0.001377669, 0.001380044, 0.001361181, 0.001354003, 
    0.001350955, 0.001348287, 0.001341799, 0.001346279, 0.001344513, 
    0.001348715, 0.001351386, 0.001350065, 0.001358222, 0.00135505, 
    0.001371773, 0.001364566, 0.001383367, 0.001378864, 0.001384446, 
    0.001381597, 0.001386479, 0.001382086, 0.001389698, 0.001391357, 
    0.001390223, 0.001394577, 0.001381842, 0.001386731, 0.001350028, 
    0.001350243, 0.001351247, 0.001346835, 0.001346565, 0.001342524, 
    0.00134612, 0.001347651, 0.001351541, 0.001353842, 0.00135603, 
    0.001360843, 0.001366221, 0.001373746, 0.001379156, 0.001382784, 
    0.001380559, 0.001382524, 0.001380328, 0.001379299, 0.001390735, 
    0.001384312, 0.001393951, 0.001393417, 0.001389054, 0.001393477, 
    0.001350394, 0.001349155, 0.001344851, 0.001348219, 0.001342084, 
    0.001345517, 0.001347492, 0.001355116, 0.001356792, 0.001358346, 
    0.001361416, 0.001365358, 0.001372277, 0.001378301, 0.001383803, 
    0.0013834, 0.001383542, 0.001384772, 0.001381726, 0.001385272, 
    0.001385867, 0.001384311, 0.001393346, 0.001390764, 0.001393406, 
    0.001391725, 0.001349557, 0.001351644, 0.001350516, 0.001352637, 
    0.001351143, 0.001357787, 0.00135978, 0.001369111, 0.00136528, 
    0.001371378, 0.001365899, 0.00136687, 0.001371577, 0.001366195, 
    0.001377969, 0.001369986, 0.00138482, 0.001376842, 0.00138532, 
    0.00138378, 0.00138633, 0.001388614, 0.001391489, 0.001396797, 
    0.001395567, 0.001400007, 0.001354755, 0.001357463, 0.001357224, 
    0.001360059, 0.001362156, 0.001366702, 0.001373998, 0.001371254, 
    0.001376293, 0.001377304, 0.001369649, 0.001374349, 0.001359276, 
    0.00136171, 0.00136026, 0.001354969, 0.001371886, 0.001363201, 
    0.001379246, 0.001374535, 0.001388289, 0.001381447, 0.001394891, 
    0.001400645, 0.001406063, 0.001412399, 0.001358941, 0.001357101, 
    0.001360396, 0.001364957, 0.001369191, 0.001374823, 0.001375399, 
    0.001376455, 0.001379189, 0.001381489, 0.001376789, 0.001382066, 
    0.001362275, 0.001372641, 0.001356405, 0.001361291, 0.001364688, 
    0.001363198, 0.00137094, 0.001372766, 0.001380189, 0.001376351, 
    0.001399225, 0.001389097, 0.001417227, 0.001409357, 0.001356458, 
    0.001358935, 0.00136756, 0.001363455, 0.001375199, 0.001378092, 
    0.001380444, 0.001383452, 0.001383777, 0.00138556, 0.001382639, 
    0.001385444, 0.001374835, 0.001379574, 0.001366573, 0.001369736, 
    0.001368281, 0.001366685, 0.001371611, 0.001376863, 0.001376975, 
    0.001378659, 0.001383408, 0.001375246, 0.001400533, 0.001384909, 
    0.001361636, 0.001366411, 0.001367092, 0.001365242, 0.001377802, 
    0.001373249, 0.001385516, 0.001382199, 0.001387635, 0.001384933, 
    0.001384536, 0.001381068, 0.001378909, 0.001373458, 0.001369025, 
    0.001365511, 0.001366328, 0.001370188, 0.001377184, 0.001383807, 
    0.001382356, 0.001387222, 0.001374347, 0.001379743, 0.001377657, 
    0.001383098, 0.001371181, 0.001381329, 0.001368589, 0.001369705, 
    0.001373159, 0.00138011, 0.001381648, 0.001383291, 0.001382277, 
    0.001377361, 0.001376556, 0.001373075, 0.001372114, 0.001369462, 
    0.001367267, 0.001369273, 0.001371379, 0.001377363, 0.00138276, 
    0.001388647, 0.001390088, 0.001396974, 0.001391369, 0.00140062, 
    0.001392755, 0.001406374, 0.001381917, 0.001392523, 0.001373316, 
    0.001375383, 0.001379124, 0.001387708, 0.001383072, 0.001388494, 
    0.001376525, 0.001370321, 0.001368717, 0.001365724, 0.001368785, 
    0.001368536, 0.001371466, 0.001370525, 0.001377562, 0.001373781, 
    0.001384526, 0.001388451, 0.001399542, 0.001406349, 0.001413282, 
    0.001416345, 0.001417278, 0.001417667,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.21443e-06, 1.224907e-06, 1.222866e-06, 1.231344e-06, 1.226637e-06, 
    1.232193e-06, 1.21655e-06, 1.225323e-06, 1.219718e-06, 1.21537e-06, 
    1.24788e-06, 1.231722e-06, 1.264784e-06, 1.254392e-06, 1.280581e-06, 
    1.263163e-06, 1.284108e-06, 1.280077e-06, 1.292231e-06, 1.288743e-06, 
    1.304352e-06, 1.293842e-06, 1.312482e-06, 1.301838e-06, 1.3035e-06, 
    1.293495e-06, 1.234966e-06, 1.245863e-06, 1.234322e-06, 1.235872e-06, 
    1.235176e-06, 1.226734e-06, 1.22249e-06, 1.21363e-06, 1.215236e-06, 
    1.221745e-06, 1.236569e-06, 1.231526e-06, 1.244255e-06, 1.243967e-06, 
    1.258216e-06, 1.251781e-06, 1.275858e-06, 1.26899e-06, 1.288888e-06, 
    1.283868e-06, 1.288651e-06, 1.2872e-06, 1.28867e-06, 1.281313e-06, 
    1.284462e-06, 1.277998e-06, 1.252986e-06, 1.260311e-06, 1.23853e-06, 
    1.225528e-06, 1.216933e-06, 1.210853e-06, 1.211711e-06, 1.213349e-06, 
    1.221783e-06, 1.229741e-06, 1.235823e-06, 1.239901e-06, 1.243925e-06, 
    1.256147e-06, 1.262642e-06, 1.277248e-06, 1.274606e-06, 1.279084e-06, 
    1.283369e-06, 1.290581e-06, 1.289393e-06, 1.292575e-06, 1.278965e-06, 
    1.288001e-06, 1.273101e-06, 1.277167e-06, 1.24502e-06, 1.232886e-06, 
    1.227746e-06, 1.223257e-06, 1.212371e-06, 1.219883e-06, 1.216919e-06, 
    1.223977e-06, 1.228473e-06, 1.226248e-06, 1.240012e-06, 1.234651e-06, 
    1.263028e-06, 1.250764e-06, 1.282869e-06, 1.275148e-06, 1.284723e-06, 
    1.279833e-06, 1.288218e-06, 1.28067e-06, 1.29376e-06, 1.29662e-06, 
    1.294665e-06, 1.302182e-06, 1.280251e-06, 1.28865e-06, 1.226187e-06, 
    1.226549e-06, 1.22824e-06, 1.220817e-06, 1.220364e-06, 1.213585e-06, 
    1.219616e-06, 1.222189e-06, 1.228734e-06, 1.232613e-06, 1.236307e-06, 
    1.244449e-06, 1.253575e-06, 1.266395e-06, 1.275647e-06, 1.281869e-06, 
    1.278052e-06, 1.281421e-06, 1.277655e-06, 1.275891e-06, 1.295547e-06, 
    1.284491e-06, 1.301099e-06, 1.300177e-06, 1.292649e-06, 1.30028e-06, 
    1.226804e-06, 1.224717e-06, 1.217487e-06, 1.223143e-06, 1.212848e-06, 
    1.218605e-06, 1.221921e-06, 1.234763e-06, 1.237594e-06, 1.240222e-06, 
    1.24542e-06, 1.252109e-06, 1.263887e-06, 1.274182e-06, 1.283618e-06, 
    1.282926e-06, 1.283169e-06, 1.285282e-06, 1.280052e-06, 1.286141e-06, 
    1.287164e-06, 1.284489e-06, 1.300053e-06, 1.295597e-06, 1.300157e-06, 
    1.297254e-06, 1.225395e-06, 1.228908e-06, 1.227009e-06, 1.230581e-06, 
    1.228063e-06, 1.239276e-06, 1.242648e-06, 1.258491e-06, 1.251977e-06, 
    1.262353e-06, 1.253029e-06, 1.254678e-06, 1.262691e-06, 1.253531e-06, 
    1.273612e-06, 1.259979e-06, 1.285364e-06, 1.271683e-06, 1.286223e-06, 
    1.283576e-06, 1.28796e-06, 1.291892e-06, 1.296848e-06, 1.306018e-06, 
    1.303891e-06, 1.31158e-06, 1.234155e-06, 1.238728e-06, 1.238326e-06, 
    1.243121e-06, 1.246674e-06, 1.254393e-06, 1.266826e-06, 1.262143e-06, 
    1.270746e-06, 1.272477e-06, 1.259409e-06, 1.267424e-06, 1.241793e-06, 
    1.245915e-06, 1.24346e-06, 1.234513e-06, 1.263219e-06, 1.248444e-06, 
    1.275799e-06, 1.267741e-06, 1.29133e-06, 1.27957e-06, 1.302721e-06, 
    1.312684e-06, 1.322097e-06, 1.33314e-06, 1.241229e-06, 1.238116e-06, 
    1.243692e-06, 1.251428e-06, 1.258628e-06, 1.268234e-06, 1.269219e-06, 
    1.271023e-06, 1.275703e-06, 1.279646e-06, 1.271593e-06, 1.280634e-06, 
    1.246872e-06, 1.264506e-06, 1.236938e-06, 1.245206e-06, 1.250969e-06, 
    1.24844e-06, 1.261606e-06, 1.26472e-06, 1.277414e-06, 1.270844e-06, 
    1.31022e-06, 1.292722e-06, 1.341582e-06, 1.327832e-06, 1.23703e-06, 
    1.241218e-06, 1.255851e-06, 1.248878e-06, 1.268876e-06, 1.273824e-06, 
    1.277854e-06, 1.283015e-06, 1.283572e-06, 1.286636e-06, 1.281617e-06, 
    1.286437e-06, 1.268253e-06, 1.276362e-06, 1.254173e-06, 1.259555e-06, 
    1.257077e-06, 1.254363e-06, 1.26275e-06, 1.271718e-06, 1.27191e-06, 
    1.274793e-06, 1.282933e-06, 1.268955e-06, 1.312486e-06, 1.285511e-06, 
    1.245793e-06, 1.253896e-06, 1.255056e-06, 1.251912e-06, 1.273327e-06, 
    1.265546e-06, 1.286561e-06, 1.280864e-06, 1.290206e-06, 1.285559e-06, 
    1.284876e-06, 1.278922e-06, 1.275222e-06, 1.265901e-06, 1.258342e-06, 
    1.252366e-06, 1.253754e-06, 1.260324e-06, 1.272267e-06, 1.283621e-06, 
    1.281129e-06, 1.289493e-06, 1.267418e-06, 1.27665e-06, 1.273077e-06, 
    1.282403e-06, 1.262018e-06, 1.279367e-06, 1.257603e-06, 1.259503e-06, 
    1.265391e-06, 1.277279e-06, 1.279917e-06, 1.282737e-06, 1.280996e-06, 
    1.272572e-06, 1.271195e-06, 1.265247e-06, 1.263607e-06, 1.259088e-06, 
    1.255352e-06, 1.258765e-06, 1.262353e-06, 1.272575e-06, 1.281823e-06, 
    1.291946e-06, 1.29443e-06, 1.306321e-06, 1.296636e-06, 1.312637e-06, 
    1.299025e-06, 1.322634e-06, 1.280377e-06, 1.29863e-06, 1.26566e-06, 
    1.26919e-06, 1.275589e-06, 1.290329e-06, 1.282361e-06, 1.291682e-06, 
    1.271141e-06, 1.260551e-06, 1.257819e-06, 1.252729e-06, 1.257935e-06, 
    1.257511e-06, 1.262502e-06, 1.260897e-06, 1.272915e-06, 1.266452e-06, 
    1.284856e-06, 1.291607e-06, 1.310771e-06, 1.322592e-06, 1.334682e-06, 
    1.340038e-06, 1.34167e-06, 1.342352e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  7.62962e-06, 7.663833e-06, 7.657164e-06, 7.684774e-06, 7.66945e-06, 
    7.687516e-06, 7.636518e-06, 7.66513e-06, 7.646854e-06, 7.632637e-06, 
    7.738333e-06, 7.685942e-06, 7.792898e-06, 7.759395e-06, 7.843597e-06, 
    7.787654e-06, 7.854883e-06, 7.841975e-06, 7.880833e-06, 7.869683e-06, 
    7.919392e-06, 7.885952e-06, 7.945202e-06, 7.911397e-06, 7.916667e-06, 
    7.884806e-06, 7.696551e-06, 7.731862e-06, 7.69444e-06, 7.699475e-06, 
    7.697209e-06, 7.669728e-06, 7.655881e-06, 7.626941e-06, 7.632183e-06, 
    7.653437e-06, 7.70168e-06, 7.685288e-06, 7.7266e-06, 7.725669e-06, 
    7.771707e-06, 7.750935e-06, 7.828442e-06, 7.806382e-06, 7.870139e-06, 
    7.854078e-06, 7.869366e-06, 7.864717e-06, 7.869403e-06, 7.845872e-06, 
    7.855933e-06, 7.83524e-06, 7.754918e-06, 7.778539e-06, 7.708093e-06, 
    7.665777e-06, 7.637736e-06, 7.617852e-06, 7.620644e-06, 7.626002e-06, 
    7.653545e-06, 7.679474e-06, 7.69925e-06, 7.712473e-06, 7.725511e-06, 
    7.765004e-06, 7.785947e-06, 7.832876e-06, 7.824408e-06, 7.838745e-06, 
    7.852473e-06, 7.875509e-06, 7.871713e-06, 7.881856e-06, 7.838332e-06, 
    7.867242e-06, 7.819513e-06, 7.832556e-06, 7.729092e-06, 7.689746e-06, 
    7.672996e-06, 7.65837e-06, 7.622798e-06, 7.647351e-06, 7.637659e-06, 
    7.660695e-06, 7.675338e-06, 7.668083e-06, 7.712826e-06, 7.695407e-06, 
    7.787176e-06, 7.747614e-06, 7.850882e-06, 7.826128e-06, 7.856793e-06, 
    7.84114e-06, 7.867944e-06, 7.843806e-06, 7.885624e-06, 7.894736e-06, 
    7.88849e-06, 7.912437e-06, 7.842415e-06, 7.869278e-06, 7.667925e-06, 
    7.669108e-06, 7.674605e-06, 7.650387e-06, 7.648907e-06, 7.626746e-06, 
    7.646447e-06, 7.654842e-06, 7.676169e-06, 7.688775e-06, 7.700769e-06, 
    7.72718e-06, 7.75668e-06, 7.797995e-06, 7.827722e-06, 7.84765e-06, 
    7.835421e-06, 7.846201e-06, 7.83413e-06, 7.828466e-06, 7.891294e-06, 
    7.855992e-06, 7.908968e-06, 7.906036e-06, 7.882031e-06, 7.906344e-06, 
    7.669922e-06, 7.663112e-06, 7.639507e-06, 7.657964e-06, 7.624319e-06, 
    7.643137e-06, 7.653946e-06, 7.695749e-06, 7.704944e-06, 7.71347e-06, 
    7.730312e-06, 7.751934e-06, 7.789917e-06, 7.822998e-06, 7.85324e-06, 
    7.851011e-06, 7.851788e-06, 7.85853e-06, 7.84179e-06, 7.861262e-06, 
    7.864518e-06, 7.855972e-06, 7.905619e-06, 7.891425e-06, 7.905941e-06, 
    7.896686e-06, 7.665313e-06, 7.676741e-06, 7.670547e-06, 7.682174e-06, 
    7.673962e-06, 7.710403e-06, 7.721325e-06, 7.772536e-06, 7.751506e-06, 
    7.784981e-06, 7.754892e-06, 7.760217e-06, 7.786025e-06, 7.756498e-06, 
    7.821137e-06, 7.777266e-06, 7.858783e-06, 7.814904e-06, 7.861517e-06, 
    7.853042e-06, 7.867047e-06, 7.879601e-06, 7.89539e-06, 7.924562e-06, 
    7.917789e-06, 7.942207e-06, 7.693799e-06, 7.708634e-06, 7.707333e-06, 
    7.722871e-06, 7.734366e-06, 7.759329e-06, 7.799381e-06, 7.784301e-06, 
    7.811968e-06, 7.817525e-06, 7.775465e-06, 7.801265e-06, 7.718498e-06, 
    7.731832e-06, 7.723888e-06, 7.694839e-06, 7.78769e-06, 7.739985e-06, 
    7.828112e-06, 7.802225e-06, 7.877786e-06, 7.840174e-06, 7.914063e-06, 
    7.945681e-06, 7.975496e-06, 8.010316e-06, 7.716741e-06, 7.706636e-06, 
    7.724708e-06, 7.749729e-06, 7.772967e-06, 7.8039e-06, 7.807061e-06, 
    7.812843e-06, 7.82786e-06, 7.840498e-06, 7.814647e-06, 7.843643e-06, 
    7.7349e-06, 7.791836e-06, 7.702704e-06, 7.729504e-06, 7.748142e-06, 
    7.739968e-06, 7.782474e-06, 7.792487e-06, 7.833243e-06, 7.81217e-06, 
    7.937842e-06, 7.882179e-06, 8.036875e-06, 7.99357e-06, 7.703098e-06, 
    7.716677e-06, 7.763999e-06, 7.741472e-06, 7.805947e-06, 7.821838e-06, 
    7.834751e-06, 7.851274e-06, 7.853047e-06, 7.862844e-06, 7.846776e-06, 
    7.862197e-06, 7.803877e-06, 7.829922e-06, 7.758506e-06, 7.775853e-06, 
    7.767866e-06, 7.759091e-06, 7.78613e-06, 7.814959e-06, 7.815579e-06, 
    7.824812e-06, 7.85085e-06, 7.806057e-06, 7.944974e-06, 7.859075e-06, 
    7.731493e-06, 7.757667e-06, 7.761417e-06, 7.751268e-06, 7.82022e-06, 
    7.795214e-06, 7.862606e-06, 7.844366e-06, 7.874229e-06, 7.859382e-06, 
    7.857178e-06, 7.838124e-06, 7.826242e-06, 7.796291e-06, 7.771928e-06, 
    7.752645e-06, 7.757111e-06, 7.778301e-06, 7.816702e-06, 7.853101e-06, 
    7.845111e-06, 7.871855e-06, 7.801097e-06, 7.830738e-06, 7.819257e-06, 
    7.849161e-06, 7.783862e-06, 7.839561e-06, 7.769627e-06, 7.775742e-06, 
    7.794693e-06, 7.832864e-06, 7.84132e-06, 7.850343e-06, 7.844761e-06, 
    7.817742e-06, 7.813313e-06, 7.794182e-06, 7.788886e-06, 7.774335e-06, 
    7.762265e-06, 7.773275e-06, 7.784816e-06, 7.817694e-06, 7.84733e-06, 
    7.879676e-06, 7.887601e-06, 7.925402e-06, 7.894592e-06, 7.945408e-06, 
    7.902154e-06, 7.977059e-06, 7.84279e-06, 7.901083e-06, 7.795563e-06, 
    7.806905e-06, 7.827432e-06, 7.874589e-06, 7.849121e-06, 7.878903e-06, 
    7.813136e-06, 7.779038e-06, 7.770233e-06, 7.753802e-06, 7.770593e-06, 
    7.769228e-06, 7.785307e-06, 7.780124e-06, 7.818763e-06, 7.797999e-06, 
    7.85701e-06, 7.878574e-06, 7.939547e-06, 7.976959e-06, 8.015115e-06, 
    8.031952e-06, 8.037081e-06, 8.039216e-06,
  3.976129e-06, 4.006499e-06, 4.00059e-06, 4.025133e-06, 4.011514e-06, 
    4.027592e-06, 3.982283e-06, 4.007704e-06, 3.99147e-06, 3.978864e-06, 
    4.072916e-06, 4.026229e-06, 4.121659e-06, 4.091719e-06, 4.167096e-06, 
    4.116991e-06, 4.177228e-06, 4.165655e-06, 4.200542e-06, 4.190537e-06, 
    4.235262e-06, 4.205163e-06, 4.258528e-06, 4.228071e-06, 4.232827e-06, 
    4.20417e-06, 4.035615e-06, 4.06709e-06, 4.033751e-06, 4.038234e-06, 
    4.036224e-06, 4.011792e-06, 3.999497e-06, 3.973817e-06, 3.978475e-06, 
    3.997342e-06, 4.04025e-06, 4.02567e-06, 4.062469e-06, 4.061636e-06, 
    4.102747e-06, 4.084191e-06, 4.153529e-06, 4.133779e-06, 4.190954e-06, 
    4.176547e-06, 4.190276e-06, 4.186112e-06, 4.19033e-06, 4.169207e-06, 
    4.178252e-06, 4.159686e-06, 4.087663e-06, 4.108778e-06, 4.045921e-06, 
    4.008294e-06, 3.983395e-06, 3.965757e-06, 3.968249e-06, 3.972999e-06, 
    3.997452e-06, 4.020503e-06, 4.038101e-06, 4.049889e-06, 4.061516e-06, 
    4.096772e-06, 4.115496e-06, 4.157524e-06, 4.149933e-06, 4.1628e-06, 
    4.175115e-06, 4.195812e-06, 4.192404e-06, 4.20153e-06, 4.162465e-06, 
    4.18841e-06, 4.145611e-06, 4.157299e-06, 4.064656e-06, 4.029602e-06, 
    4.014717e-06, 4.001725e-06, 3.970164e-06, 3.991948e-06, 3.983354e-06, 
    4.003815e-06, 4.016833e-06, 4.010394e-06, 4.050211e-06, 4.034712e-06, 
    4.116606e-06, 4.081255e-06, 4.173678e-06, 4.151491e-06, 4.179003e-06, 
    4.164957e-06, 4.189033e-06, 4.167362e-06, 4.204931e-06, 4.213125e-06, 
    4.207524e-06, 4.229063e-06, 4.166162e-06, 4.190274e-06, 4.010212e-06, 
    4.011262e-06, 4.016157e-06, 3.994656e-06, 3.993343e-06, 3.973688e-06, 
    3.991177e-06, 3.998633e-06, 4.017591e-06, 4.028816e-06, 4.0395e-06, 
    4.063029e-06, 4.089365e-06, 4.126307e-06, 4.152928e-06, 4.170808e-06, 
    4.159842e-06, 4.169523e-06, 4.158701e-06, 4.153633e-06, 4.210052e-06, 
    4.178335e-06, 4.225963e-06, 4.223323e-06, 4.201746e-06, 4.22362e-06, 
    4.012e-06, 4.005959e-06, 3.985003e-06, 4.001399e-06, 3.97155e-06, 
    3.988244e-06, 3.997854e-06, 4.035031e-06, 4.043222e-06, 4.050816e-06, 
    4.065836e-06, 4.08514e-06, 4.119086e-06, 4.148713e-06, 4.175833e-06, 
    4.173844e-06, 4.174544e-06, 4.180607e-06, 4.165589e-06, 4.183075e-06, 
    4.18601e-06, 4.178334e-06, 4.222969e-06, 4.2102e-06, 4.223266e-06, 
    4.214951e-06, 4.007923e-06, 4.018093e-06, 4.012596e-06, 4.022934e-06, 
    4.015647e-06, 4.048079e-06, 4.057822e-06, 4.103538e-06, 4.084759e-06, 
    4.114668e-06, 4.087795e-06, 4.09255e-06, 4.115635e-06, 4.089247e-06, 
    4.147073e-06, 4.107826e-06, 4.180843e-06, 4.141521e-06, 4.183312e-06, 
    4.175715e-06, 4.188298e-06, 4.199576e-06, 4.213786e-06, 4.240045e-06, 
    4.23396e-06, 4.255959e-06, 4.033275e-06, 4.046498e-06, 4.045338e-06, 
    4.059195e-06, 4.069454e-06, 4.09173e-06, 4.127549e-06, 4.114067e-06, 
    4.138835e-06, 4.143812e-06, 4.106192e-06, 4.129271e-06, 4.05536e-06, 
    4.067263e-06, 4.060178e-06, 4.034315e-06, 4.117166e-06, 4.074563e-06, 
    4.153368e-06, 4.130191e-06, 4.197967e-06, 4.164205e-06, 4.230611e-06, 
    4.259105e-06, 4.28601e-06, 4.317503e-06, 4.053727e-06, 4.044733e-06, 
    4.060846e-06, 4.08317e-06, 4.103938e-06, 4.131603e-06, 4.13444e-06, 
    4.139631e-06, 4.153093e-06, 4.164422e-06, 4.141268e-06, 4.167264e-06, 
    4.070016e-06, 4.120874e-06, 4.041331e-06, 4.065215e-06, 4.081855e-06, 
    4.074557e-06, 4.112529e-06, 4.121496e-06, 4.15801e-06, 4.139122e-06, 
    4.252062e-06, 4.201954e-06, 4.341555e-06, 4.302371e-06, 4.041592e-06, 
    4.053698e-06, 4.095932e-06, 4.075817e-06, 4.133455e-06, 4.147687e-06, 
    4.159275e-06, 4.174097e-06, 4.175702e-06, 4.184495e-06, 4.170089e-06, 
    4.183928e-06, 4.131662e-06, 4.154988e-06, 4.091102e-06, 4.106614e-06, 
    4.099476e-06, 4.09165e-06, 4.115824e-06, 4.141631e-06, 4.14219e-06, 
    4.150477e-06, 4.173849e-06, 4.133689e-06, 4.258531e-06, 4.181255e-06, 
    4.066914e-06, 4.09029e-06, 4.093642e-06, 4.084577e-06, 4.146259e-06, 
    4.123868e-06, 4.184282e-06, 4.167923e-06, 4.194741e-06, 4.181406e-06, 
    4.179445e-06, 4.162346e-06, 4.151712e-06, 4.124892e-06, 4.103121e-06, 
    4.085892e-06, 4.089896e-06, 4.108831e-06, 4.143213e-06, 4.175844e-06, 
    4.168687e-06, 4.192701e-06, 4.129265e-06, 4.155817e-06, 4.145544e-06, 
    4.172351e-06, 4.113707e-06, 4.163603e-06, 4.100988e-06, 4.106465e-06, 
    4.123424e-06, 4.157615e-06, 4.165205e-06, 4.173301e-06, 4.168306e-06, 
    4.144089e-06, 4.140129e-06, 4.123013e-06, 4.118288e-06, 4.105273e-06, 
    4.094505e-06, 4.10434e-06, 4.114678e-06, 4.144102e-06, 4.170682e-06, 
    4.199736e-06, 4.20686e-06, 4.240905e-06, 4.213173e-06, 4.258961e-06, 
    4.220005e-06, 4.287532e-06, 4.166512e-06, 4.218877e-06, 4.124199e-06, 
    4.134362e-06, 4.15276e-06, 4.195088e-06, 4.172224e-06, 4.198972e-06, 
    4.139975e-06, 4.109481e-06, 4.101614e-06, 4.086937e-06, 4.10195e-06, 
    4.100728e-06, 4.115112e-06, 4.110488e-06, 4.14508e-06, 4.126486e-06, 
    4.179394e-06, 4.198762e-06, 4.253649e-06, 4.28742e-06, 4.321911e-06, 
    4.337166e-06, 4.341813e-06, 4.343756e-06,
  3.78041e-06, 3.813993e-06, 3.807456e-06, 3.834614e-06, 3.81954e-06, 
    3.837337e-06, 3.78721e-06, 3.815328e-06, 3.797368e-06, 3.78343e-06, 
    3.887551e-06, 3.835828e-06, 3.94161e-06, 3.908388e-06, 3.992074e-06, 
    3.936429e-06, 4.003335e-06, 3.990468e-06, 4.029258e-06, 4.018129e-06, 
    4.067907e-06, 4.034398e-06, 4.093818e-06, 4.059896e-06, 4.065193e-06, 
    4.033294e-06, 3.846217e-06, 3.881094e-06, 3.844154e-06, 3.849118e-06, 
    3.846891e-06, 3.81985e-06, 3.806251e-06, 3.777851e-06, 3.783001e-06, 
    3.803865e-06, 3.851351e-06, 3.835206e-06, 3.87596e-06, 3.875038e-06, 
    3.920619e-06, 3.900039e-06, 3.976995e-06, 3.955059e-06, 4.018593e-06, 
    4.002574e-06, 4.01784e-06, 4.013209e-06, 4.0179e-06, 3.994417e-06, 
    4.004471e-06, 3.983835e-06, 3.903889e-06, 3.927311e-06, 3.85763e-06, 
    3.815984e-06, 3.78844e-06, 3.768944e-06, 3.771698e-06, 3.776949e-06, 
    3.803987e-06, 3.829487e-06, 3.848968e-06, 3.862023e-06, 3.874905e-06, 
    3.914e-06, 3.934769e-06, 3.981435e-06, 3.973e-06, 3.987298e-06, 
    4.000982e-06, 4.023997e-06, 4.020206e-06, 4.030358e-06, 3.986923e-06, 
    4.015767e-06, 3.968197e-06, 3.981183e-06, 3.878397e-06, 3.839559e-06, 
    3.823091e-06, 3.808711e-06, 3.773815e-06, 3.797898e-06, 3.788396e-06, 
    3.811022e-06, 3.825427e-06, 3.8183e-06, 3.86238e-06, 3.845217e-06, 
    3.936001e-06, 3.896786e-06, 3.999385e-06, 3.974731e-06, 4.005304e-06, 
    3.989692e-06, 4.016458e-06, 3.992365e-06, 4.034141e-06, 4.04326e-06, 
    4.037027e-06, 4.060998e-06, 3.991031e-06, 4.017838e-06, 3.818099e-06, 
    3.819261e-06, 3.824678e-06, 3.800893e-06, 3.799441e-06, 3.777709e-06, 
    3.797045e-06, 3.805291e-06, 3.826263e-06, 3.838689e-06, 3.850519e-06, 
    3.876583e-06, 3.905779e-06, 3.946765e-06, 3.976327e-06, 3.996194e-06, 
    3.984008e-06, 3.994766e-06, 3.98274e-06, 3.977109e-06, 4.039841e-06, 
    4.004564e-06, 4.057546e-06, 4.054607e-06, 4.030599e-06, 4.054938e-06, 
    3.820077e-06, 3.813393e-06, 3.790218e-06, 3.808349e-06, 3.775346e-06, 
    3.793803e-06, 3.804432e-06, 3.845572e-06, 3.85464e-06, 3.863052e-06, 
    3.879692e-06, 3.901092e-06, 3.938751e-06, 3.971646e-06, 4.001779e-06, 
    3.999568e-06, 4.000347e-06, 4.007089e-06, 3.990395e-06, 4.009833e-06, 
    4.013097e-06, 4.004562e-06, 4.054214e-06, 4.040002e-06, 4.054545e-06, 
    4.045289e-06, 3.815565e-06, 3.826819e-06, 3.820736e-06, 3.832178e-06, 
    3.824115e-06, 3.860023e-06, 3.870817e-06, 3.9215e-06, 3.900669e-06, 
    3.933848e-06, 3.904035e-06, 3.90931e-06, 3.934927e-06, 3.905644e-06, 
    3.969827e-06, 3.92626e-06, 4.007351e-06, 3.963663e-06, 4.010095e-06, 
    4.001649e-06, 4.015639e-06, 4.028184e-06, 4.043994e-06, 4.073228e-06, 
    4.066451e-06, 4.090953e-06, 3.843625e-06, 3.85827e-06, 3.856982e-06, 
    3.872334e-06, 3.883703e-06, 3.908399e-06, 3.948143e-06, 3.933179e-06, 
    3.960673e-06, 3.966202e-06, 3.924439e-06, 3.950056e-06, 3.868087e-06, 
    3.881278e-06, 3.873423e-06, 3.844778e-06, 3.936621e-06, 3.88937e-06, 
    3.976816e-06, 3.951077e-06, 4.026394e-06, 3.98886e-06, 4.062722e-06, 
    4.094465e-06, 4.124448e-06, 4.159587e-06, 3.866276e-06, 3.856313e-06, 
    3.874162e-06, 3.898911e-06, 3.921941e-06, 3.952644e-06, 3.955793e-06, 
    3.961557e-06, 3.976509e-06, 3.989097e-06, 3.963378e-06, 3.992256e-06, 
    3.884335e-06, 3.940735e-06, 3.852547e-06, 3.879009e-06, 3.897451e-06, 
    3.889359e-06, 3.93147e-06, 3.941423e-06, 3.981975e-06, 3.960991e-06, 
    4.086618e-06, 4.030833e-06, 4.186435e-06, 4.142701e-06, 3.852834e-06, 
    3.866243e-06, 3.913062e-06, 3.890756e-06, 3.954699e-06, 3.970506e-06, 
    3.983377e-06, 3.999852e-06, 4.001635e-06, 4.011412e-06, 3.995395e-06, 
    4.01078e-06, 3.952709e-06, 3.978616e-06, 3.907701e-06, 3.924909e-06, 
    3.91699e-06, 3.908309e-06, 3.935128e-06, 3.963782e-06, 3.964399e-06, 
    3.973606e-06, 3.999591e-06, 3.954959e-06, 4.093834e-06, 4.007822e-06, 
    3.880887e-06, 3.906807e-06, 3.91052e-06, 3.900466e-06, 3.968919e-06, 
    3.944057e-06, 4.011174e-06, 3.992988e-06, 4.022805e-06, 4.007976e-06, 
    4.005796e-06, 3.98679e-06, 3.974976e-06, 3.945195e-06, 3.921034e-06, 
    3.901924e-06, 3.906364e-06, 3.92737e-06, 3.965538e-06, 4.001794e-06, 
    3.99384e-06, 4.020535e-06, 3.950047e-06, 3.979538e-06, 3.968127e-06, 
    3.99791e-06, 3.93278e-06, 3.9882e-06, 3.918666e-06, 3.924742e-06, 
    3.943564e-06, 3.981539e-06, 3.989967e-06, 3.998968e-06, 3.993413e-06, 
    3.96651e-06, 3.962112e-06, 3.943107e-06, 3.937865e-06, 3.923419e-06, 
    3.911475e-06, 3.922386e-06, 3.933858e-06, 3.966523e-06, 3.996056e-06, 
    4.028363e-06, 4.036287e-06, 4.074193e-06, 4.043319e-06, 4.094315e-06, 
    4.050933e-06, 4.126156e-06, 3.991428e-06, 4.049668e-06, 3.944423e-06, 
    3.955705e-06, 3.976143e-06, 4.023197e-06, 3.997769e-06, 4.027515e-06, 
    3.96194e-06, 3.928093e-06, 3.919361e-06, 3.903084e-06, 3.919734e-06, 
    3.918379e-06, 3.934337e-06, 3.929206e-06, 3.96761e-06, 3.946961e-06, 
    4.005741e-06, 4.027281e-06, 4.088381e-06, 4.126025e-06, 4.1645e-06, 
    4.181531e-06, 4.186721e-06, 4.188891e-06,
  3.868069e-06, 3.904865e-06, 3.897699e-06, 3.927474e-06, 3.910944e-06, 
    3.93046e-06, 3.875516e-06, 3.906329e-06, 3.886645e-06, 3.871375e-06, 
    3.985568e-06, 3.928805e-06, 4.04495e-06, 4.008443e-06, 4.100456e-06, 
    4.039258e-06, 4.11285e-06, 4.098686e-06, 4.14139e-06, 4.129135e-06, 
    4.183986e-06, 4.147053e-06, 4.212558e-06, 4.175152e-06, 4.180993e-06, 
    4.145837e-06, 3.940198e-06, 3.978479e-06, 3.937935e-06, 3.943382e-06, 
    3.940937e-06, 3.911285e-06, 3.896382e-06, 3.865264e-06, 3.870904e-06, 
    3.893765e-06, 3.945832e-06, 3.928121e-06, 3.972833e-06, 3.971821e-06, 
    4.021879e-06, 3.999271e-06, 4.083861e-06, 4.059733e-06, 4.129646e-06, 
    4.112009e-06, 4.128816e-06, 4.123717e-06, 4.128883e-06, 4.103032e-06, 
    4.114098e-06, 4.091386e-06, 4.003501e-06, 4.029233e-06, 3.95272e-06, 
    3.907053e-06, 3.876864e-06, 3.85551e-06, 3.858526e-06, 3.864277e-06, 
    3.893899e-06, 3.92185e-06, 3.943215e-06, 3.957538e-06, 3.971675e-06, 
    4.014613e-06, 4.037431e-06, 4.088748e-06, 4.079465e-06, 4.095198e-06, 
    4.110257e-06, 4.135597e-06, 4.131422e-06, 4.142604e-06, 4.094783e-06, 
    4.126535e-06, 4.074181e-06, 4.088468e-06, 3.975519e-06, 3.932895e-06, 
    3.914842e-06, 3.899076e-06, 3.860845e-06, 3.887227e-06, 3.876817e-06, 
    3.901606e-06, 3.917397e-06, 3.909584e-06, 3.95793e-06, 3.9391e-06, 
    4.038785e-06, 3.9957e-06, 4.108499e-06, 4.081369e-06, 4.115014e-06, 
    4.09783e-06, 4.127296e-06, 4.100772e-06, 4.14677e-06, 4.156818e-06, 
    4.149951e-06, 4.176364e-06, 4.099304e-06, 4.128816e-06, 3.909365e-06, 
    3.910638e-06, 3.916576e-06, 3.890509e-06, 3.888917e-06, 3.865109e-06, 
    3.88629e-06, 3.895327e-06, 3.918314e-06, 3.931941e-06, 3.944916e-06, 
    3.973517e-06, 4.005577e-06, 4.050617e-06, 4.083126e-06, 4.104986e-06, 
    4.091575e-06, 4.103414e-06, 4.09018e-06, 4.083985e-06, 4.153052e-06, 
    4.114201e-06, 4.17256e-06, 4.169321e-06, 4.14287e-06, 4.169685e-06, 
    3.911533e-06, 3.904205e-06, 3.878812e-06, 3.898677e-06, 3.86252e-06, 
    3.882739e-06, 3.894387e-06, 3.939492e-06, 3.949437e-06, 3.958668e-06, 
    3.97693e-06, 4.000427e-06, 4.041807e-06, 4.077978e-06, 4.111133e-06, 
    4.1087e-06, 4.109557e-06, 4.116979e-06, 4.098604e-06, 4.12e-06, 
    4.123596e-06, 4.114197e-06, 4.168886e-06, 4.153227e-06, 4.169251e-06, 
    4.159052e-06, 3.906586e-06, 3.918925e-06, 3.912255e-06, 3.924802e-06, 
    3.91596e-06, 3.955347e-06, 3.967193e-06, 4.02285e-06, 3.999964e-06, 
    4.036418e-06, 4.00366e-06, 4.009455e-06, 4.037609e-06, 4.005427e-06, 
    4.075979e-06, 4.028081e-06, 4.117268e-06, 4.069202e-06, 4.120289e-06, 
    4.11099e-06, 4.126392e-06, 4.14021e-06, 4.157625e-06, 4.18985e-06, 
    4.182377e-06, 4.209396e-06, 3.937354e-06, 3.953422e-06, 3.952007e-06, 
    3.968853e-06, 3.981334e-06, 4.008452e-06, 4.05213e-06, 4.035679e-06, 
    4.065906e-06, 4.071987e-06, 4.026075e-06, 4.054234e-06, 3.964194e-06, 
    3.978675e-06, 3.97005e-06, 3.93862e-06, 4.039466e-06, 3.987558e-06, 
    4.083663e-06, 4.055355e-06, 4.138238e-06, 4.096918e-06, 4.178266e-06, 
    4.213275e-06, 4.246354e-06, 4.285165e-06, 3.962205e-06, 3.951272e-06, 
    3.970859e-06, 3.998035e-06, 4.023331e-06, 4.057079e-06, 4.06054e-06, 
    4.06688e-06, 4.083324e-06, 4.097175e-06, 4.068885e-06, 4.100651e-06, 
    3.982036e-06, 4.043987e-06, 3.947142e-06, 3.976184e-06, 3.996431e-06, 
    3.987544e-06, 4.033801e-06, 4.04474e-06, 4.089341e-06, 4.066256e-06, 
    4.20462e-06, 4.14313e-06, 4.314832e-06, 4.266512e-06, 3.947456e-06, 
    3.962168e-06, 4.013577e-06, 3.989077e-06, 4.059337e-06, 4.076721e-06, 
    4.090881e-06, 4.109014e-06, 4.110975e-06, 4.121739e-06, 4.104107e-06, 
    4.121042e-06, 4.057151e-06, 4.085643e-06, 4.007685e-06, 4.026593e-06, 
    4.017889e-06, 4.008353e-06, 4.037821e-06, 4.069329e-06, 4.070004e-06, 
    4.080133e-06, 4.108738e-06, 4.059623e-06, 4.212587e-06, 4.117798e-06, 
    3.978241e-06, 4.006708e-06, 4.010783e-06, 3.999739e-06, 4.074977e-06, 
    4.047637e-06, 4.121477e-06, 4.101458e-06, 4.134284e-06, 4.117956e-06, 
    4.115556e-06, 4.094637e-06, 4.081639e-06, 4.048889e-06, 4.022335e-06, 
    4.00134e-06, 4.006217e-06, 4.029297e-06, 4.07126e-06, 4.111152e-06, 
    4.102397e-06, 4.131784e-06, 4.054223e-06, 4.086659e-06, 4.074107e-06, 
    4.106875e-06, 4.035242e-06, 4.0962e-06, 4.019731e-06, 4.026408e-06, 
    4.047095e-06, 4.088863e-06, 4.098133e-06, 4.10804e-06, 4.101926e-06, 
    4.072328e-06, 4.06749e-06, 4.046592e-06, 4.040831e-06, 4.024954e-06, 
    4.011831e-06, 4.02382e-06, 4.036428e-06, 4.072341e-06, 4.104837e-06, 
    4.140406e-06, 4.149134e-06, 4.19092e-06, 4.156888e-06, 4.213117e-06, 
    4.165287e-06, 4.248252e-06, 4.099748e-06, 4.163885e-06, 4.048038e-06, 
    4.060444e-06, 4.082926e-06, 4.13472e-06, 4.106721e-06, 4.139475e-06, 
    4.0673e-06, 4.030094e-06, 4.020495e-06, 4.002614e-06, 4.020904e-06, 
    4.019415e-06, 4.036951e-06, 4.031312e-06, 4.073536e-06, 4.050829e-06, 
    4.115496e-06, 4.139216e-06, 4.20656e-06, 4.2481e-06, 4.290588e-06, 
    4.309409e-06, 4.315146e-06, 4.317545e-06,
  4.120389e-06, 4.15886e-06, 4.151365e-06, 4.182512e-06, 4.165217e-06, 
    4.185637e-06, 4.128171e-06, 4.160392e-06, 4.139806e-06, 4.123843e-06, 
    4.243343e-06, 4.183905e-06, 4.305588e-06, 4.267306e-06, 4.363847e-06, 
    4.29962e-06, 4.376864e-06, 4.361985e-06, 4.406853e-06, 4.393972e-06, 
    4.451656e-06, 4.412806e-06, 4.481728e-06, 4.442359e-06, 4.448505e-06, 
    4.411528e-06, 4.195826e-06, 4.235917e-06, 4.193458e-06, 4.19916e-06, 
    4.1966e-06, 4.165574e-06, 4.14999e-06, 4.117456e-06, 4.123351e-06, 
    4.147251e-06, 4.201725e-06, 4.183187e-06, 4.229994e-06, 4.228934e-06, 
    4.281391e-06, 4.257693e-06, 4.346419e-06, 4.321093e-06, 4.394509e-06, 
    4.375979e-06, 4.393638e-06, 4.388279e-06, 4.393708e-06, 4.366549e-06, 
    4.378173e-06, 4.354319e-06, 4.262126e-06, 4.289103e-06, 4.208935e-06, 
    4.161152e-06, 4.129582e-06, 4.107264e-06, 4.110415e-06, 4.116426e-06, 
    4.147392e-06, 4.176625e-06, 4.198983e-06, 4.213978e-06, 4.228782e-06, 
    4.273779e-06, 4.297702e-06, 4.351551e-06, 4.341803e-06, 4.358323e-06, 
    4.374137e-06, 4.400765e-06, 4.396376e-06, 4.40813e-06, 4.357886e-06, 
    4.391242e-06, 4.336256e-06, 4.351255e-06, 4.232817e-06, 4.188183e-06, 
    4.169299e-06, 4.152805e-06, 4.112839e-06, 4.140416e-06, 4.129532e-06, 
    4.15545e-06, 4.171968e-06, 4.163793e-06, 4.214388e-06, 4.194677e-06, 
    4.299122e-06, 4.253953e-06, 4.372291e-06, 4.343803e-06, 4.379136e-06, 
    4.361085e-06, 4.39204e-06, 4.364175e-06, 4.412509e-06, 4.423076e-06, 
    4.415854e-06, 4.443632e-06, 4.362633e-06, 4.393638e-06, 4.163565e-06, 
    4.164897e-06, 4.171108e-06, 4.143847e-06, 4.142182e-06, 4.117294e-06, 
    4.139435e-06, 4.148885e-06, 4.172926e-06, 4.187185e-06, 4.200765e-06, 
    4.230712e-06, 4.264304e-06, 4.311531e-06, 4.345646e-06, 4.368601e-06, 
    4.354516e-06, 4.36695e-06, 4.353053e-06, 4.346547e-06, 4.419115e-06, 
    4.378282e-06, 4.439631e-06, 4.436223e-06, 4.40841e-06, 4.436607e-06, 
    4.165833e-06, 4.158167e-06, 4.131617e-06, 4.152387e-06, 4.114589e-06, 
    4.135723e-06, 4.147903e-06, 4.195089e-06, 4.205496e-06, 4.215161e-06, 
    4.234286e-06, 4.258904e-06, 4.302289e-06, 4.340243e-06, 4.375058e-06, 
    4.372502e-06, 4.373402e-06, 4.3812e-06, 4.361899e-06, 4.384374e-06, 
    4.388153e-06, 4.378277e-06, 4.435766e-06, 4.419298e-06, 4.43615e-06, 
    4.425423e-06, 4.160658e-06, 4.173565e-06, 4.166588e-06, 4.179715e-06, 
    4.170465e-06, 4.211686e-06, 4.224091e-06, 4.282411e-06, 4.258419e-06, 
    4.296638e-06, 4.262292e-06, 4.268367e-06, 4.297891e-06, 4.264144e-06, 
    4.338146e-06, 4.287897e-06, 4.381503e-06, 4.331037e-06, 4.384678e-06, 
    4.374907e-06, 4.39109e-06, 4.405613e-06, 4.423922e-06, 4.457824e-06, 
    4.44996e-06, 4.478396e-06, 4.19285e-06, 4.20967e-06, 4.208187e-06, 
    4.225827e-06, 4.238901e-06, 4.267315e-06, 4.313118e-06, 4.29586e-06, 
    4.327571e-06, 4.333954e-06, 4.285789e-06, 4.315326e-06, 4.220949e-06, 
    4.236117e-06, 4.227081e-06, 4.194176e-06, 4.299835e-06, 4.245422e-06, 
    4.346211e-06, 4.316501e-06, 4.403541e-06, 4.36013e-06, 4.445634e-06, 
    4.482485e-06, 4.517323e-06, 4.558243e-06, 4.218866e-06, 4.207418e-06, 
    4.227927e-06, 4.2564e-06, 4.282913e-06, 4.318309e-06, 4.32194e-06, 
    4.328594e-06, 4.345854e-06, 4.360398e-06, 4.3307e-06, 4.364048e-06, 
    4.239641e-06, 4.304577e-06, 4.203096e-06, 4.233509e-06, 4.254718e-06, 
    4.245405e-06, 4.29389e-06, 4.305364e-06, 4.352173e-06, 4.327938e-06, 
    4.473375e-06, 4.408686e-06, 4.58954e-06, 4.538573e-06, 4.203423e-06, 
    4.218826e-06, 4.272688e-06, 4.247011e-06, 4.320678e-06, 4.338924e-06, 
    4.353788e-06, 4.372833e-06, 4.374891e-06, 4.386202e-06, 4.367677e-06, 
    4.385469e-06, 4.318385e-06, 4.348289e-06, 4.266511e-06, 4.286333e-06, 
    4.277207e-06, 4.26721e-06, 4.298107e-06, 4.331167e-06, 4.331873e-06, 
    4.342506e-06, 4.372554e-06, 4.320978e-06, 4.481768e-06, 4.38207e-06, 
    4.235659e-06, 4.26549e-06, 4.269758e-06, 4.258182e-06, 4.337092e-06, 
    4.308404e-06, 4.385925e-06, 4.364895e-06, 4.399383e-06, 4.382226e-06, 
    4.379705e-06, 4.357733e-06, 4.344085e-06, 4.309717e-06, 4.281869e-06, 
    4.25986e-06, 4.264972e-06, 4.289169e-06, 4.333193e-06, 4.375079e-06, 
    4.365884e-06, 4.396757e-06, 4.315312e-06, 4.349357e-06, 4.336181e-06, 
    4.370585e-06, 4.295403e-06, 4.359383e-06, 4.279137e-06, 4.286138e-06, 
    4.307836e-06, 4.351673e-06, 4.361404e-06, 4.371811e-06, 4.365387e-06, 
    4.334314e-06, 4.329234e-06, 4.307307e-06, 4.301265e-06, 4.284613e-06, 
    4.270856e-06, 4.283425e-06, 4.296648e-06, 4.334326e-06, 4.368445e-06, 
    4.40582e-06, 4.414994e-06, 4.458955e-06, 4.423153e-06, 4.482327e-06, 
    4.431993e-06, 4.519331e-06, 4.363105e-06, 4.430513e-06, 4.308824e-06, 
    4.321839e-06, 4.34544e-06, 4.399846e-06, 4.370424e-06, 4.404844e-06, 
    4.329036e-06, 4.290006e-06, 4.279939e-06, 4.261196e-06, 4.280368e-06, 
    4.278807e-06, 4.297195e-06, 4.291281e-06, 4.33558e-06, 4.311752e-06, 
    4.379642e-06, 4.404571e-06, 4.475412e-06, 4.519166e-06, 4.563958e-06, 
    4.583816e-06, 4.589871e-06, 4.592403e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.77824, 5.778221, 5.778224, 5.778209, 5.778217, 5.778207, 5.778236, 
    5.77822, 5.77823, 5.778238, 5.778179, 5.778208, 5.778149, 5.778167, 
    5.77812, 5.778152, 5.778114, 5.778121, 5.7781, 5.778106, 5.778078, 
    5.778097, 5.778064, 5.778082, 5.77808, 5.778097, 5.778203, 5.778183, 
    5.778203, 5.778201, 5.778202, 5.778217, 5.778225, 5.778241, 5.778238, 
    5.778226, 5.7782, 5.778209, 5.778185, 5.778186, 5.77816, 5.778172, 
    5.778129, 5.778141, 5.778105, 5.778114, 5.778106, 5.778108, 5.778106, 
    5.778119, 5.778113, 5.778125, 5.77817, 5.778156, 5.778196, 5.77822, 
    5.778235, 5.778246, 5.778245, 5.778242, 5.778226, 5.778212, 5.778201, 
    5.778193, 5.778186, 5.778164, 5.778152, 5.778126, 5.778131, 5.778123, 
    5.778115, 5.778102, 5.778104, 5.778099, 5.778123, 5.778107, 5.778133, 
    5.778126, 5.778184, 5.778206, 5.778215, 5.778224, 5.778244, 5.77823, 
    5.778235, 5.778223, 5.778214, 5.778218, 5.778193, 5.778203, 5.778152, 
    5.778174, 5.778116, 5.77813, 5.778113, 5.778121, 5.778107, 5.77812, 
    5.778097, 5.778091, 5.778095, 5.778082, 5.778121, 5.778106, 5.778218, 
    5.778218, 5.778214, 5.778228, 5.778229, 5.778242, 5.77823, 5.778226, 
    5.778214, 5.778207, 5.7782, 5.778185, 5.778169, 5.778145, 5.778129, 
    5.778118, 5.778125, 5.778119, 5.778125, 5.778129, 5.778093, 5.778113, 
    5.778084, 5.778085, 5.778099, 5.778085, 5.778217, 5.778221, 5.778234, 
    5.778224, 5.778243, 5.778232, 5.778226, 5.778203, 5.778198, 5.778193, 
    5.778183, 5.778171, 5.77815, 5.778131, 5.778115, 5.778116, 5.778116, 
    5.778112, 5.778121, 5.77811, 5.778109, 5.778113, 5.778086, 5.778093, 
    5.778085, 5.77809, 5.77822, 5.778214, 5.778217, 5.77821, 5.778215, 
    5.778194, 5.778188, 5.77816, 5.778172, 5.778153, 5.77817, 5.778167, 
    5.778152, 5.778169, 5.778132, 5.778157, 5.778111, 5.778136, 5.77811, 
    5.778115, 5.778107, 5.7781, 5.778091, 5.778075, 5.778079, 5.778065, 
    5.778204, 5.778195, 5.778196, 5.778188, 5.778181, 5.778167, 5.778145, 
    5.778153, 5.778138, 5.778135, 5.778158, 5.778144, 5.77819, 5.778183, 
    5.778187, 5.778203, 5.778151, 5.778178, 5.778129, 5.778143, 5.778101, 
    5.778122, 5.778081, 5.778063, 5.778047, 5.778027, 5.778191, 5.778197, 
    5.778186, 5.778172, 5.77816, 5.778142, 5.778141, 5.778137, 5.778129, 
    5.778122, 5.778136, 5.77812, 5.778181, 5.778149, 5.778199, 5.778184, 
    5.778173, 5.778178, 5.778154, 5.778149, 5.778126, 5.778138, 5.778068, 
    5.778099, 5.778013, 5.778037, 5.778199, 5.778191, 5.778164, 5.778177, 
    5.778141, 5.778132, 5.778125, 5.778116, 5.778115, 5.77811, 5.778118, 
    5.77811, 5.778142, 5.778128, 5.778168, 5.778158, 5.778162, 5.778167, 
    5.778152, 5.778136, 5.778136, 5.778131, 5.778116, 5.778141, 5.778063, 
    5.778111, 5.778183, 5.778168, 5.778166, 5.778172, 5.778133, 5.778147, 
    5.77811, 5.77812, 5.778103, 5.778111, 5.778112, 5.778123, 5.77813, 
    5.778146, 5.77816, 5.778171, 5.778168, 5.778156, 5.778135, 5.778115, 
    5.778119, 5.778104, 5.778144, 5.778127, 5.778133, 5.778117, 5.778153, 
    5.778122, 5.778162, 5.778158, 5.778147, 5.778126, 5.778121, 5.778116, 
    5.77812, 5.778134, 5.778137, 5.778148, 5.778151, 5.778159, 5.778165, 
    5.778159, 5.778153, 5.778134, 5.778118, 5.7781, 5.778095, 5.778074, 
    5.778091, 5.778063, 5.778087, 5.778046, 5.778121, 5.778088, 5.778147, 
    5.778141, 5.778129, 5.778103, 5.778117, 5.7781, 5.778137, 5.778156, 
    5.778161, 5.77817, 5.778161, 5.778162, 5.778152, 5.778155, 5.778134, 
    5.778145, 5.778112, 5.7781, 5.778067, 5.778046, 5.778025, 5.778015, 
    5.778012, 5.778011 ;

 SOIL1C_TO_SOIL2C =
  3.099197e-08, 3.112855e-08, 3.1102e-08, 3.121216e-08, 3.115106e-08, 
    3.122319e-08, 3.101967e-08, 3.113397e-08, 3.1061e-08, 3.100427e-08, 
    3.142594e-08, 3.121708e-08, 3.164294e-08, 3.150972e-08, 3.184439e-08, 
    3.162221e-08, 3.18892e-08, 3.183799e-08, 3.199213e-08, 3.194797e-08, 
    3.214512e-08, 3.201251e-08, 3.224732e-08, 3.211345e-08, 3.213439e-08, 
    3.200814e-08, 3.125912e-08, 3.139994e-08, 3.125077e-08, 3.127085e-08, 
    3.126184e-08, 3.115231e-08, 3.109712e-08, 3.098154e-08, 3.100252e-08, 
    3.108741e-08, 3.127988e-08, 3.121455e-08, 3.137922e-08, 3.13755e-08, 
    3.155882e-08, 3.147616e-08, 3.17843e-08, 3.169673e-08, 3.194982e-08, 
    3.188616e-08, 3.194683e-08, 3.192843e-08, 3.194706e-08, 3.185371e-08, 
    3.189371e-08, 3.181157e-08, 3.149164e-08, 3.158566e-08, 3.130525e-08, 
    3.113665e-08, 3.102468e-08, 3.094522e-08, 3.095645e-08, 3.097787e-08, 
    3.108791e-08, 3.119139e-08, 3.127024e-08, 3.132299e-08, 3.137496e-08, 
    3.153227e-08, 3.161555e-08, 3.180201e-08, 3.176837e-08, 3.182537e-08, 
    3.187983e-08, 3.197126e-08, 3.195622e-08, 3.19965e-08, 3.182387e-08, 
    3.19386e-08, 3.17492e-08, 3.1801e-08, 3.138907e-08, 3.123218e-08, 
    3.116547e-08, 3.110711e-08, 3.096509e-08, 3.106316e-08, 3.10245e-08, 
    3.111648e-08, 3.117493e-08, 3.114602e-08, 3.132443e-08, 3.125507e-08, 
    3.162048e-08, 3.146308e-08, 3.187348e-08, 3.177527e-08, 3.189702e-08, 
    3.18349e-08, 3.194134e-08, 3.184554e-08, 3.20115e-08, 3.204763e-08, 
    3.202294e-08, 3.21178e-08, 3.184023e-08, 3.194682e-08, 3.114521e-08, 
    3.114993e-08, 3.117189e-08, 3.107534e-08, 3.106943e-08, 3.098096e-08, 
    3.105968e-08, 3.109321e-08, 3.117832e-08, 3.122866e-08, 3.127651e-08, 
    3.138173e-08, 3.149924e-08, 3.166357e-08, 3.178164e-08, 3.186078e-08, 
    3.181225e-08, 3.18551e-08, 3.18072e-08, 3.178475e-08, 3.203409e-08, 
    3.189408e-08, 3.210416e-08, 3.209253e-08, 3.199746e-08, 3.209384e-08, 
    3.115323e-08, 3.112611e-08, 3.103191e-08, 3.110563e-08, 3.097133e-08, 
    3.10465e-08, 3.108972e-08, 3.125651e-08, 3.129317e-08, 3.132714e-08, 
    3.139426e-08, 3.148039e-08, 3.163149e-08, 3.176297e-08, 3.1883e-08, 
    3.187421e-08, 3.18773e-08, 3.190411e-08, 3.18377e-08, 3.191502e-08, 
    3.192799e-08, 3.189407e-08, 3.209098e-08, 3.203472e-08, 3.209228e-08, 
    3.205566e-08, 3.113493e-08, 3.118058e-08, 3.115591e-08, 3.120229e-08, 
    3.116961e-08, 3.131492e-08, 3.135849e-08, 3.156236e-08, 3.14787e-08, 
    3.161186e-08, 3.149222e-08, 3.151342e-08, 3.161619e-08, 3.149869e-08, 
    3.175572e-08, 3.158145e-08, 3.190516e-08, 3.173112e-08, 3.191606e-08, 
    3.188248e-08, 3.193808e-08, 3.198788e-08, 3.205053e-08, 3.216612e-08, 
    3.213936e-08, 3.223603e-08, 3.124863e-08, 3.130784e-08, 3.130263e-08, 
    3.13646e-08, 3.141042e-08, 3.150976e-08, 3.166907e-08, 3.160917e-08, 
    3.171916e-08, 3.174124e-08, 3.157414e-08, 3.167673e-08, 3.134747e-08, 
    3.140066e-08, 3.136899e-08, 3.12533e-08, 3.162296e-08, 3.143325e-08, 
    3.178359e-08, 3.168081e-08, 3.198078e-08, 3.183159e-08, 3.212462e-08, 
    3.224988e-08, 3.23678e-08, 3.250558e-08, 3.134016e-08, 3.129993e-08, 
    3.137197e-08, 3.147163e-08, 3.156412e-08, 3.168708e-08, 3.169966e-08, 
    3.172269e-08, 3.178236e-08, 3.183253e-08, 3.172997e-08, 3.18451e-08, 
    3.141299e-08, 3.163943e-08, 3.128471e-08, 3.139152e-08, 3.146576e-08, 
    3.14332e-08, 3.160232e-08, 3.164218e-08, 3.180416e-08, 3.172043e-08, 
    3.221896e-08, 3.199839e-08, 3.26105e-08, 3.243943e-08, 3.128587e-08, 
    3.134002e-08, 3.152849e-08, 3.143882e-08, 3.169529e-08, 3.175841e-08, 
    3.180974e-08, 3.187534e-08, 3.188243e-08, 3.19213e-08, 3.18576e-08, 
    3.191878e-08, 3.168734e-08, 3.179077e-08, 3.150695e-08, 3.157603e-08, 
    3.154425e-08, 3.150939e-08, 3.161697e-08, 3.173158e-08, 3.173404e-08, 
    3.177079e-08, 3.187433e-08, 3.169633e-08, 3.224742e-08, 3.190706e-08, 
    3.139907e-08, 3.150337e-08, 3.151828e-08, 3.147787e-08, 3.175209e-08, 
    3.165272e-08, 3.192035e-08, 3.184802e-08, 3.196653e-08, 3.190764e-08, 
    3.189898e-08, 3.182334e-08, 3.177625e-08, 3.165728e-08, 3.156049e-08, 
    3.148374e-08, 3.150158e-08, 3.158589e-08, 3.17386e-08, 3.188307e-08, 
    3.185142e-08, 3.195753e-08, 3.167669e-08, 3.179444e-08, 3.174893e-08, 
    3.186761e-08, 3.160757e-08, 3.182899e-08, 3.155098e-08, 3.157535e-08, 
    3.165075e-08, 3.180243e-08, 3.1836e-08, 3.187182e-08, 3.184972e-08, 
    3.174247e-08, 3.172491e-08, 3.164892e-08, 3.162794e-08, 3.157005e-08, 
    3.152211e-08, 3.156591e-08, 3.16119e-08, 3.174252e-08, 3.186024e-08, 
    3.198858e-08, 3.202e-08, 3.216995e-08, 3.204788e-08, 3.224931e-08, 
    3.207804e-08, 3.237454e-08, 3.184183e-08, 3.207301e-08, 3.165419e-08, 
    3.169931e-08, 3.178091e-08, 3.19681e-08, 3.186705e-08, 3.198523e-08, 
    3.172422e-08, 3.15888e-08, 3.155377e-08, 3.14884e-08, 3.155526e-08, 
    3.154982e-08, 3.16138e-08, 3.159325e-08, 3.174686e-08, 3.166435e-08, 
    3.189876e-08, 3.19843e-08, 3.22259e-08, 3.2374e-08, 3.252478e-08, 
    3.259135e-08, 3.261161e-08, 3.262008e-08 ;

 SOIL1C_TO_SOIL3C =
  3.675989e-10, 3.692194e-10, 3.689044e-10, 3.702115e-10, 3.694864e-10, 
    3.703423e-10, 3.679275e-10, 3.692837e-10, 3.684179e-10, 3.677448e-10, 
    3.727481e-10, 3.702698e-10, 3.753229e-10, 3.737421e-10, 3.777133e-10, 
    3.750769e-10, 3.782449e-10, 3.776373e-10, 3.794663e-10, 3.789423e-10, 
    3.812817e-10, 3.797082e-10, 3.824945e-10, 3.80906e-10, 3.811544e-10, 
    3.796563e-10, 3.707686e-10, 3.724395e-10, 3.706696e-10, 3.709079e-10, 
    3.708009e-10, 3.695014e-10, 3.688465e-10, 3.674751e-10, 3.67724e-10, 
    3.687313e-10, 3.71015e-10, 3.702398e-10, 3.721936e-10, 3.721495e-10, 
    3.743247e-10, 3.73344e-10, 3.770003e-10, 3.759611e-10, 3.789642e-10, 
    3.782089e-10, 3.789287e-10, 3.787105e-10, 3.789316e-10, 3.778239e-10, 
    3.782984e-10, 3.773238e-10, 3.735276e-10, 3.746432e-10, 3.71316e-10, 
    3.693155e-10, 3.679869e-10, 3.670441e-10, 3.671774e-10, 3.674315e-10, 
    3.687372e-10, 3.69965e-10, 3.709006e-10, 3.715265e-10, 3.721432e-10, 
    3.740097e-10, 3.749979e-10, 3.772104e-10, 3.768112e-10, 3.774875e-10, 
    3.781338e-10, 3.792188e-10, 3.790402e-10, 3.795182e-10, 3.774697e-10, 
    3.788311e-10, 3.765837e-10, 3.771984e-10, 3.723106e-10, 3.70449e-10, 
    3.696575e-10, 3.689649e-10, 3.672799e-10, 3.684435e-10, 3.679848e-10, 
    3.690762e-10, 3.697697e-10, 3.694267e-10, 3.715436e-10, 3.707206e-10, 
    3.750564e-10, 3.731888e-10, 3.780584e-10, 3.768931e-10, 3.783378e-10, 
    3.776006e-10, 3.788637e-10, 3.777269e-10, 3.796961e-10, 3.801249e-10, 
    3.798319e-10, 3.809575e-10, 3.776639e-10, 3.789287e-10, 3.694171e-10, 
    3.69473e-10, 3.697336e-10, 3.68588e-10, 3.68518e-10, 3.674682e-10, 
    3.684023e-10, 3.688001e-10, 3.698099e-10, 3.704072e-10, 3.70975e-10, 
    3.722234e-10, 3.736178e-10, 3.755677e-10, 3.769687e-10, 3.779077e-10, 
    3.773319e-10, 3.778403e-10, 3.77272e-10, 3.770056e-10, 3.799642e-10, 
    3.783029e-10, 3.807956e-10, 3.806577e-10, 3.795295e-10, 3.806733e-10, 
    3.695123e-10, 3.691904e-10, 3.680728e-10, 3.689474e-10, 3.673539e-10, 
    3.682459e-10, 3.687587e-10, 3.707377e-10, 3.711726e-10, 3.715758e-10, 
    3.723722e-10, 3.733941e-10, 3.751871e-10, 3.767471e-10, 3.781714e-10, 
    3.78067e-10, 3.781038e-10, 3.78422e-10, 3.776338e-10, 3.785513e-10, 
    3.787053e-10, 3.783027e-10, 3.806392e-10, 3.799717e-10, 3.806548e-10, 
    3.802202e-10, 3.692951e-10, 3.698367e-10, 3.69544e-10, 3.700944e-10, 
    3.697066e-10, 3.714307e-10, 3.719477e-10, 3.743668e-10, 3.73374e-10, 
    3.749541e-10, 3.735346e-10, 3.737861e-10, 3.750055e-10, 3.736113e-10, 
    3.766611e-10, 3.745933e-10, 3.784343e-10, 3.763692e-10, 3.785637e-10, 
    3.781652e-10, 3.78825e-10, 3.794159e-10, 3.801593e-10, 3.81531e-10, 
    3.812133e-10, 3.823605e-10, 3.706442e-10, 3.713467e-10, 3.712849e-10, 
    3.720202e-10, 3.725639e-10, 3.737426e-10, 3.75633e-10, 3.749221e-10, 
    3.762272e-10, 3.764893e-10, 3.745065e-10, 3.757238e-10, 3.718169e-10, 
    3.724481e-10, 3.720723e-10, 3.706996e-10, 3.750859e-10, 3.728347e-10, 
    3.769918e-10, 3.757722e-10, 3.793316e-10, 3.775614e-10, 3.810385e-10, 
    3.825249e-10, 3.839241e-10, 3.855591e-10, 3.717302e-10, 3.712528e-10, 
    3.721076e-10, 3.732902e-10, 3.743876e-10, 3.758466e-10, 3.759959e-10, 
    3.762692e-10, 3.769772e-10, 3.775725e-10, 3.763556e-10, 3.777217e-10, 
    3.725943e-10, 3.752813e-10, 3.710723e-10, 3.723396e-10, 3.732205e-10, 
    3.728342e-10, 3.748409e-10, 3.753139e-10, 3.772359e-10, 3.762423e-10, 
    3.82158e-10, 3.795406e-10, 3.868041e-10, 3.847741e-10, 3.710861e-10, 
    3.717286e-10, 3.739649e-10, 3.729008e-10, 3.75944e-10, 3.766931e-10, 
    3.773021e-10, 3.780805e-10, 3.781646e-10, 3.786258e-10, 3.7787e-10, 
    3.78596e-10, 3.758497e-10, 3.770769e-10, 3.737093e-10, 3.745289e-10, 
    3.741519e-10, 3.737383e-10, 3.750148e-10, 3.763747e-10, 3.764039e-10, 
    3.768399e-10, 3.780685e-10, 3.759563e-10, 3.824956e-10, 3.784569e-10, 
    3.724293e-10, 3.736668e-10, 3.738437e-10, 3.733643e-10, 3.76618e-10, 
    3.75439e-10, 3.786146e-10, 3.777563e-10, 3.791626e-10, 3.784638e-10, 
    3.78361e-10, 3.774635e-10, 3.769047e-10, 3.754931e-10, 3.743445e-10, 
    3.734338e-10, 3.736456e-10, 3.74646e-10, 3.764579e-10, 3.781722e-10, 
    3.777967e-10, 3.790557e-10, 3.757233e-10, 3.771206e-10, 3.765805e-10, 
    3.779888e-10, 3.749032e-10, 3.775305e-10, 3.742317e-10, 3.745209e-10, 
    3.754156e-10, 3.772153e-10, 3.776136e-10, 3.780387e-10, 3.777764e-10, 
    3.765039e-10, 3.762955e-10, 3.753939e-10, 3.751449e-10, 3.744579e-10, 
    3.738892e-10, 3.744088e-10, 3.749545e-10, 3.765045e-10, 3.779013e-10, 
    3.794243e-10, 3.79797e-10, 3.815764e-10, 3.801278e-10, 3.825181e-10, 
    3.804857e-10, 3.840041e-10, 3.776829e-10, 3.804261e-10, 3.754563e-10, 
    3.759917e-10, 3.769601e-10, 3.791812e-10, 3.779821e-10, 3.793845e-10, 
    3.762873e-10, 3.746805e-10, 3.742648e-10, 3.734892e-10, 3.742825e-10, 
    3.74218e-10, 3.749772e-10, 3.747332e-10, 3.76556e-10, 3.755769e-10, 
    3.783584e-10, 3.793734e-10, 3.822403e-10, 3.839978e-10, 3.85787e-10, 
    3.865769e-10, 3.868173e-10, 3.869178e-10 ;

 SOIL1C_vr =
  19.98109, 19.98104, 19.98105, 19.98101, 19.98103, 19.981, 19.98108, 
    19.98104, 19.98107, 19.98109, 19.98093, 19.98101, 19.98085, 19.9809, 
    19.98077, 19.98085, 19.98075, 19.98077, 19.98071, 19.98073, 19.98066, 
    19.98071, 19.98062, 19.98067, 19.98066, 19.98071, 19.98099, 19.98094, 
    19.981, 19.98099, 19.98099, 19.98103, 19.98105, 19.9811, 19.98109, 
    19.98106, 19.98098, 19.98101, 19.98095, 19.98095, 19.98088, 19.98091, 
    19.98079, 19.98083, 19.98073, 19.98075, 19.98073, 19.98074, 19.98073, 
    19.98077, 19.98075, 19.98078, 19.9809, 19.98087, 19.98097, 19.98104, 
    19.98108, 19.98111, 19.98111, 19.9811, 19.98106, 19.98102, 19.98099, 
    19.98097, 19.98095, 19.98089, 19.98086, 19.98079, 19.9808, 19.98078, 
    19.98076, 19.98072, 19.98073, 19.98071, 19.98078, 19.98074, 19.98081, 
    19.98079, 19.98094, 19.981, 19.98103, 19.98105, 19.9811, 19.98107, 
    19.98108, 19.98104, 19.98102, 19.98103, 19.98097, 19.98099, 19.98086, 
    19.98092, 19.98076, 19.9808, 19.98075, 19.98077, 19.98073, 19.98077, 
    19.98071, 19.98069, 19.9807, 19.98067, 19.98077, 19.98073, 19.98104, 
    19.98103, 19.98102, 19.98106, 19.98106, 19.9811, 19.98107, 19.98105, 
    19.98102, 19.981, 19.98099, 19.98095, 19.9809, 19.98084, 19.98079, 
    19.98076, 19.98078, 19.98077, 19.98079, 19.98079, 19.9807, 19.98075, 
    19.98067, 19.98068, 19.98071, 19.98068, 19.98103, 19.98104, 19.98108, 
    19.98105, 19.9811, 19.98107, 19.98106, 19.98099, 19.98098, 19.98097, 
    19.98094, 19.98091, 19.98085, 19.9808, 19.98076, 19.98076, 19.98076, 
    19.98075, 19.98077, 19.98075, 19.98074, 19.98075, 19.98068, 19.9807, 
    19.98068, 19.98069, 19.98104, 19.98102, 19.98103, 19.98101, 19.98103, 
    19.98097, 19.98095, 19.98088, 19.98091, 19.98086, 19.9809, 19.9809, 
    19.98086, 19.9809, 19.9808, 19.98087, 19.98075, 19.98081, 19.98074, 
    19.98076, 19.98074, 19.98072, 19.98069, 19.98065, 19.98066, 19.98062, 
    19.981, 19.98097, 19.98097, 19.98095, 19.98093, 19.9809, 19.98084, 
    19.98086, 19.98082, 19.98081, 19.98087, 19.98083, 19.98096, 19.98094, 
    19.98095, 19.98099, 19.98085, 19.98093, 19.98079, 19.98083, 19.98072, 
    19.98078, 19.98067, 19.98062, 19.98058, 19.98052, 19.98096, 19.98098, 
    19.98095, 19.98091, 19.98088, 19.98083, 19.98083, 19.98082, 19.98079, 
    19.98078, 19.98081, 19.98077, 19.98093, 19.98085, 19.98098, 19.98094, 
    19.98091, 19.98093, 19.98086, 19.98085, 19.98079, 19.98082, 19.98063, 
    19.98071, 19.98048, 19.98055, 19.98098, 19.98096, 19.98089, 19.98092, 
    19.98083, 19.9808, 19.98078, 19.98076, 19.98076, 19.98074, 19.98077, 
    19.98074, 19.98083, 19.98079, 19.9809, 19.98087, 19.98088, 19.9809, 
    19.98086, 19.98081, 19.98081, 19.9808, 19.98076, 19.98083, 19.98062, 
    19.98075, 19.98094, 19.9809, 19.98089, 19.98091, 19.98081, 19.98084, 
    19.98074, 19.98077, 19.98072, 19.98075, 19.98075, 19.98078, 19.9808, 
    19.98084, 19.98088, 19.98091, 19.9809, 19.98087, 19.98081, 19.98076, 
    19.98077, 19.98073, 19.98083, 19.98079, 19.98081, 19.98076, 19.98086, 
    19.98078, 19.98088, 19.98087, 19.98084, 19.98079, 19.98077, 19.98076, 
    19.98077, 19.98081, 19.98082, 19.98084, 19.98085, 19.98088, 19.98089, 
    19.98088, 19.98086, 19.98081, 19.98076, 19.98072, 19.98071, 19.98065, 
    19.98069, 19.98062, 19.98068, 19.98057, 19.98077, 19.98068, 19.98084, 
    19.98083, 19.98079, 19.98072, 19.98076, 19.98072, 19.98082, 19.98087, 
    19.98088, 19.98091, 19.98088, 19.98088, 19.98086, 19.98087, 19.98081, 
    19.98084, 19.98075, 19.98072, 19.98063, 19.98057, 19.98052, 19.98049, 
    19.98048, 19.98048,
  19.98328, 19.98321, 19.98323, 19.98318, 19.9832, 19.98317, 19.98326, 
    19.98321, 19.98325, 19.98327, 19.98308, 19.98317, 19.98298, 19.98304, 
    19.98288, 19.98298, 19.98286, 19.98288, 19.98281, 19.98283, 19.98274, 
    19.9828, 19.98269, 19.98276, 19.98275, 19.98281, 19.98315, 19.98309, 
    19.98316, 19.98315, 19.98315, 19.9832, 19.98323, 19.98328, 19.98327, 
    19.98323, 19.98314, 19.98317, 19.9831, 19.9831, 19.98301, 19.98305, 
    19.98291, 19.98295, 19.98283, 19.98286, 19.98283, 19.98284, 19.98283, 
    19.98288, 19.98286, 19.98289, 19.98304, 19.983, 19.98313, 19.98321, 
    19.98326, 19.9833, 19.98329, 19.98328, 19.98323, 19.98318, 19.98315, 
    19.98312, 19.9831, 19.98303, 19.98299, 19.9829, 19.98292, 19.98289, 
    19.98286, 19.98282, 19.98283, 19.98281, 19.98289, 19.98284, 19.98293, 
    19.9829, 19.98309, 19.98317, 19.9832, 19.98322, 19.98329, 19.98324, 
    19.98326, 19.98322, 19.98319, 19.98321, 19.98312, 19.98315, 19.98298, 
    19.98306, 19.98287, 19.98291, 19.98286, 19.98289, 19.98284, 19.98288, 
    19.9828, 19.98279, 19.9828, 19.98275, 19.98288, 19.98283, 19.98321, 
    19.9832, 19.98319, 19.98324, 19.98324, 19.98328, 19.98325, 19.98323, 
    19.98319, 19.98317, 19.98314, 19.9831, 19.98304, 19.98297, 19.98291, 
    19.98287, 19.98289, 19.98288, 19.9829, 19.98291, 19.98279, 19.98286, 
    19.98276, 19.98277, 19.98281, 19.98277, 19.9832, 19.98322, 19.98326, 
    19.98322, 19.98329, 19.98325, 19.98323, 19.98315, 19.98314, 19.98312, 
    19.98309, 19.98305, 19.98298, 19.98292, 19.98286, 19.98287, 19.98286, 
    19.98285, 19.98288, 19.98285, 19.98284, 19.98286, 19.98277, 19.98279, 
    19.98277, 19.98278, 19.98321, 19.98319, 19.9832, 19.98318, 19.98319, 
    19.98313, 19.98311, 19.98301, 19.98305, 19.98299, 19.98304, 19.98303, 
    19.98299, 19.98304, 19.98292, 19.983, 19.98285, 19.98293, 19.98285, 
    19.98286, 19.98284, 19.98281, 19.98278, 19.98273, 19.98274, 19.9827, 
    19.98316, 19.98313, 19.98313, 19.9831, 19.98308, 19.98304, 19.98296, 
    19.98299, 19.98294, 19.98293, 19.98301, 19.98296, 19.98311, 19.98309, 
    19.9831, 19.98316, 19.98298, 19.98307, 19.98291, 19.98296, 19.98282, 
    19.98289, 19.98275, 19.98269, 19.98264, 19.98257, 19.98312, 19.98313, 
    19.9831, 19.98305, 19.98301, 19.98295, 19.98295, 19.98294, 19.98291, 
    19.98289, 19.98293, 19.98288, 19.98308, 19.98298, 19.98314, 19.98309, 
    19.98306, 19.98307, 19.98299, 19.98298, 19.9829, 19.98294, 19.98271, 
    19.98281, 19.98252, 19.9826, 19.98314, 19.98312, 19.98303, 19.98307, 
    19.98295, 19.98292, 19.9829, 19.98287, 19.98286, 19.98285, 19.98287, 
    19.98285, 19.98295, 19.98291, 19.98304, 19.98301, 19.98302, 19.98304, 
    19.98299, 19.98293, 19.98293, 19.98291, 19.98287, 19.98295, 19.98269, 
    19.98285, 19.98309, 19.98304, 19.98303, 19.98305, 19.98292, 19.98297, 
    19.98285, 19.98288, 19.98282, 19.98285, 19.98285, 19.98289, 19.98291, 
    19.98297, 19.98301, 19.98305, 19.98304, 19.983, 19.98293, 19.98286, 
    19.98288, 19.98283, 19.98296, 19.9829, 19.98293, 19.98287, 19.98299, 
    19.98289, 19.98302, 19.98301, 19.98297, 19.9829, 19.98288, 19.98287, 
    19.98288, 19.98293, 19.98294, 19.98297, 19.98298, 19.98301, 19.98303, 
    19.98301, 19.98299, 19.98293, 19.98287, 19.98281, 19.9828, 19.98273, 
    19.98279, 19.98269, 19.98277, 19.98264, 19.98288, 19.98277, 19.98297, 
    19.98295, 19.98291, 19.98282, 19.98287, 19.98281, 19.98294, 19.983, 
    19.98302, 19.98305, 19.98302, 19.98302, 19.98299, 19.983, 19.98293, 
    19.98296, 19.98285, 19.98281, 19.9827, 19.98264, 19.98256, 19.98253, 
    19.98252, 19.98252,
  19.98426, 19.98419, 19.9842, 19.98414, 19.98418, 19.98414, 19.98424, 
    19.98418, 19.98422, 19.98425, 19.98404, 19.98414, 19.98392, 19.98399, 
    19.98382, 19.98393, 19.9838, 19.98383, 19.98375, 19.98377, 19.98367, 
    19.98374, 19.98362, 19.98368, 19.98368, 19.98374, 19.98412, 19.98405, 
    19.98413, 19.98411, 19.98412, 19.98417, 19.9842, 19.98426, 19.98425, 
    19.98421, 19.98411, 19.98414, 19.98406, 19.98406, 19.98397, 19.98401, 
    19.98385, 19.9839, 19.98377, 19.9838, 19.98377, 19.98378, 19.98377, 
    19.98382, 19.9838, 19.98384, 19.984, 19.98395, 19.9841, 19.98418, 
    19.98424, 19.98428, 19.98428, 19.98426, 19.98421, 19.98416, 19.98412, 
    19.98409, 19.98406, 19.98398, 19.98394, 19.98384, 19.98386, 19.98383, 
    19.9838, 19.98376, 19.98376, 19.98375, 19.98383, 19.98377, 19.98387, 
    19.98384, 19.98405, 19.98413, 19.98417, 19.9842, 19.98427, 19.98422, 
    19.98424, 19.98419, 19.98416, 19.98418, 19.98409, 19.98412, 19.98394, 
    19.98402, 19.98381, 19.98386, 19.9838, 19.98383, 19.98377, 19.98382, 
    19.98374, 19.98372, 19.98373, 19.98368, 19.98382, 19.98377, 19.98418, 
    19.98418, 19.98417, 19.98421, 19.98422, 19.98426, 19.98422, 19.98421, 
    19.98416, 19.98414, 19.98411, 19.98406, 19.984, 19.98391, 19.98385, 
    19.98381, 19.98384, 19.98382, 19.98384, 19.98385, 19.98372, 19.9838, 
    19.98369, 19.9837, 19.98374, 19.9837, 19.98417, 19.98419, 19.98424, 
    19.9842, 19.98427, 19.98423, 19.98421, 19.98412, 19.9841, 19.98409, 
    19.98405, 19.98401, 19.98393, 19.98386, 19.9838, 19.98381, 19.9838, 
    19.98379, 19.98383, 19.98379, 19.98378, 19.9838, 19.9837, 19.98372, 
    19.9837, 19.98372, 19.98418, 19.98416, 19.98417, 19.98415, 19.98417, 
    19.98409, 19.98407, 19.98396, 19.98401, 19.98394, 19.984, 19.98399, 
    19.98394, 19.984, 19.98387, 19.98396, 19.98379, 19.98388, 19.98379, 
    19.9838, 19.98377, 19.98375, 19.98372, 19.98366, 19.98367, 19.98362, 
    19.98413, 19.9841, 19.9841, 19.98407, 19.98404, 19.98399, 19.98391, 
    19.98394, 19.98389, 19.98388, 19.98396, 19.98391, 19.98408, 19.98405, 
    19.98406, 19.98412, 19.98393, 19.98403, 19.98385, 19.98391, 19.98375, 
    19.98383, 19.98368, 19.98362, 19.98356, 19.98349, 19.98408, 19.9841, 
    19.98406, 19.98401, 19.98396, 19.9839, 19.9839, 19.98388, 19.98385, 
    19.98383, 19.98388, 19.98382, 19.98404, 19.98393, 19.98411, 19.98405, 
    19.98401, 19.98403, 19.98395, 19.98392, 19.98384, 19.98388, 19.98363, 
    19.98374, 19.98343, 19.98352, 19.98411, 19.98408, 19.98398, 19.98403, 
    19.9839, 19.98387, 19.98384, 19.98381, 19.9838, 19.98378, 19.98382, 
    19.98378, 19.9839, 19.98385, 19.98399, 19.98396, 19.98397, 19.98399, 
    19.98394, 19.98388, 19.98388, 19.98386, 19.98381, 19.9839, 19.98362, 
    19.98379, 19.98405, 19.984, 19.98399, 19.98401, 19.98387, 19.98392, 
    19.98378, 19.98382, 19.98376, 19.98379, 19.9838, 19.98383, 19.98386, 
    19.98392, 19.98397, 19.984, 19.984, 19.98395, 19.98388, 19.9838, 
    19.98382, 19.98376, 19.98391, 19.98385, 19.98387, 19.98381, 19.98394, 
    19.98383, 19.98397, 19.98396, 19.98392, 19.98384, 19.98383, 19.98381, 
    19.98382, 19.98387, 19.98388, 19.98392, 19.98393, 19.98396, 19.98399, 
    19.98396, 19.98394, 19.98387, 19.98381, 19.98375, 19.98373, 19.98366, 
    19.98372, 19.98362, 19.9837, 19.98355, 19.98382, 19.98371, 19.98392, 
    19.9839, 19.98385, 19.98376, 19.98381, 19.98375, 19.98388, 19.98395, 
    19.98397, 19.984, 19.98397, 19.98397, 19.98394, 19.98395, 19.98387, 
    19.98391, 19.9838, 19.98375, 19.98363, 19.98355, 19.98348, 19.98344, 
    19.98343, 19.98343,
  19.98501, 19.98494, 19.98495, 19.98489, 19.98492, 19.98489, 19.98499, 
    19.98493, 19.98497, 19.985, 19.98478, 19.98489, 19.98467, 19.98474, 
    19.98456, 19.98468, 19.98454, 19.98457, 19.98449, 19.98451, 19.98441, 
    19.98448, 19.98435, 19.98442, 19.98441, 19.98448, 19.98487, 19.98479, 
    19.98487, 19.98486, 19.98487, 19.98492, 19.98495, 19.98501, 19.985, 
    19.98496, 19.98486, 19.98489, 19.9848, 19.98481, 19.98471, 19.98475, 
    19.98459, 19.98464, 19.98451, 19.98454, 19.98451, 19.98452, 19.98451, 
    19.98456, 19.98454, 19.98458, 19.98475, 19.9847, 19.98484, 19.98493, 
    19.98499, 19.98503, 19.98503, 19.98501, 19.98496, 19.9849, 19.98486, 
    19.98483, 19.98481, 19.98473, 19.98468, 19.98458, 19.9846, 19.98457, 
    19.98454, 19.9845, 19.9845, 19.98448, 19.98457, 19.98451, 19.98461, 
    19.98458, 19.9848, 19.98488, 19.98492, 19.98495, 19.98502, 19.98497, 
    19.98499, 19.98494, 19.98491, 19.98493, 19.98483, 19.98487, 19.98468, 
    19.98476, 19.98455, 19.9846, 19.98454, 19.98457, 19.98451, 19.98456, 
    19.98448, 19.98446, 19.98447, 19.98442, 19.98457, 19.98451, 19.98493, 
    19.98492, 19.98491, 19.98496, 19.98497, 19.98501, 19.98497, 19.98495, 
    19.98491, 19.98488, 19.98486, 19.9848, 19.98474, 19.98466, 19.9846, 
    19.98455, 19.98458, 19.98456, 19.98458, 19.98459, 19.98446, 19.98454, 
    19.98443, 19.98443, 19.98448, 19.98443, 19.98492, 19.98494, 19.98499, 
    19.98495, 19.98502, 19.98498, 19.98496, 19.98487, 19.98485, 19.98483, 
    19.9848, 19.98475, 19.98467, 19.98461, 19.98454, 19.98455, 19.98454, 
    19.98453, 19.98457, 19.98453, 19.98452, 19.98454, 19.98443, 19.98446, 
    19.98443, 19.98445, 19.98493, 19.98491, 19.98492, 19.9849, 19.98491, 
    19.98484, 19.98482, 19.98471, 19.98475, 19.98468, 19.98475, 19.98474, 
    19.98468, 19.98474, 19.98461, 19.9847, 19.98453, 19.98462, 19.98453, 
    19.98454, 19.98451, 19.98449, 19.98446, 19.9844, 19.98441, 19.98436, 
    19.98487, 19.98484, 19.98484, 19.98481, 19.98479, 19.98474, 19.98465, 
    19.98469, 19.98463, 19.98462, 19.9847, 19.98465, 19.98482, 19.98479, 
    19.98481, 19.98487, 19.98468, 19.98478, 19.98459, 19.98465, 19.98449, 
    19.98457, 19.98442, 19.98435, 19.98429, 19.98422, 19.98483, 19.98485, 
    19.98481, 19.98476, 19.98471, 19.98464, 19.98464, 19.98463, 19.98459, 
    19.98457, 19.98462, 19.98456, 19.98479, 19.98467, 19.98485, 19.9848, 
    19.98476, 19.98478, 19.98469, 19.98467, 19.98458, 19.98463, 19.98437, 
    19.98448, 19.98417, 19.98425, 19.98485, 19.98483, 19.98473, 19.98477, 
    19.98464, 19.98461, 19.98458, 19.98455, 19.98454, 19.98452, 19.98456, 
    19.98452, 19.98464, 19.98459, 19.98474, 19.9847, 19.98472, 19.98474, 
    19.98468, 19.98462, 19.98462, 19.9846, 19.98455, 19.98464, 19.98435, 
    19.98453, 19.98479, 19.98474, 19.98473, 19.98475, 19.98461, 19.98466, 
    19.98452, 19.98456, 19.9845, 19.98453, 19.98454, 19.98457, 19.9846, 
    19.98466, 19.98471, 19.98475, 19.98474, 19.9847, 19.98462, 19.98454, 
    19.98456, 19.9845, 19.98465, 19.98459, 19.98461, 19.98455, 19.98469, 
    19.98457, 19.98472, 19.9847, 19.98466, 19.98458, 19.98457, 19.98455, 
    19.98456, 19.98462, 19.98462, 19.98466, 19.98468, 19.9847, 19.98473, 
    19.98471, 19.98468, 19.98462, 19.98455, 19.98449, 19.98447, 19.98439, 
    19.98446, 19.98435, 19.98444, 19.98429, 19.98456, 19.98444, 19.98466, 
    19.98464, 19.9846, 19.9845, 19.98455, 19.98449, 19.98462, 19.9847, 
    19.98471, 19.98475, 19.98471, 19.98472, 19.98468, 19.98469, 19.98461, 
    19.98466, 19.98454, 19.98449, 19.98436, 19.98429, 19.98421, 19.98417, 
    19.98416, 19.98416,
  19.98609, 19.98602, 19.98603, 19.98598, 19.98601, 19.98598, 19.98607, 
    19.98602, 19.98605, 19.98608, 19.98588, 19.98598, 19.98577, 19.98584, 
    19.98568, 19.98579, 19.98566, 19.98568, 19.98561, 19.98563, 19.98554, 
    19.9856, 19.98549, 19.98555, 19.98554, 19.9856, 19.98596, 19.98589, 
    19.98596, 19.98595, 19.98596, 19.98601, 19.98603, 19.98609, 19.98608, 
    19.98604, 19.98595, 19.98598, 19.9859, 19.9859, 19.98582, 19.98586, 
    19.98571, 19.98575, 19.98563, 19.98566, 19.98563, 19.98564, 19.98563, 
    19.98568, 19.98566, 19.98569, 19.98585, 19.9858, 19.98594, 19.98602, 
    19.98607, 19.98611, 19.9861, 19.98609, 19.98604, 19.98599, 19.98595, 
    19.98593, 19.9859, 19.98583, 19.98579, 19.9857, 19.98572, 19.98569, 
    19.98566, 19.98562, 19.98563, 19.98561, 19.98569, 19.98564, 19.98573, 
    19.9857, 19.9859, 19.98597, 19.986, 19.98603, 19.9861, 19.98605, 
    19.98607, 19.98603, 19.986, 19.98601, 19.98593, 19.98596, 19.98579, 
    19.98586, 19.98567, 19.98571, 19.98565, 19.98568, 19.98563, 19.98568, 
    19.9856, 19.98558, 19.98559, 19.98555, 19.98568, 19.98563, 19.98601, 
    19.98601, 19.986, 19.98605, 19.98605, 19.98609, 19.98605, 19.98604, 
    19.986, 19.98597, 19.98595, 19.9859, 19.98584, 19.98577, 19.98571, 
    19.98567, 19.98569, 19.98567, 19.9857, 19.98571, 19.98559, 19.98566, 
    19.98556, 19.98556, 19.98561, 19.98556, 19.98601, 19.98602, 19.98607, 
    19.98603, 19.9861, 19.98606, 19.98604, 19.98596, 19.98594, 19.98593, 
    19.98589, 19.98585, 19.98578, 19.98572, 19.98566, 19.98567, 19.98566, 
    19.98565, 19.98568, 19.98565, 19.98564, 19.98566, 19.98556, 19.98559, 
    19.98556, 19.98558, 19.98602, 19.986, 19.98601, 19.98598, 19.986, 
    19.98593, 19.98591, 19.98581, 19.98585, 19.98579, 19.98585, 19.98584, 
    19.98579, 19.98584, 19.98572, 19.98581, 19.98565, 19.98573, 19.98565, 
    19.98566, 19.98564, 19.98561, 19.98558, 19.98553, 19.98554, 19.98549, 
    19.98596, 19.98594, 19.98594, 19.98591, 19.98589, 19.98584, 19.98576, 
    19.98579, 19.98574, 19.98573, 19.98581, 19.98576, 19.98592, 19.98589, 
    19.98591, 19.98596, 19.98578, 19.98588, 19.98571, 19.98576, 19.98561, 
    19.98569, 19.98555, 19.98549, 19.98543, 19.98536, 19.98592, 19.98594, 
    19.9859, 19.98586, 19.98581, 19.98575, 19.98575, 19.98574, 19.98571, 
    19.98569, 19.98573, 19.98568, 19.98589, 19.98578, 19.98595, 19.9859, 
    19.98586, 19.98588, 19.9858, 19.98578, 19.9857, 19.98574, 19.9855, 
    19.98561, 19.98531, 19.9854, 19.98594, 19.98592, 19.98583, 19.98587, 
    19.98575, 19.98572, 19.9857, 19.98566, 19.98566, 19.98564, 19.98567, 
    19.98564, 19.98575, 19.9857, 19.98584, 19.98581, 19.98582, 19.98584, 
    19.98579, 19.98573, 19.98573, 19.98571, 19.98567, 19.98575, 19.98549, 
    19.98565, 19.98589, 19.98584, 19.98583, 19.98586, 19.98572, 19.98577, 
    19.98564, 19.98568, 19.98562, 19.98565, 19.98565, 19.98569, 19.98571, 
    19.98577, 19.98582, 19.98585, 19.98584, 19.9858, 19.98573, 19.98566, 
    19.98568, 19.98563, 19.98576, 19.9857, 19.98573, 19.98567, 19.98579, 
    19.98569, 19.98582, 19.98581, 19.98577, 19.9857, 19.98568, 19.98567, 
    19.98568, 19.98573, 19.98574, 19.98577, 19.98578, 19.98581, 19.98583, 
    19.98581, 19.98579, 19.98573, 19.98567, 19.98561, 19.9856, 19.98553, 
    19.98558, 19.98549, 19.98557, 19.98543, 19.98568, 19.98557, 19.98577, 
    19.98575, 19.98571, 19.98562, 19.98567, 19.98561, 19.98574, 19.9858, 
    19.98582, 19.98585, 19.98582, 19.98582, 19.98579, 19.9858, 19.98573, 
    19.98577, 19.98565, 19.98561, 19.9855, 19.98543, 19.98536, 19.98532, 
    19.98531, 19.98531,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.72228, 0.7222776, 0.7222781, 0.7222761, 0.7222772, 0.7222759, 0.7222795, 
    0.7222775, 0.7222788, 0.7222798, 0.7222724, 0.722276, 0.7222686, 
    0.7222709, 0.722265, 0.7222689, 0.7222642, 0.7222651, 0.7222624, 
    0.7222632, 0.7222598, 0.7222621, 0.722258, 0.7222603, 0.7222599, 
    0.7222621, 0.7222753, 0.7222728, 0.7222754, 0.7222751, 0.7222753, 
    0.7222772, 0.7222781, 0.7222801, 0.7222798, 0.7222783, 0.722275, 
    0.7222761, 0.7222732, 0.7222732, 0.72227, 0.7222715, 0.7222661, 
    0.7222676, 0.7222632, 0.7222643, 0.7222632, 0.7222635, 0.7222632, 
    0.7222648, 0.7222642, 0.7222656, 0.7222712, 0.7222695, 0.7222745, 
    0.7222775, 0.7222794, 0.7222808, 0.7222806, 0.7222803, 0.7222783, 
    0.7222765, 0.7222751, 0.7222742, 0.7222733, 0.7222705, 0.7222691, 
    0.7222658, 0.7222664, 0.7222654, 0.7222644, 0.7222628, 0.722263, 
    0.7222623, 0.7222654, 0.7222633, 0.7222667, 0.7222658, 0.722273, 
    0.7222758, 0.7222769, 0.7222779, 0.7222804, 0.7222787, 0.7222794, 
    0.7222778, 0.7222767, 0.7222773, 0.7222741, 0.7222754, 0.7222689, 
    0.7222717, 0.7222645, 0.7222663, 0.7222641, 0.7222652, 0.7222633, 
    0.722265, 0.7222621, 0.7222614, 0.7222619, 0.7222602, 0.7222651, 
    0.7222632, 0.7222773, 0.7222772, 0.7222768, 0.7222785, 0.7222787, 
    0.7222802, 0.7222788, 0.7222782, 0.7222767, 0.7222759, 0.722275, 
    0.7222732, 0.7222711, 0.7222682, 0.7222661, 0.7222647, 0.7222656, 
    0.7222648, 0.7222657, 0.7222661, 0.7222617, 0.7222642, 0.7222605, 
    0.7222607, 0.7222623, 0.7222607, 0.7222772, 0.7222776, 0.7222793, 
    0.722278, 0.7222803, 0.722279, 0.7222783, 0.7222753, 0.7222747, 
    0.7222741, 0.7222729, 0.7222714, 0.7222688, 0.7222664, 0.7222643, 
    0.7222645, 0.7222645, 0.722264, 0.7222651, 0.7222638, 0.7222636, 
    0.7222642, 0.7222607, 0.7222617, 0.7222607, 0.7222613, 0.7222775, 
    0.7222767, 0.7222771, 0.7222763, 0.7222769, 0.7222743, 0.7222735, 
    0.72227, 0.7222714, 0.7222691, 0.7222712, 0.7222708, 0.722269, 0.7222711, 
    0.7222666, 0.7222697, 0.7222639, 0.722267, 0.7222638, 0.7222643, 
    0.7222634, 0.7222625, 0.7222614, 0.7222593, 0.7222598, 0.7222582, 
    0.7222755, 0.7222744, 0.7222745, 0.7222735, 0.7222726, 0.7222709, 
    0.7222681, 0.7222692, 0.7222672, 0.7222669, 0.7222698, 0.722268, 
    0.7222738, 0.7222728, 0.7222733, 0.7222754, 0.7222689, 0.7222722, 
    0.7222661, 0.7222679, 0.7222626, 0.7222652, 0.7222601, 0.7222579, 
    0.7222558, 0.7222534, 0.7222739, 0.7222746, 0.7222733, 0.7222716, 
    0.72227, 0.7222678, 0.7222676, 0.7222672, 0.7222661, 0.7222652, 0.722267, 
    0.722265, 0.7222726, 0.7222686, 0.7222748, 0.722273, 0.7222717, 
    0.7222722, 0.7222693, 0.7222686, 0.7222657, 0.7222672, 0.7222584, 
    0.7222623, 0.7222516, 0.7222546, 0.7222748, 0.7222739, 0.7222705, 
    0.7222722, 0.7222676, 0.7222666, 0.7222656, 0.7222645, 0.7222643, 
    0.7222637, 0.7222648, 0.7222637, 0.7222677, 0.722266, 0.722271, 
    0.7222697, 0.7222703, 0.7222709, 0.722269, 0.722267, 0.722267, 0.7222663, 
    0.7222645, 0.7222676, 0.7222579, 0.7222639, 0.7222728, 0.722271, 
    0.7222707, 0.7222714, 0.7222666, 0.7222684, 0.7222637, 0.7222649, 
    0.7222629, 0.7222639, 0.7222641, 0.7222654, 0.7222662, 0.7222683, 
    0.72227, 0.7222713, 0.722271, 0.7222695, 0.7222669, 0.7222643, 0.7222649, 
    0.722263, 0.722268, 0.7222659, 0.7222667, 0.7222646, 0.7222692, 
    0.7222653, 0.7222702, 0.7222697, 0.7222684, 0.7222658, 0.7222652, 
    0.7222645, 0.7222649, 0.7222668, 0.7222671, 0.7222685, 0.7222688, 
    0.7222698, 0.7222707, 0.7222699, 0.7222691, 0.7222668, 0.7222648, 
    0.7222625, 0.7222619, 0.7222593, 0.7222614, 0.7222579, 0.7222609, 
    0.7222557, 0.7222651, 0.722261, 0.7222683, 0.7222676, 0.7222661, 
    0.7222629, 0.7222646, 0.7222626, 0.7222672, 0.7222695, 0.7222701, 
    0.7222713, 0.7222701, 0.7222702, 0.7222691, 0.7222694, 0.7222667, 
    0.7222682, 0.7222641, 0.7222626, 0.7222583, 0.7222557, 0.7222531, 
    0.7222519, 0.7222515, 0.7222514 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  2.055969e-20, -2.055969e-20, -1.541976e-20, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 2.055969e-20, 3.083953e-20, -5.139921e-21, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, -2.055969e-20, -1.541976e-20, 
    1.541976e-20, 1.027984e-20, 0, 1.541976e-20, 4.111937e-20, -5.139921e-21, 
    -5.139921e-21, 2.055969e-20, 1.541976e-20, 1.541976e-20, 2.006177e-36, 
    -1.027984e-20, -1.541976e-20, 3.083953e-20, 2.055969e-20, 2.055969e-20, 
    -5.139921e-21, -3.083953e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    2.006177e-36, -1.027984e-20, -4.625929e-20, 2.055969e-20, 2.569961e-20, 
    0, -5.139921e-21, 3.597945e-20, -2.055969e-20, 0, -5.139921e-20, 
    -2.055969e-20, -2.055969e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    0, 5.139921e-21, -4.111937e-20, -1.541976e-20, -3.597945e-20, 
    -3.083953e-20, -5.139921e-21, 2.569961e-20, -2.569961e-20, -2.569961e-20, 
    -1.027984e-20, -1.541976e-20, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    -5.653913e-20, -1.027984e-20, -1.027984e-20, 5.139921e-21, 2.569961e-20, 
    2.569961e-20, 2.055969e-20, -5.139921e-21, 2.569961e-20, 5.139921e-21, 
    3.083953e-20, -5.139921e-21, -5.139921e-21, 2.006177e-36, -2.055969e-20, 
    5.139921e-21, -3.597945e-20, -5.139921e-21, 2.055969e-20, 5.139921e-21, 
    3.597945e-20, 3.597945e-20, -3.083953e-20, 1.541976e-20, -1.027984e-20, 
    1.541976e-20, -1.541976e-20, 2.006177e-36, -1.027984e-20, -2.569961e-20, 
    -5.139921e-21, 0, 4.625929e-20, 1.541976e-20, -1.027984e-20, 
    -1.027984e-20, 1.541976e-20, -5.139921e-21, -2.055969e-20, 2.055969e-20, 
    5.139921e-21, 2.055969e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, 0, 
    0, -1.027984e-20, 2.055969e-20, -2.569961e-20, 0, -1.027984e-20, 
    -2.006177e-36, 2.055969e-20, -5.139921e-21, -2.055969e-20, -2.055969e-20, 
    1.027984e-20, -5.139921e-21, 2.055969e-20, 2.055969e-20, -5.139921e-21, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -2.569961e-20, 1.541976e-20, 
    1.541976e-20, -1.541976e-20, 5.139921e-21, 0, -3.083953e-20, 
    -5.139921e-21, 2.006177e-36, -1.541976e-20, 4.111937e-20, 1.541976e-20, 
    5.139921e-21, -3.083953e-20, 1.541976e-20, -2.569961e-20, -1.027984e-20, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 1.541976e-20, 3.597945e-20, 
    -5.139921e-21, -1.027984e-20, 1.541976e-20, 3.083953e-20, 2.006177e-36, 
    0, 1.541976e-20, -1.027984e-20, 0, -2.569961e-20, 2.569961e-20, 
    2.006177e-36, 0, -3.083953e-20, -1.541976e-20, 0, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, 
    2.006177e-36, -2.569961e-20, -1.027984e-20, 2.055969e-20, 0, 
    2.055969e-20, 1.541976e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 2.569961e-20, 2.569961e-20, 2.569961e-20, 3.083953e-20, 
    -2.006177e-36, 1.027984e-20, 2.055969e-20, 1.541976e-20, 2.006177e-36, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, 3.083953e-20, -2.055969e-20, 
    2.569961e-20, -1.541976e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 2.055969e-20, 
    -1.027984e-20, -5.139921e-21, 0, 0, -2.569961e-20, -5.653913e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, -2.569961e-20, 
    5.139921e-21, 4.111937e-20, 1.541976e-20, -2.055969e-20, 5.139921e-21, 
    1.027984e-20, 2.055969e-20, 2.055969e-20, -2.569961e-20, 0, 2.055969e-20, 
    4.111937e-20, 1.541976e-20, -5.139921e-21, 2.055969e-20, -1.541976e-20, 
    1.541976e-20, 1.541976e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -2.055969e-20, -2.569961e-20, 1.541976e-20, 2.055969e-20, 2.055969e-20, 
    -1.541976e-20, -5.139921e-21, -2.006177e-36, 5.139921e-21, 0, 
    2.569961e-20, 2.569961e-20, 2.006177e-36, -3.597945e-20, 5.139921e-21, 
    -4.111937e-20, 0, 1.027984e-20, 0, -2.055969e-20, 2.055969e-20, 
    3.597945e-20, 0, -5.139921e-21, -5.139921e-21, 2.569961e-20, 
    -1.027984e-20, -1.541976e-20, 2.569961e-20, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -2.055969e-20, 3.597945e-20, 1.541976e-20, 5.139921e-21, 4.625929e-20, 
    -2.006177e-36, 2.006177e-36, -1.027984e-20, -3.597945e-20, 3.083953e-20, 
    -2.055969e-20, -2.055969e-20, -2.006177e-36, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, -1.027984e-20, -3.597945e-20, -2.569961e-20, 3.083953e-20, 
    1.541976e-20, -5.139921e-21, 2.569961e-20, 2.569961e-20, 5.139921e-21, 
    -2.006177e-36, -5.139921e-21, 1.541976e-20, 0, 2.055969e-20, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, 1.541976e-20, 2.569961e-20, 
    1.541976e-20, 2.055969e-20, 5.139921e-21, -2.006177e-36, -1.541976e-20, 
    1.541976e-20, -3.597945e-20, 2.569961e-20, 5.139921e-21, -2.006177e-36, 
    1.541976e-20, -3.083953e-20, -5.139921e-21, -2.055969e-20, 2.569961e-20, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 3.597945e-20, 
    0, 5.139921e-21, -5.139921e-21, -5.139921e-21,
  2.055969e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 2.055969e-20, 
    1.027984e-20, 0, -1.027984e-20, -2.569961e-20, -1.027984e-20, 0, 
    3.083953e-20, -1.541976e-20, 2.055969e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, -3.083953e-20, 
    5.139921e-21, -4.111937e-20, 5.139921e-21, 1.027984e-20, 2.055969e-20, 
    2.055969e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 0, 
    -2.569961e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, -2.006177e-36, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.055969e-20, 
    -1.027984e-20, 0, -2.569961e-20, -5.139921e-21, -1.027984e-20, 0, 
    2.006177e-36, 2.006177e-36, -4.111937e-20, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 2.006177e-36, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, -2.569961e-20, 
    -5.139921e-21, -4.111937e-20, 1.541976e-20, 2.006177e-36, -1.541976e-20, 
    -2.055969e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    2.006177e-36, 5.139921e-21, 2.569961e-20, -3.083953e-20, -2.055969e-20, 
    -2.569961e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 3.083953e-20, 
    2.569961e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -2.006177e-36, 3.083953e-20, 5.139921e-21, -2.006177e-36, 1.541976e-20, 
    -2.055969e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -2.055969e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 1.027984e-20, 5.139921e-20, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, 3.083953e-20, -1.541976e-20, 0, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, 2.569961e-20, 5.139921e-21, 
    -3.597945e-20, 0, 1.027984e-20, -1.027984e-20, 4.111937e-20, 
    -2.055969e-20, 1.541976e-20, 1.541976e-20, -1.027984e-20, 0, 
    -1.027984e-20, 0, -1.541976e-20, -1.541976e-20, 0, -3.083953e-20, 
    5.139921e-21, -1.541976e-20, 1.541976e-20, -1.027984e-20, 2.055969e-20, 
    5.139921e-21, 0, -5.139921e-21, -2.569961e-20, 2.055969e-20, 
    1.027984e-20, 2.006177e-36, 2.055969e-20, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, -2.055969e-20, 5.139921e-21, 1.541976e-20, 
    2.569961e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 0, 1.541976e-20, 
    0, -2.569961e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, -1.027984e-20, 4.625929e-20, -1.027984e-20, 0, 
    -5.139921e-21, -2.055969e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    -2.006177e-36, -5.139921e-21, 1.541976e-20, -1.027984e-20, 5.139921e-21, 
    -4.111937e-20, 5.139921e-21, 1.027984e-20, 2.055969e-20, 2.055969e-20, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, 0, -1.541976e-20, 
    -2.055969e-20, -2.055969e-20, 5.139921e-21, 0, -4.625929e-20, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, 0, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 0, 
    2.569961e-20, 1.541976e-20, -5.139921e-21, -2.055969e-20, -1.027984e-20, 
    1.027984e-20, 2.569961e-20, 2.055969e-20, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, -2.569961e-20, -1.027984e-20, 0, -2.569961e-20, 
    2.055969e-20, -5.139921e-21, -1.027984e-20, 0, -5.139921e-21, 
    1.541976e-20, 0, 1.541976e-20, 0, 0, 0, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 2.055969e-20, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -3.597945e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 0, 
    5.139921e-21, 5.139921e-21, 0, 1.541976e-20, -2.055969e-20, 
    -2.569961e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-20, 5.139921e-20, 2.055969e-20, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 0, 5.139921e-21, -2.569961e-20, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, -1.541976e-20, -3.597945e-20, -1.541976e-20, 0, 
    1.027984e-20, 5.139921e-21, -2.055969e-20, 2.006177e-36, -1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 0, 1.027984e-20, 1.027984e-20, 
    -2.569961e-20, 0, 1.027984e-20, 1.027984e-20, 0, 0, 2.569961e-20, 
    -1.027984e-20, 2.055969e-20, -2.569961e-20, -1.027984e-20, 0, 
    5.139921e-21, 0, -5.139921e-21, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, -3.083953e-20, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, -4.111937e-20, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, -2.055969e-20, 1.027984e-20, -1.541976e-20, 
    -1.541976e-20, 3.083953e-20, 0, 0, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -2.055969e-20, 1.027984e-20,
  2.006177e-36, -2.569961e-20, 1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -2.569961e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, 3.597945e-20, 
    5.139921e-21, 0, 5.139921e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-20, 2.006177e-36, 1.027984e-20, 
    4.111937e-20, -2.569961e-20, -5.139921e-21, -2.055969e-20, 0, 
    3.597945e-20, 0, 0, 1.541976e-20, 0, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, 5.139921e-21, 0, -2.055969e-20, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, -3.083953e-20, 5.139921e-21, 
    -2.569961e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, 1.027984e-20, 
    5.139921e-21, 0, 1.027984e-20, 4.111937e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 3.083953e-20, 5.139921e-21, 2.569961e-20, 0, 
    -1.027984e-20, 1.541976e-20, -1.027984e-20, 2.055969e-20, -2.569961e-20, 
    -1.027984e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -3.083953e-20, 5.139921e-21, -1.541976e-20, 4.625929e-20, 
    0, 5.139921e-20, 5.139921e-21, 2.006177e-36, -1.027984e-20, 
    -2.055969e-20, -2.006177e-36, 2.569961e-20, -1.541976e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, -2.006177e-36, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -1.541976e-20, 2.569961e-20, -2.569961e-20, 
    1.027984e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, 0, 1.541976e-20, -5.139921e-21, 2.006177e-36, 
    -5.139921e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    2.006177e-36, 1.027984e-20, 2.569961e-20, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, -1.027984e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -2.055969e-20, -2.006177e-36, 3.083953e-20, 0, 
    1.027984e-20, 2.006177e-36, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -3.083953e-20, 0, 
    -5.139921e-21, 5.139921e-21, -2.006177e-36, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 2.055969e-20, 2.055969e-20, -1.541976e-20, 2.055969e-20, 
    2.006177e-36, 5.139921e-21, 1.027984e-20, 2.055969e-20, 3.083953e-20, 
    2.006177e-36, -5.139921e-21, -1.027984e-20, 1.541976e-20, 1.541976e-20, 
    2.055969e-20, 2.055969e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, 
    0, 5.139921e-21, -3.597945e-20, 5.139921e-21, -5.139921e-21, 
    2.055969e-20, -2.569961e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, -1.541976e-20, -1.541976e-20, 
    5.139921e-21, 1.027984e-20, 2.055969e-20, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 0, 1.027984e-20, -1.027984e-20, 2.006177e-36, 
    -5.139921e-21, -2.055969e-20, -2.006177e-36, 1.541976e-20, 0, 
    -5.139921e-21, 2.006177e-36, 5.139921e-21, -1.541976e-20, -4.111937e-20, 
    5.139921e-21, 2.055969e-20, 2.055969e-20, -3.597945e-20, -5.139921e-21, 
    2.055969e-20, -1.541976e-20, -2.006177e-36, 0, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, -3.597945e-20, 1.541976e-20, 
    3.083953e-20, 1.027984e-20, 5.139921e-21, 4.625929e-20, 4.111937e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, 3.083953e-20, 0, 0, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, 3.597945e-20, 2.055969e-20, 
    2.055969e-20, -2.569961e-20, -2.569961e-20, -2.006177e-36, 5.139921e-21, 
    -3.083953e-20, 2.569961e-20, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, -5.139921e-21, 
    0, 0, -5.139921e-21, 2.055969e-20, 2.569961e-20, 2.055969e-20, 
    5.139921e-21, -5.139921e-21, 0, -1.027984e-20, 0, -3.597945e-20, 
    -5.139921e-21, 1.541976e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, 3.597945e-20, 1.027984e-20, 0, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, -2.006177e-36, 
    -5.139921e-21, 2.055969e-20, 0, 5.139921e-21, -7.709882e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, -2.569961e-20, -2.055969e-20, 
    1.541976e-20, 0, 4.111937e-20, 5.139921e-21, 2.006177e-36, 0, 
    -1.541976e-20, -3.083953e-20, -1.027984e-20, -2.569961e-20, 
    -2.006177e-36, -1.027984e-20, -2.055969e-20, 1.541976e-20, 2.006177e-36, 
    3.083953e-20, -3.083953e-20, 0, -5.139921e-21, -1.541976e-20, 
    -2.006177e-36, 2.055969e-20, 2.006177e-36, 2.055969e-20, -1.027984e-20, 
    -1.541976e-20, 4.625929e-20, -1.541976e-20, 2.006177e-36, 2.055969e-20, 
    -5.139921e-21, 2.006177e-36, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, 2.055969e-20, -2.055969e-20, -5.139921e-21, -2.006177e-36, 
    5.139921e-21,
  -5.139921e-21, 2.569961e-20, 5.139921e-21, 1.541976e-20, 2.055969e-20, 
    -5.139921e-21, 2.569961e-20, -2.569961e-20, -2.055969e-20, -2.006177e-36, 
    1.541976e-20, 0, 2.055969e-20, 1.541976e-20, 1.541976e-20, -2.055969e-20, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 3.597945e-20, 
    -1.541976e-20, 0, 1.027984e-20, 3.597945e-20, 1.027984e-20, 
    -3.597945e-20, 5.139921e-21, -5.139921e-21, 0, -2.569961e-20, 
    1.027984e-20, -2.569961e-20, -3.083953e-20, -5.139921e-21, -1.541976e-20, 
    -1.541976e-20, 1.541976e-20, 0, -2.569961e-20, 1.541976e-20, 
    -2.006177e-36, 2.569961e-20, -1.541976e-20, -1.541976e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, -2.055969e-20, 3.083953e-20, -2.006177e-36, 
    2.006177e-36, -2.055969e-20, 1.027984e-20, 2.006177e-36, 4.111937e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -2.569961e-20, 2.055969e-20, -1.027984e-20, 5.139921e-21, -2.569961e-20, 
    -1.027984e-20, 2.569961e-20, 2.569961e-20, -5.139921e-21, -2.006177e-36, 
    1.541976e-20, -2.006177e-36, -2.569961e-20, 2.569961e-20, 3.083953e-20, 
    2.569961e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 0, 3.083953e-20, 
    1.541976e-20, -2.055969e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    4.625929e-20, 0, -4.111937e-20, 5.139921e-21, -3.083953e-20, 
    -1.027984e-20, 1.027984e-20, -2.055969e-20, -5.139921e-21, -2.006177e-36, 
    5.139921e-21, 2.006177e-36, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    3.083953e-20, 0, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, -1.027984e-20, 0, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, 5.139921e-21, -2.569961e-20, 
    1.027984e-20, -2.055969e-20, 0, -1.027984e-20, -2.055969e-20, 
    -1.541976e-20, -3.597945e-20, 3.597945e-20, -1.541976e-20, 0, 
    2.569961e-20, -2.055969e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, 0, 1.027984e-20, -1.541976e-20, 0, -1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 3.083953e-20, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, -3.597945e-20, 3.083953e-20, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -2.569961e-20, -5.139921e-21, 
    -3.083953e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    2.055969e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, -5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -3.083953e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    4.111937e-20, -5.139921e-21, -1.027984e-20, 2.055969e-20, 2.569961e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 4.111937e-20, 2.055969e-20, 
    2.006177e-36, 2.055969e-20, 2.055969e-20, -1.027984e-20, 0, 1.541976e-20, 
    -2.569961e-20, -5.139921e-21, 0, 1.541976e-20, 4.111937e-20, 
    -2.006177e-36, 5.139921e-21, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -3.597945e-20, -2.006177e-36, -5.139921e-21, -2.006177e-36, 2.055969e-20, 
    1.541976e-20, -1.027984e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 
    2.569961e-20, 2.569961e-20, 1.541976e-20, -1.027984e-20, -2.055969e-20, 
    -1.541976e-20, 1.027984e-20, 1.027984e-20, 4.111937e-20, 3.083953e-20, 
    -2.055969e-20, -3.597945e-20, 3.083953e-20, -1.027984e-20, 1.541976e-20, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, -2.055969e-20, 2.569961e-20, 
    0, -5.139921e-21, -2.055969e-20, -5.139921e-21, 3.597945e-20, 
    -1.027984e-20, 0, -1.027984e-20, -5.139921e-21, -4.625929e-20, 
    3.597945e-20, 5.139921e-21, -1.541976e-20, 2.569961e-20, 5.139921e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, -4.625929e-20, 
    -4.625929e-20, 2.569961e-20, 1.027984e-20, 5.139921e-21, 0, 1.541976e-20, 
    -1.541976e-20, -1.541976e-20, 2.569961e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 1.541976e-20, 5.139921e-21, -1.541976e-20, 1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, 2.055969e-20, -1.541976e-20, 
    0, 2.569961e-20, 2.569961e-20, 0, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 0, -1.541976e-20, 
    -2.055969e-20, 1.541976e-20, -1.027984e-20, 1.541976e-20, -1.541976e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, -3.083953e-20, 
    2.569961e-20, 5.139921e-21, 3.083953e-20, -1.541976e-20, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.055969e-20, 1.541976e-20, 3.083953e-20, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, -1.541976e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    3.083953e-20, -5.139921e-21, 1.541976e-20, -2.055969e-20, 1.541976e-20, 
    1.027984e-20, 1.027984e-20, 5.139921e-21, -3.597945e-20, 3.083953e-20, 
    -1.027984e-20, 2.569961e-20, -1.541976e-20, -3.083953e-20,
  -1.541976e-20, 3.597945e-20, 1.541976e-20, 2.569961e-20, 1.541976e-20, 
    -3.083953e-20, 5.139921e-21, 1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, 2.055969e-20, 5.139921e-21, 
    1.541976e-20, -2.055969e-20, 5.139921e-21, -1.541976e-20, 0, 
    -2.055969e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, -4.111937e-20, 1.027984e-20, 3.083953e-20, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, -5.139921e-21, -2.006177e-36, 
    2.055969e-20, -5.139921e-21, -2.055969e-20, 2.006177e-36, -2.055969e-20, 
    -1.027984e-20, 2.006177e-36, -1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -2.055969e-20, 0, 1.541976e-20, -1.541976e-20, 1.027984e-20, 0, 
    3.083953e-20, 2.055969e-20, 3.083953e-20, 1.027984e-20, 0, -2.055969e-20, 
    -5.139921e-21, -1.027984e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    -2.055969e-20, -2.006177e-36, 2.055969e-20, 2.055969e-20, -1.027984e-20, 
    2.055969e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.055969e-20, 
    2.569961e-20, 1.027984e-20, 0, 1.027984e-20, 0, 2.055969e-20, 0, 
    5.139921e-21, -5.139921e-21, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    2.055969e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 2.055969e-20, 5.139921e-21, -3.083953e-20, 
    -1.541976e-20, 3.597945e-20, -3.597945e-20, -5.139921e-21, -4.111937e-20, 
    1.027984e-20, -2.055969e-20, 0, -2.569961e-20, -3.083953e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 2.055969e-20, 1.027984e-20, 
    1.027984e-20, -2.055969e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, -5.139921e-20, 2.569961e-20, -2.006177e-36, -2.055969e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 2.055969e-20, 
    5.139921e-21, -2.055969e-20, -2.569961e-20, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, -3.597945e-20, 2.055969e-20, -4.111937e-20, -5.139921e-21, 
    3.083953e-20, 2.569961e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -1.541976e-20, 1.541976e-20, -1.541976e-20, 2.569961e-20, 0, 
    -5.139921e-21, -2.569961e-20, -3.083953e-20, -5.139921e-21, 1.541976e-20, 
    2.055969e-20, 0, -1.027984e-20, 3.083953e-20, -2.006177e-36, 
    2.055969e-20, 1.541976e-20, 1.027984e-20, 2.006177e-36, -5.139921e-21, 
    -2.569961e-20, -5.139921e-21, 5.139921e-21, 0, 1.027984e-20, 
    -4.111937e-20, -1.027984e-20, 2.569961e-20, -1.027984e-20, 1.027984e-20, 
    -3.083953e-20, -3.083953e-20, 1.541976e-20, 2.569961e-20, -2.055969e-20, 
    2.006177e-36, 1.027984e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, 0, -2.569961e-20, 
    1.541976e-20, 5.139921e-21, 4.111937e-20, 2.055969e-20, 1.541976e-20, 0, 
    0, 0, -5.139921e-21, 1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, 0, -1.027984e-20, 
    5.139921e-21, 2.006177e-36, 1.027984e-20, 0, 0, 2.055969e-20, 
    4.625929e-20, 1.027984e-20, -2.055969e-20, 2.569961e-20, -5.139921e-21, 
    -1.027984e-20, 0, -1.027984e-20, 3.597945e-20, 3.083953e-20, 
    -2.006177e-36, 0, 5.139921e-21, 5.139921e-21, -2.055969e-20, 
    -3.597945e-20, -1.541976e-20, 2.055969e-20, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -2.055969e-20, 2.055969e-20, -3.083953e-20, 2.569961e-20, 
    -1.541976e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    5.139921e-21, 5.139921e-21, -2.055969e-20, 2.569961e-20, -1.027984e-20, 
    -5.139921e-21, 0, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    2.055969e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, 
    1.027984e-20, 5.139921e-21, 0, -5.139921e-21, 2.055969e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, -4.625929e-20, -5.139921e-21, -2.055969e-20, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, 0, -1.541976e-20, 
    -5.139921e-21, -2.055969e-20, -1.027984e-20, 1.027984e-20, -2.055969e-20, 
    3.083953e-20, 5.139921e-21, -2.569961e-20, -1.541976e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, 4.111937e-20, 2.055969e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -3.597945e-20, -2.569961e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -2.569961e-20, 1.541976e-20, 
    5.139921e-21, 2.006177e-36, -1.027984e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 0, 2.006177e-36, 2.055969e-20, 
    -1.541976e-20, -3.083953e-20, 3.083953e-20, 0, 1.027984e-20, 
    3.083953e-20, -2.055969e-20, 0, 2.055969e-20, 1.027984e-20, 0, 
    -2.569961e-20, 3.083953e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 3.083953e-20, -5.139921e-21, 3.083953e-20, 4.111937e-20, 
    2.006177e-36, 5.139921e-21, -5.139921e-21, -2.569961e-20, 5.139921e-21, 
    -2.055969e-20, -2.055969e-20, 0, 1.027984e-20, -2.006177e-36, 
    5.139921e-21, 3.083953e-20, 0, 2.569961e-20,
  8.598827e-29, 8.598799e-29, 8.598805e-29, 8.598782e-29, 8.598795e-29, 
    8.598779e-29, 8.598822e-29, 8.598798e-29, 8.598813e-29, 8.598825e-29, 
    8.598739e-29, 8.598781e-29, 8.598694e-29, 8.598721e-29, 8.598652e-29, 
    8.598698e-29, 8.598643e-29, 8.598654e-29, 8.598622e-29, 8.598631e-29, 
    8.598591e-29, 8.598618e-29, 8.59857e-29, 8.598597e-29, 8.598593e-29, 
    8.598619e-29, 8.598772e-29, 8.598743e-29, 8.598774e-29, 8.59877e-29, 
    8.598772e-29, 8.598794e-29, 8.598805e-29, 8.598829e-29, 8.598825e-29, 
    8.598808e-29, 8.598768e-29, 8.598781e-29, 8.598748e-29, 8.598749e-29, 
    8.598711e-29, 8.598728e-29, 8.598665e-29, 8.598683e-29, 8.598631e-29, 
    8.598644e-29, 8.598631e-29, 8.598635e-29, 8.598631e-29, 8.598651e-29, 
    8.598642e-29, 8.598659e-29, 8.598725e-29, 8.598705e-29, 8.598763e-29, 
    8.598798e-29, 8.59882e-29, 8.598837e-29, 8.598834e-29, 8.59883e-29, 
    8.598807e-29, 8.598786e-29, 8.59877e-29, 8.59876e-29, 8.598749e-29, 
    8.598716e-29, 8.598699e-29, 8.598662e-29, 8.598668e-29, 8.598657e-29, 
    8.598645e-29, 8.598627e-29, 8.59863e-29, 8.598621e-29, 8.598657e-29, 
    8.598633e-29, 8.598672e-29, 8.598662e-29, 8.598746e-29, 8.598778e-29, 
    8.598792e-29, 8.598804e-29, 8.598832e-29, 8.598813e-29, 8.59882e-29, 
    8.598802e-29, 8.59879e-29, 8.598796e-29, 8.598759e-29, 8.598773e-29, 
    8.598698e-29, 8.598731e-29, 8.598646e-29, 8.598667e-29, 8.598642e-29, 
    8.598654e-29, 8.598633e-29, 8.598652e-29, 8.598618e-29, 8.598611e-29, 
    8.598616e-29, 8.598597e-29, 8.598654e-29, 8.598631e-29, 8.598796e-29, 
    8.598795e-29, 8.59879e-29, 8.59881e-29, 8.598811e-29, 8.598829e-29, 
    8.598813e-29, 8.598807e-29, 8.598789e-29, 8.598779e-29, 8.598769e-29, 
    8.598748e-29, 8.598723e-29, 8.59869e-29, 8.598665e-29, 8.598649e-29, 
    8.598659e-29, 8.59865e-29, 8.59866e-29, 8.598665e-29, 8.598613e-29, 
    8.598642e-29, 8.5986e-29, 8.598602e-29, 8.598621e-29, 8.598601e-29, 
    8.598794e-29, 8.598799e-29, 8.598819e-29, 8.598804e-29, 8.598831e-29, 
    8.598816e-29, 8.598807e-29, 8.598773e-29, 8.598766e-29, 8.598758e-29, 
    8.598745e-29, 8.598727e-29, 8.598696e-29, 8.598669e-29, 8.598645e-29, 
    8.598646e-29, 8.598646e-29, 8.59864e-29, 8.598654e-29, 8.598638e-29, 
    8.598636e-29, 8.598642e-29, 8.598602e-29, 8.598613e-29, 8.598602e-29, 
    8.598609e-29, 8.598798e-29, 8.598788e-29, 8.598793e-29, 8.598784e-29, 
    8.598791e-29, 8.598761e-29, 8.598752e-29, 8.59871e-29, 8.598728e-29, 
    8.5987e-29, 8.598725e-29, 8.59872e-29, 8.598699e-29, 8.598723e-29, 
    8.598671e-29, 8.598707e-29, 8.59864e-29, 8.598676e-29, 8.598638e-29, 
    8.598645e-29, 8.598633e-29, 8.598623e-29, 8.59861e-29, 8.598586e-29, 
    8.598592e-29, 8.598572e-29, 8.598775e-29, 8.598763e-29, 8.598763e-29, 
    8.598751e-29, 8.598742e-29, 8.598721e-29, 8.598689e-29, 8.598701e-29, 
    8.598678e-29, 8.598674e-29, 8.598708e-29, 8.598687e-29, 8.598754e-29, 
    8.598743e-29, 8.59875e-29, 8.598773e-29, 8.598698e-29, 8.598737e-29, 
    8.598665e-29, 8.598686e-29, 8.598625e-29, 8.598655e-29, 8.598595e-29, 
    8.598569e-29, 8.598545e-29, 8.598516e-29, 8.598756e-29, 8.598764e-29, 
    8.598749e-29, 8.598729e-29, 8.59871e-29, 8.598685e-29, 8.598682e-29, 
    8.598678e-29, 8.598665e-29, 8.598655e-29, 8.598676e-29, 8.598652e-29, 
    8.598741e-29, 8.598695e-29, 8.598767e-29, 8.598745e-29, 8.59873e-29, 
    8.598737e-29, 8.598702e-29, 8.598694e-29, 8.598661e-29, 8.598678e-29, 
    8.598575e-29, 8.598621e-29, 8.598495e-29, 8.59853e-29, 8.598767e-29, 
    8.598756e-29, 8.598717e-29, 8.598736e-29, 8.598683e-29, 8.59867e-29, 
    8.59866e-29, 8.598646e-29, 8.598645e-29, 8.598637e-29, 8.59865e-29, 
    8.598637e-29, 8.598685e-29, 8.598663e-29, 8.598722e-29, 8.598707e-29, 
    8.598714e-29, 8.598721e-29, 8.598699e-29, 8.598676e-29, 8.598675e-29, 
    8.598668e-29, 8.598646e-29, 8.598683e-29, 8.59857e-29, 8.59864e-29, 
    8.598744e-29, 8.598722e-29, 8.598719e-29, 8.598728e-29, 8.598672e-29, 
    8.598692e-29, 8.598637e-29, 8.598652e-29, 8.598627e-29, 8.59864e-29, 
    8.598642e-29, 8.598657e-29, 8.598666e-29, 8.598691e-29, 8.598711e-29, 
    8.598727e-29, 8.598723e-29, 8.598705e-29, 8.598674e-29, 8.598645e-29, 
    8.598651e-29, 8.59863e-29, 8.598687e-29, 8.598663e-29, 8.598672e-29, 
    8.598648e-29, 8.598701e-29, 8.598655e-29, 8.598713e-29, 8.598708e-29, 
    8.598692e-29, 8.598661e-29, 8.598654e-29, 8.598647e-29, 8.598651e-29, 
    8.598674e-29, 8.598677e-29, 8.598693e-29, 8.598697e-29, 8.598709e-29, 
    8.598719e-29, 8.59871e-29, 8.5987e-29, 8.598674e-29, 8.598649e-29, 
    8.598623e-29, 8.598616e-29, 8.598586e-29, 8.598611e-29, 8.598569e-29, 
    8.598604e-29, 8.598544e-29, 8.598653e-29, 8.598606e-29, 8.598692e-29, 
    8.598683e-29, 8.598666e-29, 8.598627e-29, 8.598648e-29, 8.598624e-29, 
    8.598677e-29, 8.598705e-29, 8.598712e-29, 8.598725e-29, 8.598712e-29, 
    8.598713e-29, 8.5987e-29, 8.598704e-29, 8.598672e-29, 8.598689e-29, 
    8.598642e-29, 8.598624e-29, 8.598574e-29, 8.598544e-29, 8.598513e-29, 
    8.598499e-29, 8.598495e-29, 8.598493e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.135276e-08, 1.140281e-08, 1.139308e-08, 1.143345e-08, 1.141105e-08, 
    1.143749e-08, 1.136291e-08, 1.140479e-08, 1.137805e-08, 1.135727e-08, 
    1.151178e-08, 1.143525e-08, 1.15913e-08, 1.154248e-08, 1.166513e-08, 
    1.158371e-08, 1.168155e-08, 1.166278e-08, 1.171927e-08, 1.170308e-08, 
    1.177533e-08, 1.172674e-08, 1.181279e-08, 1.176373e-08, 1.17714e-08, 
    1.172513e-08, 1.145065e-08, 1.150225e-08, 1.144759e-08, 1.145495e-08, 
    1.145165e-08, 1.141152e-08, 1.139129e-08, 1.134894e-08, 1.135662e-08, 
    1.138773e-08, 1.145826e-08, 1.143432e-08, 1.149466e-08, 1.14933e-08, 
    1.156048e-08, 1.153019e-08, 1.164311e-08, 1.161101e-08, 1.170376e-08, 
    1.168043e-08, 1.170266e-08, 1.169592e-08, 1.170275e-08, 1.166854e-08, 
    1.16832e-08, 1.16531e-08, 1.153586e-08, 1.157031e-08, 1.146756e-08, 
    1.140577e-08, 1.136474e-08, 1.133563e-08, 1.133974e-08, 1.134759e-08, 
    1.138791e-08, 1.142583e-08, 1.145473e-08, 1.147406e-08, 1.14931e-08, 
    1.155075e-08, 1.158127e-08, 1.16496e-08, 1.163727e-08, 1.165815e-08, 
    1.167811e-08, 1.171162e-08, 1.170611e-08, 1.172087e-08, 1.165761e-08, 
    1.169965e-08, 1.163024e-08, 1.164923e-08, 1.149827e-08, 1.144078e-08, 
    1.141634e-08, 1.139495e-08, 1.134291e-08, 1.137885e-08, 1.136468e-08, 
    1.139838e-08, 1.14198e-08, 1.140921e-08, 1.147459e-08, 1.144917e-08, 
    1.158307e-08, 1.152539e-08, 1.167579e-08, 1.16398e-08, 1.168441e-08, 
    1.166165e-08, 1.170065e-08, 1.166555e-08, 1.172636e-08, 1.173961e-08, 
    1.173056e-08, 1.176532e-08, 1.16636e-08, 1.170266e-08, 1.140891e-08, 
    1.141064e-08, 1.141869e-08, 1.138331e-08, 1.138114e-08, 1.134872e-08, 
    1.137757e-08, 1.138986e-08, 1.142104e-08, 1.143949e-08, 1.145703e-08, 
    1.149558e-08, 1.153864e-08, 1.159886e-08, 1.164213e-08, 1.167113e-08, 
    1.165335e-08, 1.166905e-08, 1.16515e-08, 1.164327e-08, 1.173464e-08, 
    1.168334e-08, 1.176032e-08, 1.175606e-08, 1.172122e-08, 1.175654e-08, 
    1.141185e-08, 1.140191e-08, 1.13674e-08, 1.139441e-08, 1.134519e-08, 
    1.137274e-08, 1.138858e-08, 1.14497e-08, 1.146313e-08, 1.147558e-08, 
    1.150017e-08, 1.153174e-08, 1.158711e-08, 1.163529e-08, 1.167928e-08, 
    1.167605e-08, 1.167719e-08, 1.168701e-08, 1.166267e-08, 1.169101e-08, 
    1.169576e-08, 1.168333e-08, 1.175549e-08, 1.173487e-08, 1.175597e-08, 
    1.174255e-08, 1.140514e-08, 1.142187e-08, 1.141283e-08, 1.142983e-08, 
    1.141785e-08, 1.14711e-08, 1.148707e-08, 1.156177e-08, 1.153112e-08, 
    1.157991e-08, 1.153607e-08, 1.154384e-08, 1.15815e-08, 1.153844e-08, 
    1.163263e-08, 1.156877e-08, 1.168739e-08, 1.162362e-08, 1.169139e-08, 
    1.167909e-08, 1.169946e-08, 1.171771e-08, 1.174067e-08, 1.178303e-08, 
    1.177322e-08, 1.180865e-08, 1.144681e-08, 1.146851e-08, 1.14666e-08, 
    1.14893e-08, 1.15061e-08, 1.15425e-08, 1.160088e-08, 1.157893e-08, 
    1.161923e-08, 1.162732e-08, 1.156609e-08, 1.160369e-08, 1.148303e-08, 
    1.150252e-08, 1.149091e-08, 1.144852e-08, 1.158398e-08, 1.151446e-08, 
    1.164284e-08, 1.160518e-08, 1.171511e-08, 1.166044e-08, 1.176782e-08, 
    1.181373e-08, 1.185694e-08, 1.190743e-08, 1.148035e-08, 1.146561e-08, 
    1.1492e-08, 1.152853e-08, 1.156242e-08, 1.160748e-08, 1.161209e-08, 
    1.162053e-08, 1.164239e-08, 1.166078e-08, 1.16232e-08, 1.166539e-08, 
    1.150704e-08, 1.159002e-08, 1.146003e-08, 1.149917e-08, 1.152637e-08, 
    1.151444e-08, 1.157642e-08, 1.159103e-08, 1.165038e-08, 1.16197e-08, 
    1.180239e-08, 1.172156e-08, 1.194588e-08, 1.188319e-08, 1.146045e-08, 
    1.14803e-08, 1.154936e-08, 1.15165e-08, 1.161049e-08, 1.163362e-08, 
    1.165243e-08, 1.167647e-08, 1.167906e-08, 1.169331e-08, 1.166997e-08, 
    1.169239e-08, 1.160757e-08, 1.164547e-08, 1.154147e-08, 1.156678e-08, 
    1.155514e-08, 1.154237e-08, 1.158179e-08, 1.162379e-08, 1.162469e-08, 
    1.163815e-08, 1.16761e-08, 1.161087e-08, 1.181282e-08, 1.168809e-08, 
    1.150194e-08, 1.154016e-08, 1.154562e-08, 1.153081e-08, 1.16313e-08, 
    1.159489e-08, 1.169296e-08, 1.166646e-08, 1.170989e-08, 1.16883e-08, 
    1.168513e-08, 1.165741e-08, 1.164016e-08, 1.159656e-08, 1.156109e-08, 
    1.153296e-08, 1.15395e-08, 1.15704e-08, 1.162636e-08, 1.16793e-08, 
    1.16677e-08, 1.170659e-08, 1.160367e-08, 1.164682e-08, 1.163014e-08, 
    1.167363e-08, 1.157834e-08, 1.165948e-08, 1.15576e-08, 1.156654e-08, 
    1.159417e-08, 1.164975e-08, 1.166205e-08, 1.167518e-08, 1.166708e-08, 
    1.162778e-08, 1.162134e-08, 1.15935e-08, 1.158581e-08, 1.156459e-08, 
    1.154703e-08, 1.156307e-08, 1.157993e-08, 1.162779e-08, 1.167093e-08, 
    1.171797e-08, 1.172948e-08, 1.178443e-08, 1.17397e-08, 1.181352e-08, 
    1.175075e-08, 1.185941e-08, 1.166419e-08, 1.174891e-08, 1.159543e-08, 
    1.161196e-08, 1.164186e-08, 1.171046e-08, 1.167343e-08, 1.171674e-08, 
    1.162109e-08, 1.157146e-08, 1.155863e-08, 1.153467e-08, 1.155917e-08, 
    1.155718e-08, 1.158063e-08, 1.157309e-08, 1.162938e-08, 1.159915e-08, 
    1.168505e-08, 1.17164e-08, 1.180493e-08, 1.185921e-08, 1.191447e-08, 
    1.193887e-08, 1.194629e-08, 1.194939e-08 ;

 SOIL1N_TO_SOIL3N =
  1.347056e-10, 1.352997e-10, 1.351842e-10, 1.356634e-10, 1.353976e-10, 
    1.357113e-10, 1.348261e-10, 1.353233e-10, 1.350059e-10, 1.347591e-10, 
    1.365932e-10, 1.356847e-10, 1.375371e-10, 1.369577e-10, 1.384134e-10, 
    1.374469e-10, 1.386083e-10, 1.383856e-10, 1.390561e-10, 1.38864e-10, 
    1.397216e-10, 1.391448e-10, 1.401663e-10, 1.395839e-10, 1.39675e-10, 
    1.391258e-10, 1.358676e-10, 1.364801e-10, 1.358313e-10, 1.359186e-10, 
    1.358794e-10, 1.35403e-10, 1.35163e-10, 1.346603e-10, 1.347515e-10, 
    1.351208e-10, 1.359579e-10, 1.356738e-10, 1.3639e-10, 1.363738e-10, 
    1.371712e-10, 1.368117e-10, 1.381521e-10, 1.377711e-10, 1.38872e-10, 
    1.385951e-10, 1.38859e-10, 1.38779e-10, 1.388601e-10, 1.38454e-10, 
    1.38628e-10, 1.382707e-10, 1.36879e-10, 1.37288e-10, 1.360683e-10, 
    1.353349e-10, 1.348479e-10, 1.345023e-10, 1.345511e-10, 1.346443e-10, 
    1.351229e-10, 1.35573e-10, 1.35916e-10, 1.361454e-10, 1.363715e-10, 
    1.370557e-10, 1.37418e-10, 1.382291e-10, 1.380827e-10, 1.383307e-10, 
    1.385676e-10, 1.389654e-10, 1.388999e-10, 1.390751e-10, 1.383242e-10, 
    1.388232e-10, 1.379994e-10, 1.382247e-10, 1.364329e-10, 1.357504e-10, 
    1.354603e-10, 1.352064e-10, 1.345887e-10, 1.350153e-10, 1.348471e-10, 
    1.352472e-10, 1.355014e-10, 1.353757e-10, 1.361517e-10, 1.3585e-10, 
    1.374395e-10, 1.367548e-10, 1.3854e-10, 1.381128e-10, 1.386424e-10, 
    1.383721e-10, 1.388352e-10, 1.384184e-10, 1.391404e-10, 1.392975e-10, 
    1.391901e-10, 1.396028e-10, 1.383953e-10, 1.38859e-10, 1.353722e-10, 
    1.353927e-10, 1.354882e-10, 1.350682e-10, 1.350425e-10, 1.346577e-10, 
    1.350001e-10, 1.35146e-10, 1.355162e-10, 1.357351e-10, 1.359433e-10, 
    1.364009e-10, 1.369121e-10, 1.376269e-10, 1.381405e-10, 1.384847e-10, 
    1.382736e-10, 1.3846e-10, 1.382517e-10, 1.38154e-10, 1.392386e-10, 
    1.386296e-10, 1.395434e-10, 1.394929e-10, 1.390793e-10, 1.394986e-10, 
    1.354071e-10, 1.352891e-10, 1.348794e-10, 1.352e-10, 1.346158e-10, 
    1.349428e-10, 1.351308e-10, 1.358563e-10, 1.360157e-10, 1.361635e-10, 
    1.364554e-10, 1.368301e-10, 1.374873e-10, 1.380593e-10, 1.385814e-10, 
    1.385431e-10, 1.385566e-10, 1.386732e-10, 1.383843e-10, 1.387207e-10, 
    1.387771e-10, 1.386295e-10, 1.394861e-10, 1.392414e-10, 1.394918e-10, 
    1.393325e-10, 1.353274e-10, 1.35526e-10, 1.354187e-10, 1.356204e-10, 
    1.354783e-10, 1.361103e-10, 1.362998e-10, 1.371866e-10, 1.368227e-10, 
    1.374019e-10, 1.368815e-10, 1.369738e-10, 1.374208e-10, 1.369097e-10, 
    1.380277e-10, 1.372697e-10, 1.386778e-10, 1.379207e-10, 1.387252e-10, 
    1.385791e-10, 1.38821e-10, 1.390376e-10, 1.393102e-10, 1.39813e-10, 
    1.396966e-10, 1.401172e-10, 1.35822e-10, 1.360795e-10, 1.360569e-10, 
    1.363264e-10, 1.365257e-10, 1.369578e-10, 1.376508e-10, 1.373902e-10, 
    1.378687e-10, 1.379647e-10, 1.372378e-10, 1.376841e-10, 1.362519e-10, 
    1.364833e-10, 1.363455e-10, 1.358423e-10, 1.374502e-10, 1.36625e-10, 
    1.38149e-10, 1.377018e-10, 1.390067e-10, 1.383578e-10, 1.396325e-10, 
    1.401774e-10, 1.406904e-10, 1.412898e-10, 1.362201e-10, 1.360451e-10, 
    1.363585e-10, 1.36792e-10, 1.371943e-10, 1.377291e-10, 1.377839e-10, 
    1.378841e-10, 1.381436e-10, 1.383618e-10, 1.379157e-10, 1.384165e-10, 
    1.365369e-10, 1.375219e-10, 1.359789e-10, 1.364435e-10, 1.367664e-10, 
    1.366248e-10, 1.373604e-10, 1.375338e-10, 1.382384e-10, 1.378742e-10, 
    1.400429e-10, 1.390834e-10, 1.417463e-10, 1.41002e-10, 1.35984e-10, 
    1.362195e-10, 1.370393e-10, 1.366492e-10, 1.377648e-10, 1.380394e-10, 
    1.382627e-10, 1.385481e-10, 1.385789e-10, 1.38748e-10, 1.384709e-10, 
    1.38737e-10, 1.377303e-10, 1.381802e-10, 1.369456e-10, 1.372461e-10, 
    1.371079e-10, 1.369562e-10, 1.374242e-10, 1.379227e-10, 1.379334e-10, 
    1.380933e-10, 1.385437e-10, 1.377694e-10, 1.401667e-10, 1.38686e-10, 
    1.364764e-10, 1.3693e-10, 1.369949e-10, 1.368191e-10, 1.380119e-10, 
    1.375797e-10, 1.387439e-10, 1.384292e-10, 1.389448e-10, 1.386886e-10, 
    1.386509e-10, 1.383219e-10, 1.38117e-10, 1.375995e-10, 1.371785e-10, 
    1.368446e-10, 1.369223e-10, 1.37289e-10, 1.379532e-10, 1.385817e-10, 
    1.38444e-10, 1.389056e-10, 1.376839e-10, 1.381962e-10, 1.379982e-10, 
    1.385144e-10, 1.373833e-10, 1.383464e-10, 1.371371e-10, 1.372431e-10, 
    1.375711e-10, 1.382309e-10, 1.383769e-10, 1.385328e-10, 1.384366e-10, 
    1.379701e-10, 1.378937e-10, 1.375632e-10, 1.374719e-10, 1.372201e-10, 
    1.370116e-10, 1.37202e-10, 1.374021e-10, 1.379703e-10, 1.384824e-10, 
    1.390407e-10, 1.391774e-10, 1.398297e-10, 1.392986e-10, 1.401749e-10, 
    1.394298e-10, 1.407197e-10, 1.384023e-10, 1.39408e-10, 1.375861e-10, 
    1.377823e-10, 1.381373e-10, 1.389516e-10, 1.38512e-10, 1.390261e-10, 
    1.378907e-10, 1.373016e-10, 1.371493e-10, 1.368649e-10, 1.371557e-10, 
    1.371321e-10, 1.374104e-10, 1.37321e-10, 1.379892e-10, 1.376302e-10, 
    1.386499e-10, 1.390221e-10, 1.400731e-10, 1.407174e-10, 1.413734e-10, 
    1.416629e-10, 1.417511e-10, 1.417879e-10 ;

 SOIL1N_vr =
  2.497637, 2.49763, 2.497631, 2.497626, 2.497629, 2.497626, 2.497635, 
    2.49763, 2.497633, 2.497636, 2.497616, 2.497626, 2.497606, 2.497612, 
    2.497596, 2.497607, 2.497594, 2.497597, 2.497589, 2.497591, 2.497582, 
    2.497588, 2.497577, 2.497584, 2.497583, 2.497589, 2.497624, 2.497617, 
    2.497624, 2.497623, 2.497624, 2.497629, 2.497632, 2.497637, 2.497636, 
    2.497632, 2.497623, 2.497626, 2.497618, 2.497618, 2.49761, 2.497614, 
    2.497599, 2.497603, 2.497591, 2.497594, 2.497591, 2.497592, 2.497591, 
    2.497596, 2.497594, 2.497598, 2.497613, 2.497608, 2.497622, 2.49763, 
    2.497635, 2.497639, 2.497638, 2.497637, 2.497632, 2.497627, 2.497623, 
    2.497621, 2.497618, 2.497611, 2.497607, 2.497598, 2.4976, 2.497597, 
    2.497595, 2.49759, 2.497591, 2.497589, 2.497597, 2.497592, 2.497601, 
    2.497598, 2.497618, 2.497625, 2.497628, 2.497631, 2.497638, 2.497633, 
    2.497635, 2.497631, 2.497628, 2.497629, 2.497621, 2.497624, 2.497607, 
    2.497614, 2.497595, 2.4976, 2.497594, 2.497597, 2.497592, 2.497596, 
    2.497589, 2.497587, 2.497588, 2.497584, 2.497597, 2.497591, 2.497629, 
    2.497629, 2.497628, 2.497633, 2.497633, 2.497637, 2.497633, 2.497632, 
    2.497628, 2.497625, 2.497623, 2.497618, 2.497613, 2.497605, 2.497599, 
    2.497596, 2.497598, 2.497596, 2.497598, 2.497599, 2.497587, 2.497594, 
    2.497584, 2.497585, 2.497589, 2.497585, 2.497629, 2.49763, 2.497635, 
    2.497631, 2.497638, 2.497634, 2.497632, 2.497624, 2.497622, 2.497621, 
    2.497617, 2.497613, 2.497606, 2.4976, 2.497595, 2.497595, 2.497595, 
    2.497594, 2.497597, 2.497593, 2.497592, 2.497594, 2.497585, 2.497587, 
    2.497585, 2.497586, 2.49763, 2.497628, 2.497629, 2.497627, 2.497628, 
    2.497621, 2.497619, 2.49761, 2.497614, 2.497607, 2.497613, 2.497612, 
    2.497607, 2.497613, 2.497601, 2.497609, 2.497593, 2.497602, 2.497593, 
    2.497595, 2.497592, 2.49759, 2.497587, 2.497581, 2.497582, 2.497578, 
    2.497624, 2.497622, 2.497622, 2.497619, 2.497617, 2.497612, 2.497605, 
    2.497607, 2.497602, 2.497601, 2.497609, 2.497604, 2.49762, 2.497617, 
    2.497619, 2.497624, 2.497607, 2.497616, 2.497599, 2.497604, 2.49759, 
    2.497597, 2.497583, 2.497577, 2.497572, 2.497566, 2.49762, 2.497622, 
    2.497619, 2.497614, 2.49761, 2.497604, 2.497603, 2.497602, 2.497599, 
    2.497597, 2.497602, 2.497596, 2.497617, 2.497606, 2.497623, 2.497618, 
    2.497614, 2.497616, 2.497608, 2.497606, 2.497598, 2.497602, 2.497579, 
    2.497589, 2.497561, 2.497569, 2.497623, 2.49762, 2.497611, 2.497615, 
    2.497603, 2.4976, 2.497598, 2.497595, 2.497595, 2.497593, 2.497596, 
    2.497593, 2.497604, 2.497599, 2.497612, 2.497609, 2.497611, 2.497612, 
    2.497607, 2.497602, 2.497602, 2.4976, 2.497595, 2.497603, 2.497577, 
    2.497593, 2.497617, 2.497612, 2.497612, 2.497614, 2.497601, 2.497605, 
    2.497593, 2.497596, 2.497591, 2.497593, 2.497594, 2.497597, 2.4976, 
    2.497605, 2.49761, 2.497613, 2.497612, 2.497608, 2.497601, 2.497595, 
    2.497596, 2.497591, 2.497604, 2.497599, 2.497601, 2.497595, 2.497607, 
    2.497597, 2.49761, 2.497609, 2.497606, 2.497598, 2.497597, 2.497595, 
    2.497596, 2.497601, 2.497602, 2.497606, 2.497607, 2.497609, 2.497612, 
    2.497609, 2.497607, 2.497601, 2.497596, 2.49759, 2.497588, 2.497581, 
    2.497587, 2.497577, 2.497585, 2.497571, 2.497597, 2.497586, 2.497605, 
    2.497603, 2.497599, 2.497591, 2.497595, 2.49759, 2.497602, 2.497608, 
    2.49761, 2.497613, 2.49761, 2.49761, 2.497607, 2.497608, 2.497601, 
    2.497605, 2.497594, 2.49759, 2.497578, 2.497571, 2.497565, 2.497561, 
    2.497561, 2.49756,
  2.49791, 2.497902, 2.497903, 2.497897, 2.4979, 2.497896, 2.497908, 
    2.497901, 2.497906, 2.497909, 2.497885, 2.497897, 2.497872, 2.49788, 
    2.49786, 2.497873, 2.497858, 2.49786, 2.497851, 2.497854, 2.497843, 
    2.49785, 2.497837, 2.497844, 2.497843, 2.497851, 2.497894, 2.497886, 
    2.497895, 2.497893, 2.497894, 2.4979, 2.497904, 2.49791, 2.497909, 
    2.497904, 2.497893, 2.497897, 2.497887, 2.497887, 2.497877, 2.497881, 
    2.497864, 2.497869, 2.497854, 2.497858, 2.497854, 2.497855, 2.497854, 
    2.497859, 2.497857, 2.497862, 2.49788, 2.497875, 2.497891, 2.497901, 
    2.497908, 2.497912, 2.497912, 2.49791, 2.497904, 2.497898, 2.497894, 
    2.49789, 2.497887, 2.497878, 2.497873, 2.497863, 2.497864, 2.497861, 
    2.497858, 2.497853, 2.497854, 2.497851, 2.497861, 2.497854, 2.497866, 
    2.497863, 2.497887, 2.497896, 2.4979, 2.497903, 2.497911, 2.497905, 
    2.497908, 2.497902, 2.497899, 2.497901, 2.49789, 2.497894, 2.497873, 
    2.497882, 2.497858, 2.497864, 2.497857, 2.497861, 2.497854, 2.49786, 
    2.49785, 2.497848, 2.49785, 2.497844, 2.49786, 2.497854, 2.497901, 
    2.4979, 2.497899, 2.497905, 2.497905, 2.49791, 2.497906, 2.497904, 
    2.497899, 2.497896, 2.497893, 2.497887, 2.49788, 2.497871, 2.497864, 
    2.497859, 2.497862, 2.497859, 2.497862, 2.497864, 2.497849, 2.497857, 
    2.497845, 2.497846, 2.497851, 2.497846, 2.4979, 2.497902, 2.497907, 
    2.497903, 2.497911, 2.497906, 2.497904, 2.497894, 2.497892, 2.49789, 
    2.497886, 2.497881, 2.497872, 2.497865, 2.497858, 2.497858, 2.497858, 
    2.497857, 2.49786, 2.497856, 2.497855, 2.497857, 2.497846, 2.497849, 
    2.497846, 2.497848, 2.497901, 2.497899, 2.4979, 2.497897, 2.497899, 
    2.497891, 2.497888, 2.497876, 2.497881, 2.497874, 2.49788, 2.497879, 
    2.497873, 2.49788, 2.497865, 2.497875, 2.497857, 2.497867, 2.497856, 
    2.497858, 2.497855, 2.497852, 2.497848, 2.497841, 2.497843, 2.497837, 
    2.497895, 2.497891, 2.497892, 2.497888, 2.497885, 2.49788, 2.49787, 
    2.497874, 2.497867, 2.497866, 2.497876, 2.49787, 2.497889, 2.497886, 
    2.497888, 2.497895, 2.497873, 2.497884, 2.497864, 2.497869, 2.497852, 
    2.497861, 2.497844, 2.497837, 2.49783, 2.497822, 2.49789, 2.497892, 
    2.497888, 2.497882, 2.497876, 2.497869, 2.497869, 2.497867, 2.497864, 
    2.497861, 2.497867, 2.49786, 2.497885, 2.497872, 2.497893, 2.497886, 
    2.497882, 2.497884, 2.497874, 2.497872, 2.497862, 2.497867, 2.497838, 
    2.497851, 2.497816, 2.497826, 2.497893, 2.49789, 2.497878, 2.497884, 
    2.497869, 2.497865, 2.497862, 2.497858, 2.497858, 2.497856, 2.497859, 
    2.497856, 2.497869, 2.497863, 2.49788, 2.497876, 2.497878, 2.49788, 
    2.497873, 2.497867, 2.497866, 2.497864, 2.497858, 2.497869, 2.497837, 
    2.497856, 2.497886, 2.49788, 2.497879, 2.497881, 2.497865, 2.497871, 
    2.497856, 2.49786, 2.497853, 2.497856, 2.497857, 2.497861, 2.497864, 
    2.497871, 2.497877, 2.497881, 2.49788, 2.497875, 2.497866, 2.497858, 
    2.49786, 2.497854, 2.49787, 2.497863, 2.497866, 2.497859, 2.497874, 
    2.497861, 2.497877, 2.497876, 2.497871, 2.497863, 2.49786, 2.497859, 
    2.49786, 2.497866, 2.497867, 2.497871, 2.497873, 2.497876, 2.497879, 
    2.497876, 2.497874, 2.497866, 2.497859, 2.497852, 2.49785, 2.497841, 
    2.497848, 2.497837, 2.497847, 2.497829, 2.49786, 2.497847, 2.497871, 
    2.497869, 2.497864, 2.497853, 2.497859, 2.497852, 2.497867, 2.497875, 
    2.497877, 2.497881, 2.497877, 2.497877, 2.497874, 2.497875, 2.497866, 
    2.49787, 2.497857, 2.497852, 2.497838, 2.497829, 2.497821, 2.497817, 
    2.497816, 2.497815,
  2.498032, 2.498024, 2.498025, 2.498018, 2.498022, 2.498017, 2.49803, 
    2.498023, 2.498028, 2.498031, 2.498004, 2.498018, 2.497991, 2.497999, 
    2.497978, 2.497992, 2.497975, 2.497978, 2.497968, 2.497971, 2.497959, 
    2.497967, 2.497952, 2.497961, 2.497959, 2.497967, 2.498015, 2.498006, 
    2.498016, 2.498014, 2.498015, 2.498022, 2.498025, 2.498033, 2.498031, 
    2.498026, 2.498014, 2.498018, 2.498007, 2.498008, 2.497996, 2.498001, 
    2.497982, 2.497987, 2.497971, 2.497975, 2.497971, 2.497972, 2.497971, 
    2.497977, 2.497975, 2.49798, 2.498, 2.497994, 2.498012, 2.498023, 
    2.49803, 2.498035, 2.498034, 2.498033, 2.498026, 2.498019, 2.498014, 
    2.498011, 2.498008, 2.497998, 2.497992, 2.49798, 2.497983, 2.497979, 
    2.497976, 2.49797, 2.497971, 2.497968, 2.497979, 2.497972, 2.497984, 
    2.497981, 2.498007, 2.498017, 2.498021, 2.498025, 2.498034, 2.498028, 
    2.49803, 2.498024, 2.49802, 2.498022, 2.498011, 2.498015, 2.497992, 
    2.498002, 2.497976, 2.497982, 2.497974, 2.497978, 2.497972, 2.497978, 
    2.497967, 2.497965, 2.497966, 2.49796, 2.497978, 2.497971, 2.498022, 
    2.498022, 2.498021, 2.498027, 2.498027, 2.498033, 2.498028, 2.498026, 
    2.49802, 2.498017, 2.498014, 2.498007, 2.498, 2.497989, 2.497982, 
    2.497977, 2.49798, 2.497977, 2.49798, 2.497982, 2.497966, 2.497975, 
    2.497961, 2.497962, 2.497968, 2.497962, 2.498022, 2.498024, 2.498029, 
    2.498025, 2.498034, 2.498029, 2.498026, 2.498015, 2.498013, 2.498011, 
    2.498006, 2.498001, 2.497991, 2.497983, 2.497975, 2.497976, 2.497976, 
    2.497974, 2.497978, 2.497973, 2.497972, 2.497975, 2.497962, 2.497966, 
    2.497962, 2.497964, 2.498023, 2.49802, 2.498022, 2.498019, 2.498021, 
    2.498012, 2.498009, 2.497996, 2.498001, 2.497993, 2.498, 2.497999, 
    2.497992, 2.498, 2.497983, 2.497994, 2.497974, 2.497985, 2.497973, 
    2.497975, 2.497972, 2.497969, 2.497965, 2.497957, 2.497959, 2.497953, 
    2.498016, 2.498012, 2.498012, 2.498008, 2.498005, 2.497999, 2.497989, 
    2.497993, 2.497986, 2.497984, 2.497995, 2.497988, 2.498009, 2.498006, 
    2.498008, 2.498015, 2.497992, 2.498004, 2.497982, 2.497988, 2.497969, 
    2.497979, 2.49796, 2.497952, 2.497945, 2.497936, 2.49801, 2.498013, 
    2.498008, 2.498002, 2.497996, 2.497988, 2.497987, 2.497986, 2.497982, 
    2.497978, 2.497985, 2.497978, 2.498005, 2.497991, 2.498013, 2.498007, 
    2.498002, 2.498004, 2.497993, 2.497991, 2.49798, 2.497986, 2.497954, 
    2.497968, 2.497929, 2.49794, 2.498013, 2.49801, 2.497998, 2.498003, 
    2.497987, 2.497983, 2.49798, 2.497976, 2.497975, 2.497973, 2.497977, 
    2.497973, 2.497988, 2.497981, 2.497999, 2.497995, 2.497997, 2.497999, 
    2.497992, 2.497985, 2.497985, 2.497983, 2.497976, 2.497987, 2.497952, 
    2.497974, 2.498006, 2.497999, 2.497998, 2.498001, 2.497984, 2.49799, 
    2.497973, 2.497977, 2.49797, 2.497974, 2.497974, 2.497979, 2.497982, 
    2.49799, 2.497996, 2.498001, 2.498, 2.497994, 2.497984, 2.497975, 
    2.497977, 2.497971, 2.497988, 2.497981, 2.497984, 2.497976, 2.497993, 
    2.497979, 2.497996, 2.497995, 2.49799, 2.49798, 2.497978, 2.497976, 
    2.497977, 2.497984, 2.497985, 2.49799, 2.497992, 2.497995, 2.497998, 
    2.497995, 2.497993, 2.497984, 2.497977, 2.497969, 2.497967, 2.497957, 
    2.497965, 2.497952, 2.497963, 2.497944, 2.497978, 2.497963, 2.49799, 
    2.497987, 2.497982, 2.49797, 2.497976, 2.497969, 2.497985, 2.497994, 
    2.497996, 2.498, 2.497996, 2.497997, 2.497993, 2.497994, 2.497984, 
    2.497989, 2.497974, 2.497969, 2.497953, 2.497944, 2.497935, 2.49793, 
    2.497929, 2.497928,
  2.498126, 2.498117, 2.498119, 2.498111, 2.498116, 2.498111, 2.498124, 
    2.498116, 2.498121, 2.498125, 2.498098, 2.498111, 2.498083, 2.498092, 
    2.49807, 2.498085, 2.498067, 2.498071, 2.498061, 2.498064, 2.498051, 
    2.49806, 2.498044, 2.498053, 2.498051, 2.49806, 2.498108, 2.498099, 
    2.498109, 2.498108, 2.498108, 2.498115, 2.498119, 2.498127, 2.498125, 
    2.49812, 2.498107, 2.498111, 2.498101, 2.498101, 2.498089, 2.498094, 
    2.498074, 2.49808, 2.498064, 2.498068, 2.498064, 2.498065, 2.498064, 
    2.49807, 2.498067, 2.498072, 2.498093, 2.498087, 2.498106, 2.498116, 
    2.498124, 2.498129, 2.498128, 2.498127, 2.49812, 2.498113, 2.498108, 
    2.498104, 2.498101, 2.498091, 2.498085, 2.498073, 2.498075, 2.498072, 
    2.498068, 2.498062, 2.498063, 2.49806, 2.498072, 2.498064, 2.498076, 
    2.498073, 2.4981, 2.49811, 2.498115, 2.498118, 2.498128, 2.498121, 
    2.498124, 2.498118, 2.498114, 2.498116, 2.498104, 2.498109, 2.498085, 
    2.498095, 2.498069, 2.498075, 2.498067, 2.498071, 2.498064, 2.49807, 
    2.49806, 2.498057, 2.498059, 2.498053, 2.498071, 2.498064, 2.498116, 
    2.498116, 2.498114, 2.49812, 2.498121, 2.498127, 2.498122, 2.498119, 
    2.498114, 2.498111, 2.498107, 2.498101, 2.498093, 2.498082, 2.498075, 
    2.498069, 2.498072, 2.49807, 2.498073, 2.498074, 2.498058, 2.498067, 
    2.498054, 2.498054, 2.49806, 2.498054, 2.498115, 2.498117, 2.498123, 
    2.498118, 2.498127, 2.498122, 2.49812, 2.498109, 2.498106, 2.498104, 
    2.4981, 2.498094, 2.498084, 2.498076, 2.498068, 2.498068, 2.498068, 
    2.498066, 2.498071, 2.498066, 2.498065, 2.498067, 2.498054, 2.498058, 
    2.498054, 2.498057, 2.498116, 2.498114, 2.498115, 2.498112, 2.498114, 
    2.498105, 2.498102, 2.498089, 2.498094, 2.498085, 2.498093, 2.498092, 
    2.498085, 2.498093, 2.498076, 2.498087, 2.498066, 2.498078, 2.498066, 
    2.498068, 2.498064, 2.498061, 2.498057, 2.498049, 2.498051, 2.498045, 
    2.498109, 2.498105, 2.498106, 2.498101, 2.498099, 2.498092, 2.498082, 
    2.498086, 2.498079, 2.498077, 2.498088, 2.498081, 2.498103, 2.498099, 
    2.498101, 2.498109, 2.498085, 2.498097, 2.498074, 2.498081, 2.498061, 
    2.498071, 2.498052, 2.498044, 2.498036, 2.498027, 2.498103, 2.498106, 
    2.498101, 2.498095, 2.498089, 2.49808, 2.49808, 2.498078, 2.498074, 
    2.498071, 2.498078, 2.49807, 2.498098, 2.498084, 2.498107, 2.4981, 
    2.498095, 2.498097, 2.498086, 2.498084, 2.498073, 2.498078, 2.498046, 
    2.49806, 2.498021, 2.498032, 2.498107, 2.498103, 2.498091, 2.498097, 
    2.49808, 2.498076, 2.498073, 2.498068, 2.498068, 2.498065, 2.49807, 
    2.498065, 2.49808, 2.498074, 2.498092, 2.498088, 2.49809, 2.498092, 
    2.498085, 2.498078, 2.498078, 2.498075, 2.498068, 2.49808, 2.498044, 
    2.498066, 2.498099, 2.498093, 2.498091, 2.498094, 2.498076, 2.498083, 
    2.498065, 2.49807, 2.498062, 2.498066, 2.498067, 2.498072, 2.498075, 
    2.498083, 2.498089, 2.498094, 2.498093, 2.498087, 2.498077, 2.498068, 
    2.49807, 2.498063, 2.498081, 2.498074, 2.498077, 2.498069, 2.498086, 
    2.498071, 2.49809, 2.498088, 2.498083, 2.498073, 2.498071, 2.498069, 
    2.49807, 2.498077, 2.498078, 2.498083, 2.498085, 2.498088, 2.498091, 
    2.498088, 2.498085, 2.498077, 2.498069, 2.498061, 2.498059, 2.498049, 
    2.498057, 2.498044, 2.498055, 2.498036, 2.49807, 2.498055, 2.498083, 
    2.49808, 2.498075, 2.498062, 2.498069, 2.498061, 2.498078, 2.498087, 
    2.498089, 2.498094, 2.498089, 2.49809, 2.498085, 2.498087, 2.498077, 
    2.498082, 2.498067, 2.498061, 2.498045, 2.498036, 2.498026, 2.498022, 
    2.49802, 2.49802,
  2.498261, 2.498253, 2.498254, 2.498248, 2.498251, 2.498247, 2.498259, 
    2.498252, 2.498256, 2.49826, 2.498235, 2.498247, 2.498222, 2.49823, 
    2.49821, 2.498223, 2.498207, 2.49821, 2.498201, 2.498204, 2.498192, 
    2.4982, 2.498186, 2.498194, 2.498193, 2.4982, 2.498245, 2.498236, 
    2.498245, 2.498244, 2.498245, 2.498251, 2.498254, 2.498261, 2.49826, 
    2.498255, 2.498244, 2.498247, 2.498238, 2.498238, 2.498227, 2.498232, 
    2.498214, 2.498219, 2.498204, 2.498208, 2.498204, 2.498205, 2.498204, 
    2.498209, 2.498207, 2.498212, 2.498231, 2.498225, 2.498242, 2.498252, 
    2.498259, 2.498263, 2.498263, 2.498261, 2.498255, 2.498249, 2.498244, 
    2.498241, 2.498238, 2.498229, 2.498224, 2.498213, 2.498214, 2.498211, 
    2.498208, 2.498202, 2.498203, 2.498201, 2.498211, 2.498204, 2.498216, 
    2.498213, 2.498237, 2.498246, 2.49825, 2.498254, 2.498262, 2.498256, 
    2.498259, 2.498253, 2.49825, 2.498251, 2.498241, 2.498245, 2.498223, 
    2.498233, 2.498208, 2.498214, 2.498207, 2.49821, 2.498204, 2.49821, 
    2.4982, 2.498198, 2.498199, 2.498194, 2.49821, 2.498204, 2.498251, 
    2.498251, 2.49825, 2.498256, 2.498256, 2.498261, 2.498257, 2.498255, 
    2.49825, 2.498247, 2.498244, 2.498238, 2.49823, 2.498221, 2.498214, 
    2.498209, 2.498212, 2.498209, 2.498212, 2.498214, 2.498199, 2.498207, 
    2.498194, 2.498195, 2.498201, 2.498195, 2.498251, 2.498253, 2.498258, 
    2.498254, 2.498262, 2.498257, 2.498255, 2.498245, 2.498243, 2.498241, 
    2.498237, 2.498232, 2.498223, 2.498215, 2.498208, 2.498208, 2.498208, 
    2.498206, 2.49821, 2.498206, 2.498205, 2.498207, 2.498195, 2.498199, 
    2.498195, 2.498197, 2.498252, 2.49825, 2.498251, 2.498248, 2.49825, 
    2.498241, 2.498239, 2.498227, 2.498232, 2.498224, 2.498231, 2.49823, 
    2.498224, 2.49823, 2.498215, 2.498226, 2.498206, 2.498217, 2.498206, 
    2.498208, 2.498204, 2.498201, 2.498198, 2.498191, 2.498192, 2.498187, 
    2.498245, 2.498242, 2.498242, 2.498239, 2.498236, 2.49823, 2.49822, 
    2.498224, 2.498217, 2.498216, 2.498226, 2.49822, 2.49824, 2.498236, 
    2.498238, 2.498245, 2.498223, 2.498235, 2.498214, 2.49822, 2.498202, 
    2.498211, 2.498193, 2.498186, 2.498179, 2.498171, 2.49824, 2.498242, 
    2.498238, 2.498232, 2.498227, 2.498219, 2.498219, 2.498217, 2.498214, 
    2.498211, 2.498217, 2.49821, 2.498236, 2.498222, 2.498243, 2.498237, 
    2.498233, 2.498235, 2.498224, 2.498222, 2.498212, 2.498217, 2.498188, 
    2.498201, 2.498164, 2.498174, 2.498243, 2.49824, 2.498229, 2.498234, 
    2.498219, 2.498215, 2.498212, 2.498208, 2.498208, 2.498205, 2.498209, 
    2.498205, 2.498219, 2.498213, 2.49823, 2.498226, 2.498228, 2.49823, 
    2.498224, 2.498217, 2.498217, 2.498214, 2.498208, 2.498219, 2.498186, 
    2.498206, 2.498236, 2.49823, 2.498229, 2.498232, 2.498215, 2.498221, 
    2.498205, 2.49821, 2.498203, 2.498206, 2.498207, 2.498211, 2.498214, 
    2.498221, 2.498227, 2.498231, 2.49823, 2.498225, 2.498216, 2.498208, 
    2.498209, 2.498203, 2.49822, 2.498213, 2.498216, 2.498209, 2.498224, 
    2.498211, 2.498227, 2.498226, 2.498221, 2.498213, 2.49821, 2.498208, 
    2.49821, 2.498216, 2.498217, 2.498222, 2.498223, 2.498226, 2.498229, 
    2.498227, 2.498224, 2.498216, 2.498209, 2.498201, 2.498199, 2.498191, 
    2.498198, 2.498186, 2.498196, 2.498178, 2.49821, 2.498196, 2.498221, 
    2.498219, 2.498214, 2.498203, 2.498209, 2.498202, 2.498217, 2.498225, 
    2.498227, 2.498231, 2.498227, 2.498228, 2.498224, 2.498225, 2.498216, 
    2.498221, 2.498207, 2.498202, 2.498187, 2.498178, 2.498169, 2.498165, 
    2.498164, 2.498164,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  5.98301e-08, 6.00939e-08, 6.004262e-08, 6.02554e-08, 6.013737e-08, 
    6.02767e-08, 5.988359e-08, 6.010438e-08, 5.996343e-08, 5.985386e-08, 
    6.066833e-08, 6.02649e-08, 6.108748e-08, 6.083015e-08, 6.147663e-08, 
    6.104744e-08, 6.156317e-08, 6.146426e-08, 6.176201e-08, 6.167671e-08, 
    6.205753e-08, 6.180138e-08, 6.225498e-08, 6.199637e-08, 6.203682e-08, 
    6.179292e-08, 6.03461e-08, 6.06181e-08, 6.032997e-08, 6.036876e-08, 
    6.035136e-08, 6.01398e-08, 6.003319e-08, 5.980995e-08, 5.985048e-08, 
    6.001445e-08, 6.038621e-08, 6.026001e-08, 6.057807e-08, 6.057089e-08, 
    6.0925e-08, 6.076534e-08, 6.136055e-08, 6.119138e-08, 6.168027e-08, 
    6.155731e-08, 6.167449e-08, 6.163896e-08, 6.167495e-08, 6.149462e-08, 
    6.157188e-08, 6.141321e-08, 6.079524e-08, 6.097684e-08, 6.043521e-08, 
    6.010954e-08, 5.989327e-08, 5.97398e-08, 5.97615e-08, 5.980285e-08, 
    6.001541e-08, 6.021527e-08, 6.036758e-08, 6.046947e-08, 6.056986e-08, 
    6.087372e-08, 6.103458e-08, 6.139475e-08, 6.132976e-08, 6.143987e-08, 
    6.154508e-08, 6.17217e-08, 6.169263e-08, 6.177045e-08, 6.143697e-08, 
    6.16586e-08, 6.129274e-08, 6.13928e-08, 6.059711e-08, 6.029406e-08, 
    6.016522e-08, 6.005248e-08, 5.977817e-08, 5.99676e-08, 5.989293e-08, 
    6.007059e-08, 6.018348e-08, 6.012765e-08, 6.047225e-08, 6.033828e-08, 
    6.104411e-08, 6.074007e-08, 6.153281e-08, 6.13431e-08, 6.157828e-08, 
    6.145827e-08, 6.166389e-08, 6.147884e-08, 6.179941e-08, 6.186922e-08, 
    6.182151e-08, 6.200477e-08, 6.146858e-08, 6.167448e-08, 6.012608e-08, 
    6.013519e-08, 6.017761e-08, 5.999112e-08, 5.997972e-08, 5.980883e-08, 
    5.996089e-08, 6.002564e-08, 6.019003e-08, 6.028726e-08, 6.037969e-08, 
    6.058293e-08, 6.080991e-08, 6.112733e-08, 6.13554e-08, 6.150827e-08, 
    6.141454e-08, 6.14973e-08, 6.140478e-08, 6.136142e-08, 6.184305e-08, 
    6.15726e-08, 6.197841e-08, 6.195595e-08, 6.17723e-08, 6.195848e-08, 
    6.014158e-08, 6.008919e-08, 5.990725e-08, 6.004963e-08, 5.979022e-08, 
    5.993542e-08, 6.001891e-08, 6.034107e-08, 6.041186e-08, 6.04775e-08, 
    6.060714e-08, 6.077351e-08, 6.106537e-08, 6.131934e-08, 6.15512e-08, 
    6.153422e-08, 6.154019e-08, 6.159198e-08, 6.146369e-08, 6.161305e-08, 
    6.163811e-08, 6.157257e-08, 6.195295e-08, 6.184428e-08, 6.195548e-08, 
    6.188472e-08, 6.010622e-08, 6.019439e-08, 6.014675e-08, 6.023634e-08, 
    6.017321e-08, 6.045389e-08, 6.053804e-08, 6.093184e-08, 6.077023e-08, 
    6.102744e-08, 6.079636e-08, 6.08373e-08, 6.103582e-08, 6.080885e-08, 
    6.130533e-08, 6.096871e-08, 6.1594e-08, 6.125781e-08, 6.161507e-08, 
    6.15502e-08, 6.16576e-08, 6.175379e-08, 6.187481e-08, 6.209811e-08, 
    6.204641e-08, 6.223316e-08, 6.032585e-08, 6.044021e-08, 6.043015e-08, 
    6.054984e-08, 6.063836e-08, 6.083022e-08, 6.113797e-08, 6.102225e-08, 
    6.123471e-08, 6.127735e-08, 6.095458e-08, 6.115275e-08, 6.051675e-08, 
    6.061949e-08, 6.055833e-08, 6.033486e-08, 6.10489e-08, 6.068244e-08, 
    6.135917e-08, 6.116063e-08, 6.174007e-08, 6.145189e-08, 6.201794e-08, 
    6.225992e-08, 6.248771e-08, 6.275387e-08, 6.050263e-08, 6.042492e-08, 
    6.056407e-08, 6.075658e-08, 6.093524e-08, 6.117273e-08, 6.119704e-08, 
    6.124154e-08, 6.135679e-08, 6.14537e-08, 6.12556e-08, 6.1478e-08, 
    6.064331e-08, 6.108071e-08, 6.039554e-08, 6.060183e-08, 6.074524e-08, 
    6.068234e-08, 6.100902e-08, 6.108602e-08, 6.13989e-08, 6.123716e-08, 
    6.220019e-08, 6.17741e-08, 6.295657e-08, 6.262609e-08, 6.039777e-08, 
    6.050237e-08, 6.086641e-08, 6.06932e-08, 6.118859e-08, 6.131054e-08, 
    6.140968e-08, 6.15364e-08, 6.155009e-08, 6.162517e-08, 6.150213e-08, 
    6.162032e-08, 6.117324e-08, 6.137303e-08, 6.082481e-08, 6.095823e-08, 
    6.089685e-08, 6.082953e-08, 6.103733e-08, 6.125871e-08, 6.126346e-08, 
    6.133444e-08, 6.153446e-08, 6.11906e-08, 6.225516e-08, 6.159767e-08, 
    6.061643e-08, 6.08179e-08, 6.084669e-08, 6.076864e-08, 6.129832e-08, 
    6.110638e-08, 6.162335e-08, 6.148363e-08, 6.171256e-08, 6.15988e-08, 
    6.158206e-08, 6.143595e-08, 6.134499e-08, 6.111519e-08, 6.092822e-08, 
    6.077996e-08, 6.081444e-08, 6.097729e-08, 6.127226e-08, 6.155133e-08, 
    6.149019e-08, 6.169516e-08, 6.115268e-08, 6.138013e-08, 6.129222e-08, 
    6.152147e-08, 6.101917e-08, 6.144686e-08, 6.090985e-08, 6.095693e-08, 
    6.110258e-08, 6.139555e-08, 6.14604e-08, 6.15296e-08, 6.14869e-08, 
    6.127975e-08, 6.124581e-08, 6.109904e-08, 6.105851e-08, 6.094668e-08, 
    6.085409e-08, 6.093868e-08, 6.102752e-08, 6.127984e-08, 6.150723e-08, 
    6.175516e-08, 6.181584e-08, 6.210551e-08, 6.186968e-08, 6.225882e-08, 
    6.192796e-08, 6.250072e-08, 6.147167e-08, 6.191825e-08, 6.110921e-08, 
    6.119637e-08, 6.1354e-08, 6.171559e-08, 6.152039e-08, 6.174868e-08, 
    6.124449e-08, 6.09829e-08, 6.091524e-08, 6.078897e-08, 6.091813e-08, 
    6.090762e-08, 6.103121e-08, 6.09915e-08, 6.128822e-08, 6.112883e-08, 
    6.158164e-08, 6.174688e-08, 6.221359e-08, 6.249969e-08, 6.279098e-08, 
    6.291957e-08, 6.295871e-08, 6.297508e-08 ;

 SOIL1_HR_S3 =
  7.100462e-10, 7.131781e-10, 7.125693e-10, 7.150954e-10, 7.136942e-10, 
    7.153482e-10, 7.106812e-10, 7.133024e-10, 7.116291e-10, 7.103282e-10, 
    7.199978e-10, 7.152081e-10, 7.249742e-10, 7.219191e-10, 7.295943e-10, 
    7.244987e-10, 7.306219e-10, 7.294475e-10, 7.329826e-10, 7.319699e-10, 
    7.364914e-10, 7.334501e-10, 7.388357e-10, 7.357652e-10, 7.362455e-10, 
    7.333497e-10, 7.161721e-10, 7.194014e-10, 7.159808e-10, 7.164412e-10, 
    7.162346e-10, 7.13723e-10, 7.124573e-10, 7.098069e-10, 7.102881e-10, 
    7.122348e-10, 7.166483e-10, 7.151502e-10, 7.189263e-10, 7.18841e-10, 
    7.230451e-10, 7.211495e-10, 7.282162e-10, 7.262076e-10, 7.320121e-10, 
    7.305523e-10, 7.319435e-10, 7.315217e-10, 7.31949e-10, 7.29808e-10, 
    7.307253e-10, 7.288414e-10, 7.215045e-10, 7.236606e-10, 7.172301e-10, 
    7.133637e-10, 7.107961e-10, 7.089741e-10, 7.092317e-10, 7.097227e-10, 
    7.122462e-10, 7.14619e-10, 7.164273e-10, 7.176368e-10, 7.188287e-10, 
    7.224362e-10, 7.24346e-10, 7.286223e-10, 7.278507e-10, 7.29158e-10, 
    7.304071e-10, 7.325041e-10, 7.321589e-10, 7.330828e-10, 7.291236e-10, 
    7.317548e-10, 7.274111e-10, 7.285991e-10, 7.191522e-10, 7.155544e-10, 
    7.140247e-10, 7.126863e-10, 7.094297e-10, 7.116786e-10, 7.10792e-10, 
    7.129013e-10, 7.142416e-10, 7.135787e-10, 7.176699e-10, 7.160793e-10, 
    7.244592e-10, 7.208495e-10, 7.302614e-10, 7.28009e-10, 7.308013e-10, 
    7.293765e-10, 7.318177e-10, 7.296206e-10, 7.334268e-10, 7.342555e-10, 
    7.336892e-10, 7.358649e-10, 7.294988e-10, 7.319435e-10, 7.135601e-10, 
    7.136682e-10, 7.141719e-10, 7.119579e-10, 7.118224e-10, 7.097937e-10, 
    7.115989e-10, 7.123676e-10, 7.143193e-10, 7.154736e-10, 7.16571e-10, 
    7.189839e-10, 7.216787e-10, 7.254473e-10, 7.28155e-10, 7.299701e-10, 
    7.288572e-10, 7.298397e-10, 7.287413e-10, 7.282265e-10, 7.339449e-10, 
    7.307339e-10, 7.35552e-10, 7.352854e-10, 7.331048e-10, 7.353154e-10, 
    7.137441e-10, 7.131221e-10, 7.109621e-10, 7.126524e-10, 7.095728e-10, 
    7.112965e-10, 7.122877e-10, 7.161124e-10, 7.169529e-10, 7.177322e-10, 
    7.192713e-10, 7.212465e-10, 7.247117e-10, 7.277269e-10, 7.304797e-10, 
    7.302781e-10, 7.303491e-10, 7.30964e-10, 7.294407e-10, 7.312141e-10, 
    7.315116e-10, 7.307335e-10, 7.352496e-10, 7.339594e-10, 7.352797e-10, 
    7.344396e-10, 7.133243e-10, 7.143711e-10, 7.138054e-10, 7.148691e-10, 
    7.141197e-10, 7.174518e-10, 7.184509e-10, 7.231263e-10, 7.212076e-10, 
    7.242614e-10, 7.215178e-10, 7.220039e-10, 7.243608e-10, 7.216661e-10, 
    7.275606e-10, 7.23564e-10, 7.309879e-10, 7.269965e-10, 7.31238e-10, 
    7.304679e-10, 7.317431e-10, 7.328851e-10, 7.34322e-10, 7.369732e-10, 
    7.363593e-10, 7.385766e-10, 7.159317e-10, 7.172895e-10, 7.1717e-10, 
    7.18591e-10, 7.196419e-10, 7.219199e-10, 7.255736e-10, 7.241996e-10, 
    7.267221e-10, 7.272285e-10, 7.233963e-10, 7.257491e-10, 7.181982e-10, 
    7.19418e-10, 7.186918e-10, 7.160387e-10, 7.245161e-10, 7.201653e-10, 
    7.281998e-10, 7.258426e-10, 7.327223e-10, 7.293007e-10, 7.360214e-10, 
    7.388944e-10, 7.415989e-10, 7.447592e-10, 7.180306e-10, 7.17108e-10, 
    7.1876e-10, 7.210456e-10, 7.231666e-10, 7.259863e-10, 7.262749e-10, 
    7.268032e-10, 7.281716e-10, 7.293222e-10, 7.269701e-10, 7.296106e-10, 
    7.197007e-10, 7.248938e-10, 7.167591e-10, 7.192084e-10, 7.209109e-10, 
    7.201642e-10, 7.240427e-10, 7.249568e-10, 7.286716e-10, 7.267513e-10, 
    7.381852e-10, 7.331262e-10, 7.471659e-10, 7.43242e-10, 7.167856e-10, 
    7.180274e-10, 7.223495e-10, 7.20293e-10, 7.261747e-10, 7.276225e-10, 
    7.287995e-10, 7.303041e-10, 7.304666e-10, 7.31358e-10, 7.298972e-10, 
    7.313004e-10, 7.259924e-10, 7.283644e-10, 7.218556e-10, 7.234396e-10, 
    7.227109e-10, 7.219116e-10, 7.243787e-10, 7.270071e-10, 7.270634e-10, 
    7.279062e-10, 7.30281e-10, 7.261985e-10, 7.388379e-10, 7.310315e-10, 
    7.193816e-10, 7.217735e-10, 7.221153e-10, 7.211887e-10, 7.274773e-10, 
    7.251986e-10, 7.313363e-10, 7.296775e-10, 7.323955e-10, 7.310449e-10, 
    7.308462e-10, 7.291115e-10, 7.280315e-10, 7.253031e-10, 7.230833e-10, 
    7.213232e-10, 7.217324e-10, 7.236659e-10, 7.271679e-10, 7.304812e-10, 
    7.297554e-10, 7.32189e-10, 7.257482e-10, 7.284487e-10, 7.274049e-10, 
    7.301267e-10, 7.241631e-10, 7.292409e-10, 7.228652e-10, 7.234242e-10, 
    7.251534e-10, 7.286318e-10, 7.294017e-10, 7.302233e-10, 7.297163e-10, 
    7.272569e-10, 7.26854e-10, 7.251114e-10, 7.246302e-10, 7.233025e-10, 
    7.222032e-10, 7.232075e-10, 7.242623e-10, 7.27258e-10, 7.299577e-10, 
    7.329013e-10, 7.336218e-10, 7.37061e-10, 7.342611e-10, 7.388813e-10, 
    7.34953e-10, 7.417535e-10, 7.295355e-10, 7.348377e-10, 7.252322e-10, 
    7.262669e-10, 7.281385e-10, 7.324315e-10, 7.30114e-10, 7.328244e-10, 
    7.268382e-10, 7.237325e-10, 7.229292e-10, 7.214301e-10, 7.229635e-10, 
    7.228387e-10, 7.243061e-10, 7.238345e-10, 7.273575e-10, 7.254651e-10, 
    7.308411e-10, 7.32803e-10, 7.383442e-10, 7.417413e-10, 7.451998e-10, 
    7.467267e-10, 7.471914e-10, 7.473857e-10 ;

 SOIL2C =
  5.783957, 5.783963, 5.783962, 5.783967, 5.783964, 5.783967, 5.783958, 
    5.783963, 5.78396, 5.783957, 5.783976, 5.783967, 5.783985, 5.783979, 
    5.783994, 5.783985, 5.783996, 5.783994, 5.784001, 5.783999, 5.784008, 
    5.784002, 5.784012, 5.784006, 5.784007, 5.784001, 5.783968, 5.783975, 
    5.783968, 5.783969, 5.783968, 5.783964, 5.783961, 5.783956, 5.783957, 
    5.783961, 5.783969, 5.783967, 5.783974, 5.783974, 5.783982, 5.783978, 
    5.783992, 5.783988, 5.783999, 5.783996, 5.783999, 5.783998, 5.783999, 
    5.783995, 5.783997, 5.783993, 5.783979, 5.783983, 5.78397, 5.783963, 
    5.783958, 5.783955, 5.783955, 5.783956, 5.783961, 5.783966, 5.783969, 
    5.783971, 5.783974, 5.78398, 5.783984, 5.783992, 5.783991, 5.783993, 
    5.783996, 5.784, 5.783999, 5.784001, 5.783993, 5.783998, 5.78399, 
    5.783992, 5.783974, 5.783967, 5.783964, 5.783962, 5.783956, 5.78396, 
    5.783958, 5.783962, 5.783965, 5.783964, 5.783971, 5.783968, 5.783984, 
    5.783978, 5.783996, 5.783991, 5.783997, 5.783994, 5.783998, 5.783994, 
    5.784002, 5.784003, 5.784002, 5.784006, 5.783994, 5.783999, 5.783964, 
    5.783964, 5.783965, 5.78396, 5.78396, 5.783956, 5.78396, 5.783961, 
    5.783965, 5.783967, 5.783969, 5.783974, 5.783979, 5.783986, 5.783991, 
    5.783995, 5.783993, 5.783995, 5.783993, 5.783992, 5.784003, 5.783997, 
    5.784006, 5.784005, 5.784001, 5.784005, 5.783964, 5.783963, 5.783958, 
    5.783962, 5.783956, 5.783959, 5.783961, 5.783968, 5.78397, 5.783971, 
    5.783975, 5.783978, 5.783985, 5.783991, 5.783996, 5.783996, 5.783996, 
    5.783997, 5.783994, 5.783998, 5.783998, 5.783997, 5.784005, 5.784003, 
    5.784005, 5.784004, 5.783963, 5.783965, 5.783964, 5.783966, 5.783965, 
    5.783971, 5.783973, 5.783982, 5.783978, 5.783984, 5.783979, 5.78398, 
    5.783984, 5.783979, 5.78399, 5.783983, 5.783997, 5.783989, 5.783998, 
    5.783996, 5.783998, 5.784, 5.784003, 5.784009, 5.784007, 5.784011, 
    5.783968, 5.783971, 5.78397, 5.783973, 5.783975, 5.783979, 5.783987, 
    5.783984, 5.783989, 5.78399, 5.783982, 5.783987, 5.783972, 5.783975, 
    5.783973, 5.783968, 5.783985, 5.783976, 5.783991, 5.783987, 5.784, 
    5.783994, 5.784007, 5.784012, 5.784017, 5.784023, 5.783972, 5.78397, 
    5.783973, 5.783978, 5.783982, 5.783988, 5.783988, 5.783989, 5.783991, 
    5.783994, 5.783989, 5.783994, 5.783975, 5.783985, 5.783969, 5.783974, 
    5.783978, 5.783976, 5.783984, 5.783985, 5.783992, 5.783989, 5.784011, 
    5.784001, 5.784028, 5.78402, 5.78397, 5.783972, 5.78398, 5.783977, 
    5.783988, 5.78399, 5.783993, 5.783996, 5.783996, 5.783998, 5.783995, 
    5.783998, 5.783988, 5.783992, 5.783979, 5.783982, 5.783981, 5.783979, 
    5.783984, 5.783989, 5.783989, 5.783991, 5.783996, 5.783988, 5.784012, 
    5.783997, 5.783975, 5.783979, 5.78398, 5.783978, 5.78399, 5.783986, 
    5.783998, 5.783994, 5.783999, 5.783997, 5.783997, 5.783993, 5.783991, 
    5.783986, 5.783982, 5.783978, 5.783979, 5.783983, 5.783989, 5.783996, 
    5.783995, 5.783999, 5.783987, 5.783992, 5.78399, 5.783995, 5.783984, 
    5.783994, 5.783981, 5.783982, 5.783986, 5.783992, 5.783994, 5.783996, 
    5.783995, 5.78399, 5.783989, 5.783986, 5.783985, 5.783982, 5.78398, 
    5.783982, 5.783984, 5.78399, 5.783995, 5.784, 5.784002, 5.784009, 
    5.784003, 5.784012, 5.784005, 5.784018, 5.783994, 5.784004, 5.783986, 
    5.783988, 5.783991, 5.784, 5.783995, 5.784, 5.783989, 5.783983, 5.783981, 
    5.783978, 5.783981, 5.783981, 5.783984, 5.783983, 5.78399, 5.783986, 
    5.783997, 5.784, 5.784011, 5.784018, 5.784024, 5.784027, 5.784028, 
    5.784029 ;

 SOIL2C_TO_SOIL1C =
  1.058451e-09, 1.063122e-09, 1.062214e-09, 1.065981e-09, 1.063891e-09, 
    1.066358e-09, 1.059398e-09, 1.063307e-09, 1.060812e-09, 1.058872e-09, 
    1.073291e-09, 1.066149e-09, 1.080712e-09, 1.076156e-09, 1.087601e-09, 
    1.080003e-09, 1.089134e-09, 1.087383e-09, 1.092654e-09, 1.091144e-09, 
    1.097886e-09, 1.093351e-09, 1.101382e-09, 1.096803e-09, 1.097519e-09, 
    1.093201e-09, 1.067586e-09, 1.072402e-09, 1.067301e-09, 1.067988e-09, 
    1.06768e-09, 1.063934e-09, 1.062047e-09, 1.058095e-09, 1.058812e-09, 
    1.061715e-09, 1.068297e-09, 1.066062e-09, 1.071693e-09, 1.071566e-09, 
    1.077835e-09, 1.075009e-09, 1.085546e-09, 1.082551e-09, 1.091207e-09, 
    1.08903e-09, 1.091104e-09, 1.090475e-09, 1.091113e-09, 1.08792e-09, 
    1.089288e-09, 1.086479e-09, 1.075538e-09, 1.078753e-09, 1.069164e-09, 
    1.063398e-09, 1.05957e-09, 1.056853e-09, 1.057237e-09, 1.057969e-09, 
    1.061732e-09, 1.06527e-09, 1.067967e-09, 1.069771e-09, 1.071548e-09, 
    1.076927e-09, 1.079775e-09, 1.086152e-09, 1.085001e-09, 1.086951e-09, 
    1.088813e-09, 1.09194e-09, 1.091426e-09, 1.092803e-09, 1.086899e-09, 
    1.090823e-09, 1.084346e-09, 1.086117e-09, 1.07203e-09, 1.066665e-09, 
    1.064384e-09, 1.062388e-09, 1.057532e-09, 1.060886e-09, 1.059564e-09, 
    1.062709e-09, 1.064708e-09, 1.063719e-09, 1.06982e-09, 1.067448e-09, 
    1.079944e-09, 1.074561e-09, 1.088596e-09, 1.085238e-09, 1.089401e-09, 
    1.087277e-09, 1.090917e-09, 1.087641e-09, 1.093316e-09, 1.094552e-09, 
    1.093707e-09, 1.096952e-09, 1.087459e-09, 1.091104e-09, 1.063691e-09, 
    1.063853e-09, 1.064604e-09, 1.061302e-09, 1.0611e-09, 1.058075e-09, 
    1.060767e-09, 1.061913e-09, 1.064823e-09, 1.066545e-09, 1.068181e-09, 
    1.071779e-09, 1.075798e-09, 1.081418e-09, 1.085455e-09, 1.088162e-09, 
    1.086502e-09, 1.087967e-09, 1.086329e-09, 1.085562e-09, 1.094089e-09, 
    1.089301e-09, 1.096485e-09, 1.096088e-09, 1.092836e-09, 1.096132e-09, 
    1.063966e-09, 1.063038e-09, 1.059817e-09, 1.062338e-09, 1.057745e-09, 
    1.060316e-09, 1.061794e-09, 1.067497e-09, 1.068751e-09, 1.069913e-09, 
    1.072208e-09, 1.075153e-09, 1.080321e-09, 1.084817e-09, 1.088922e-09, 
    1.088621e-09, 1.088727e-09, 1.089644e-09, 1.087372e-09, 1.090017e-09, 
    1.09046e-09, 1.0893e-09, 1.096034e-09, 1.09411e-09, 1.096079e-09, 
    1.094827e-09, 1.06334e-09, 1.064901e-09, 1.064057e-09, 1.065643e-09, 
    1.064526e-09, 1.069495e-09, 1.070985e-09, 1.077957e-09, 1.075095e-09, 
    1.079649e-09, 1.075558e-09, 1.076283e-09, 1.079797e-09, 1.075779e-09, 
    1.084569e-09, 1.078609e-09, 1.089679e-09, 1.083728e-09, 1.090052e-09, 
    1.088904e-09, 1.090806e-09, 1.092509e-09, 1.094651e-09, 1.098604e-09, 
    1.097689e-09, 1.100995e-09, 1.067228e-09, 1.069253e-09, 1.069074e-09, 
    1.071193e-09, 1.072761e-09, 1.076157e-09, 1.081606e-09, 1.079557e-09, 
    1.083319e-09, 1.084074e-09, 1.078359e-09, 1.081867e-09, 1.070608e-09, 
    1.072427e-09, 1.071344e-09, 1.067388e-09, 1.080029e-09, 1.073541e-09, 
    1.085522e-09, 1.082007e-09, 1.092266e-09, 1.087164e-09, 1.097185e-09, 
    1.101469e-09, 1.105502e-09, 1.110214e-09, 1.070358e-09, 1.068982e-09, 
    1.071445e-09, 1.074854e-09, 1.078017e-09, 1.082221e-09, 1.082652e-09, 
    1.083439e-09, 1.08548e-09, 1.087196e-09, 1.083688e-09, 1.087626e-09, 
    1.072848e-09, 1.080592e-09, 1.068462e-09, 1.072114e-09, 1.074653e-09, 
    1.073539e-09, 1.079323e-09, 1.080686e-09, 1.086225e-09, 1.083362e-09, 
    1.100412e-09, 1.092868e-09, 1.113803e-09, 1.107952e-09, 1.068501e-09, 
    1.070353e-09, 1.076798e-09, 1.073732e-09, 1.082502e-09, 1.084661e-09, 
    1.086416e-09, 1.08866e-09, 1.088902e-09, 1.090231e-09, 1.088053e-09, 
    1.090145e-09, 1.08223e-09, 1.085767e-09, 1.076062e-09, 1.078424e-09, 
    1.077337e-09, 1.076145e-09, 1.079824e-09, 1.083743e-09, 1.083827e-09, 
    1.085084e-09, 1.088625e-09, 1.082538e-09, 1.101385e-09, 1.089745e-09, 
    1.072372e-09, 1.075939e-09, 1.076449e-09, 1.075067e-09, 1.084445e-09, 
    1.081047e-09, 1.090199e-09, 1.087725e-09, 1.091778e-09, 1.089764e-09, 
    1.089468e-09, 1.086881e-09, 1.085271e-09, 1.081202e-09, 1.077892e-09, 
    1.075268e-09, 1.075878e-09, 1.078761e-09, 1.083983e-09, 1.088924e-09, 
    1.087842e-09, 1.09147e-09, 1.081866e-09, 1.085893e-09, 1.084337e-09, 
    1.088395e-09, 1.079503e-09, 1.087075e-09, 1.077567e-09, 1.078401e-09, 
    1.080979e-09, 1.086166e-09, 1.087314e-09, 1.088539e-09, 1.087783e-09, 
    1.084116e-09, 1.083515e-09, 1.080917e-09, 1.080199e-09, 1.078219e-09, 
    1.07658e-09, 1.078078e-09, 1.07965e-09, 1.084118e-09, 1.088143e-09, 
    1.092533e-09, 1.093607e-09, 1.098735e-09, 1.09456e-09, 1.10145e-09, 
    1.095592e-09, 1.105732e-09, 1.087514e-09, 1.09542e-09, 1.081097e-09, 
    1.08264e-09, 1.085431e-09, 1.091832e-09, 1.088376e-09, 1.092418e-09, 
    1.083492e-09, 1.07886e-09, 1.077663e-09, 1.075427e-09, 1.077714e-09, 
    1.077528e-09, 1.079716e-09, 1.079013e-09, 1.084266e-09, 1.081444e-09, 
    1.089461e-09, 1.092386e-09, 1.100649e-09, 1.105714e-09, 1.110871e-09, 
    1.113148e-09, 1.113841e-09, 1.114131e-09 ;

 SOIL2C_TO_SOIL3C =
  7.560366e-11, 7.593726e-11, 7.587241e-11, 7.614148e-11, 7.599223e-11, 
    7.616841e-11, 7.56713e-11, 7.59505e-11, 7.577227e-11, 7.563371e-11, 
    7.666366e-11, 7.615349e-11, 7.719372e-11, 7.68683e-11, 7.768582e-11, 
    7.714307e-11, 7.779526e-11, 7.767018e-11, 7.804671e-11, 7.793884e-11, 
    7.842043e-11, 7.809649e-11, 7.867012e-11, 7.834308e-11, 7.839423e-11, 
    7.808581e-11, 7.625617e-11, 7.660014e-11, 7.623579e-11, 7.628484e-11, 
    7.626283e-11, 7.599531e-11, 7.586048e-11, 7.557818e-11, 7.562943e-11, 
    7.583678e-11, 7.630689e-11, 7.614732e-11, 7.654953e-11, 7.654045e-11, 
    7.698824e-11, 7.678633e-11, 7.753903e-11, 7.73251e-11, 7.794334e-11, 
    7.778785e-11, 7.793603e-11, 7.78911e-11, 7.793662e-11, 7.770858e-11, 
    7.780628e-11, 7.760563e-11, 7.682414e-11, 7.70538e-11, 7.636886e-11, 
    7.595703e-11, 7.568354e-11, 7.548947e-11, 7.551691e-11, 7.55692e-11, 
    7.5838e-11, 7.609074e-11, 7.628335e-11, 7.641218e-11, 7.653914e-11, 
    7.692338e-11, 7.712681e-11, 7.758228e-11, 7.75001e-11, 7.763934e-11, 
    7.777239e-11, 7.799574e-11, 7.795898e-11, 7.805738e-11, 7.763568e-11, 
    7.791594e-11, 7.745328e-11, 7.757982e-11, 7.657359e-11, 7.619037e-11, 
    7.602744e-11, 7.588487e-11, 7.5538e-11, 7.577754e-11, 7.568311e-11, 
    7.590778e-11, 7.605053e-11, 7.597994e-11, 7.641571e-11, 7.624629e-11, 
    7.713886e-11, 7.675439e-11, 7.775686e-11, 7.751697e-11, 7.781437e-11, 
    7.766261e-11, 7.792263e-11, 7.768862e-11, 7.809401e-11, 7.818228e-11, 
    7.812196e-11, 7.83537e-11, 7.767564e-11, 7.793603e-11, 7.597795e-11, 
    7.598946e-11, 7.604312e-11, 7.580728e-11, 7.579287e-11, 7.557677e-11, 
    7.576905e-11, 7.585094e-11, 7.605882e-11, 7.618177e-11, 7.629866e-11, 
    7.655566e-11, 7.68427e-11, 7.724411e-11, 7.753252e-11, 7.772585e-11, 
    7.76073e-11, 7.771196e-11, 7.759497e-11, 7.754013e-11, 7.81492e-11, 
    7.780719e-11, 7.832037e-11, 7.829198e-11, 7.805972e-11, 7.829518e-11, 
    7.599756e-11, 7.593129e-11, 7.570122e-11, 7.588127e-11, 7.555324e-11, 
    7.573685e-11, 7.584242e-11, 7.624981e-11, 7.633934e-11, 7.642234e-11, 
    7.658628e-11, 7.679667e-11, 7.716576e-11, 7.748692e-11, 7.778013e-11, 
    7.775864e-11, 7.776621e-11, 7.78317e-11, 7.766946e-11, 7.785834e-11, 
    7.789003e-11, 7.780716e-11, 7.828817e-11, 7.815074e-11, 7.829137e-11, 
    7.82019e-11, 7.595283e-11, 7.606433e-11, 7.600408e-11, 7.611738e-11, 
    7.603756e-11, 7.639248e-11, 7.64989e-11, 7.699689e-11, 7.679252e-11, 
    7.711779e-11, 7.682557e-11, 7.687734e-11, 7.712838e-11, 7.684137e-11, 
    7.74692e-11, 7.704352e-11, 7.783425e-11, 7.740911e-11, 7.786089e-11, 
    7.777886e-11, 7.791468e-11, 7.803632e-11, 7.818936e-11, 7.847174e-11, 
    7.840636e-11, 7.864253e-11, 7.623056e-11, 7.637518e-11, 7.636246e-11, 
    7.651382e-11, 7.662575e-11, 7.686839e-11, 7.725756e-11, 7.711122e-11, 
    7.737989e-11, 7.743383e-11, 7.702565e-11, 7.727625e-11, 7.647198e-11, 
    7.660191e-11, 7.652456e-11, 7.624196e-11, 7.714492e-11, 7.66815e-11, 
    7.753728e-11, 7.728621e-11, 7.801897e-11, 7.765454e-11, 7.837036e-11, 
    7.867636e-11, 7.896443e-11, 7.930102e-11, 7.645412e-11, 7.635585e-11, 
    7.653182e-11, 7.677527e-11, 7.700118e-11, 7.730153e-11, 7.733226e-11, 
    7.738853e-11, 7.753428e-11, 7.765683e-11, 7.740631e-11, 7.768755e-11, 
    7.663202e-11, 7.718515e-11, 7.631869e-11, 7.657958e-11, 7.676092e-11, 
    7.668138e-11, 7.70945e-11, 7.719186e-11, 7.758753e-11, 7.7383e-11, 
    7.860083e-11, 7.8062e-11, 7.955735e-11, 7.913942e-11, 7.632152e-11, 
    7.645379e-11, 7.691416e-11, 7.669511e-11, 7.732158e-11, 7.747579e-11, 
    7.760116e-11, 7.776142e-11, 7.777872e-11, 7.787367e-11, 7.771808e-11, 
    7.786753e-11, 7.730216e-11, 7.755481e-11, 7.686154e-11, 7.703026e-11, 
    7.695265e-11, 7.686751e-11, 7.713029e-11, 7.741024e-11, 7.741625e-11, 
    7.750602e-11, 7.775895e-11, 7.732412e-11, 7.867034e-11, 7.78389e-11, 
    7.659803e-11, 7.68528e-11, 7.688921e-11, 7.679051e-11, 7.746033e-11, 
    7.721762e-11, 7.787136e-11, 7.769468e-11, 7.798417e-11, 7.784032e-11, 
    7.781915e-11, 7.763439e-11, 7.751936e-11, 7.722874e-11, 7.699231e-11, 
    7.680483e-11, 7.684842e-11, 7.705436e-11, 7.742738e-11, 7.778028e-11, 
    7.770298e-11, 7.796218e-11, 7.727616e-11, 7.75638e-11, 7.745262e-11, 
    7.774253e-11, 7.710733e-11, 7.764818e-11, 7.696908e-11, 7.702862e-11, 
    7.721281e-11, 7.75833e-11, 7.76653e-11, 7.775282e-11, 7.769881e-11, 
    7.743685e-11, 7.739394e-11, 7.720833e-11, 7.715708e-11, 7.701566e-11, 
    7.689857e-11, 7.700555e-11, 7.711789e-11, 7.743697e-11, 7.772452e-11, 
    7.803805e-11, 7.811479e-11, 7.848109e-11, 7.818288e-11, 7.867498e-11, 
    7.825657e-11, 7.898089e-11, 7.767955e-11, 7.824429e-11, 7.722119e-11, 
    7.733141e-11, 7.753075e-11, 7.7988e-11, 7.774117e-11, 7.802985e-11, 
    7.739226e-11, 7.706146e-11, 7.69759e-11, 7.681623e-11, 7.697955e-11, 
    7.696627e-11, 7.712255e-11, 7.707233e-11, 7.744756e-11, 7.7246e-11, 
    7.781861e-11, 7.802758e-11, 7.861777e-11, 7.897959e-11, 7.934794e-11, 
    7.951056e-11, 7.956006e-11, 7.958075e-11 ;

 SOIL2C_vr =
  20.00591, 20.00593, 20.00593, 20.00594, 20.00593, 20.00594, 20.00592, 
    20.00593, 20.00592, 20.00591, 20.00596, 20.00594, 20.00599, 20.00597, 
    20.00601, 20.00599, 20.00602, 20.00601, 20.00603, 20.00603, 20.00605, 
    20.00603, 20.00606, 20.00604, 20.00605, 20.00603, 20.00594, 20.00596, 
    20.00594, 20.00595, 20.00595, 20.00593, 20.00592, 20.00591, 20.00591, 
    20.00592, 20.00595, 20.00594, 20.00596, 20.00596, 20.00598, 20.00597, 
    20.00601, 20.00599, 20.00603, 20.00602, 20.00603, 20.00602, 20.00603, 
    20.00601, 20.00602, 20.00601, 20.00597, 20.00598, 20.00595, 20.00593, 
    20.00592, 20.00591, 20.00591, 20.00591, 20.00592, 20.00594, 20.00595, 
    20.00595, 20.00596, 20.00598, 20.00599, 20.00601, 20.006, 20.00601, 
    20.00602, 20.00603, 20.00603, 20.00603, 20.00601, 20.00602, 20.006, 
    20.00601, 20.00596, 20.00594, 20.00593, 20.00593, 20.00591, 20.00592, 
    20.00592, 20.00593, 20.00593, 20.00593, 20.00595, 20.00594, 20.00599, 
    20.00597, 20.00602, 20.006, 20.00602, 20.00601, 20.00602, 20.00601, 
    20.00603, 20.00604, 20.00603, 20.00604, 20.00601, 20.00603, 20.00593, 
    20.00593, 20.00593, 20.00592, 20.00592, 20.00591, 20.00592, 20.00592, 
    20.00593, 20.00594, 20.00595, 20.00596, 20.00597, 20.00599, 20.00601, 
    20.00601, 20.00601, 20.00601, 20.00601, 20.00601, 20.00603, 20.00602, 
    20.00604, 20.00604, 20.00603, 20.00604, 20.00593, 20.00593, 20.00592, 
    20.00593, 20.00591, 20.00592, 20.00592, 20.00594, 20.00595, 20.00595, 
    20.00596, 20.00597, 20.00599, 20.006, 20.00602, 20.00602, 20.00602, 
    20.00602, 20.00601, 20.00602, 20.00602, 20.00602, 20.00604, 20.00603, 
    20.00604, 20.00604, 20.00593, 20.00593, 20.00593, 20.00594, 20.00593, 
    20.00595, 20.00595, 20.00598, 20.00597, 20.00599, 20.00597, 20.00597, 
    20.00599, 20.00597, 20.006, 20.00598, 20.00602, 20.006, 20.00602, 
    20.00602, 20.00602, 20.00603, 20.00604, 20.00605, 20.00605, 20.00606, 
    20.00594, 20.00595, 20.00595, 20.00596, 20.00596, 20.00597, 20.00599, 
    20.00599, 20.006, 20.006, 20.00598, 20.00599, 20.00595, 20.00596, 
    20.00596, 20.00594, 20.00599, 20.00596, 20.00601, 20.00599, 20.00603, 
    20.00601, 20.00605, 20.00606, 20.00607, 20.00609, 20.00595, 20.00595, 
    20.00596, 20.00597, 20.00598, 20.00599, 20.006, 20.006, 20.00601, 
    20.00601, 20.006, 20.00601, 20.00596, 20.00599, 20.00595, 20.00596, 
    20.00597, 20.00596, 20.00599, 20.00599, 20.00601, 20.006, 20.00606, 
    20.00603, 20.0061, 20.00608, 20.00595, 20.00595, 20.00598, 20.00596, 
    20.00599, 20.006, 20.00601, 20.00602, 20.00602, 20.00602, 20.00601, 
    20.00602, 20.00599, 20.00601, 20.00597, 20.00598, 20.00598, 20.00597, 
    20.00599, 20.006, 20.006, 20.006, 20.00602, 20.00599, 20.00606, 20.00602, 
    20.00596, 20.00597, 20.00597, 20.00597, 20.006, 20.00599, 20.00602, 
    20.00601, 20.00603, 20.00602, 20.00602, 20.00601, 20.006, 20.00599, 
    20.00598, 20.00597, 20.00597, 20.00598, 20.006, 20.00602, 20.00601, 
    20.00603, 20.00599, 20.00601, 20.006, 20.00602, 20.00599, 20.00601, 
    20.00598, 20.00598, 20.00599, 20.00601, 20.00601, 20.00602, 20.00601, 
    20.006, 20.006, 20.00599, 20.00599, 20.00598, 20.00598, 20.00598, 
    20.00599, 20.006, 20.00601, 20.00603, 20.00603, 20.00605, 20.00604, 
    20.00606, 20.00604, 20.00607, 20.00601, 20.00604, 20.00599, 20.006, 
    20.00601, 20.00603, 20.00602, 20.00603, 20.006, 20.00598, 20.00598, 
    20.00597, 20.00598, 20.00598, 20.00599, 20.00598, 20.006, 20.00599, 
    20.00602, 20.00603, 20.00606, 20.00607, 20.00609, 20.0061, 20.0061, 
    20.0061,
  20.00534, 20.00536, 20.00536, 20.00538, 20.00537, 20.00538, 20.00535, 
    20.00537, 20.00535, 20.00535, 20.00541, 20.00538, 20.00544, 20.00542, 
    20.00547, 20.00544, 20.00548, 20.00547, 20.00549, 20.00549, 20.00552, 
    20.0055, 20.00553, 20.00551, 20.00551, 20.0055, 20.00538, 20.0054, 
    20.00538, 20.00538, 20.00538, 20.00537, 20.00536, 20.00534, 20.00534, 
    20.00536, 20.00539, 20.00538, 20.0054, 20.0054, 20.00543, 20.00541, 
    20.00546, 20.00545, 20.00549, 20.00548, 20.00549, 20.00548, 20.00549, 
    20.00547, 20.00548, 20.00547, 20.00542, 20.00543, 20.00539, 20.00537, 
    20.00535, 20.00534, 20.00534, 20.00534, 20.00536, 20.00537, 20.00538, 
    20.00539, 20.0054, 20.00542, 20.00544, 20.00546, 20.00546, 20.00547, 
    20.00548, 20.00549, 20.00549, 20.00549, 20.00547, 20.00548, 20.00546, 
    20.00546, 20.0054, 20.00538, 20.00537, 20.00536, 20.00534, 20.00535, 
    20.00535, 20.00536, 20.00537, 20.00537, 20.00539, 20.00538, 20.00544, 
    20.00541, 20.00547, 20.00546, 20.00548, 20.00547, 20.00549, 20.00547, 
    20.0055, 20.0055, 20.0055, 20.00551, 20.00547, 20.00549, 20.00537, 
    20.00537, 20.00537, 20.00536, 20.00536, 20.00534, 20.00535, 20.00536, 
    20.00537, 20.00538, 20.00539, 20.0054, 20.00542, 20.00544, 20.00546, 
    20.00547, 20.00547, 20.00547, 20.00546, 20.00546, 20.0055, 20.00548, 
    20.00551, 20.00551, 20.00549, 20.00551, 20.00537, 20.00536, 20.00535, 
    20.00536, 20.00534, 20.00535, 20.00536, 20.00538, 20.00539, 20.00539, 
    20.0054, 20.00542, 20.00544, 20.00546, 20.00548, 20.00547, 20.00548, 
    20.00548, 20.00547, 20.00548, 20.00548, 20.00548, 20.00551, 20.0055, 
    20.00551, 20.0055, 20.00537, 20.00537, 20.00537, 20.00537, 20.00537, 
    20.00539, 20.0054, 20.00543, 20.00542, 20.00544, 20.00542, 20.00542, 
    20.00544, 20.00542, 20.00546, 20.00543, 20.00548, 20.00545, 20.00548, 
    20.00548, 20.00548, 20.00549, 20.0055, 20.00552, 20.00551, 20.00553, 
    20.00538, 20.00539, 20.00539, 20.0054, 20.00541, 20.00542, 20.00545, 
    20.00544, 20.00545, 20.00546, 20.00543, 20.00545, 20.0054, 20.00541, 
    20.0054, 20.00538, 20.00544, 20.00541, 20.00546, 20.00545, 20.00549, 
    20.00547, 20.00551, 20.00553, 20.00555, 20.00557, 20.0054, 20.00539, 
    20.0054, 20.00541, 20.00543, 20.00545, 20.00545, 20.00545, 20.00546, 
    20.00547, 20.00545, 20.00547, 20.00541, 20.00544, 20.00539, 20.0054, 
    20.00541, 20.00541, 20.00543, 20.00544, 20.00546, 20.00545, 20.00553, 
    20.00549, 20.00558, 20.00556, 20.00539, 20.0054, 20.00542, 20.00541, 
    20.00545, 20.00546, 20.00546, 20.00548, 20.00548, 20.00548, 20.00547, 
    20.00548, 20.00545, 20.00546, 20.00542, 20.00543, 20.00543, 20.00542, 
    20.00544, 20.00545, 20.00546, 20.00546, 20.00547, 20.00545, 20.00553, 
    20.00548, 20.0054, 20.00542, 20.00542, 20.00542, 20.00546, 20.00544, 
    20.00548, 20.00547, 20.00549, 20.00548, 20.00548, 20.00547, 20.00546, 
    20.00544, 20.00543, 20.00542, 20.00542, 20.00543, 20.00546, 20.00548, 
    20.00547, 20.00549, 20.00545, 20.00546, 20.00546, 20.00547, 20.00544, 
    20.00547, 20.00543, 20.00543, 20.00544, 20.00546, 20.00547, 20.00547, 
    20.00547, 20.00546, 20.00545, 20.00544, 20.00544, 20.00543, 20.00542, 
    20.00543, 20.00544, 20.00546, 20.00547, 20.00549, 20.0055, 20.00552, 
    20.0055, 20.00553, 20.0055, 20.00555, 20.00547, 20.0055, 20.00544, 
    20.00545, 20.00546, 20.00549, 20.00547, 20.00549, 20.00545, 20.00543, 
    20.00543, 20.00542, 20.00543, 20.00543, 20.00544, 20.00543, 20.00546, 
    20.00544, 20.00548, 20.00549, 20.00553, 20.00555, 20.00557, 20.00558, 
    20.00558, 20.00558,
  20.00503, 20.00505, 20.00505, 20.00507, 20.00506, 20.00507, 20.00504, 
    20.00505, 20.00504, 20.00503, 20.0051, 20.00507, 20.00514, 20.00512, 
    20.00517, 20.00513, 20.00518, 20.00517, 20.00519, 20.00519, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00522, 20.0052, 20.00507, 20.0051, 
    20.00507, 20.00508, 20.00508, 20.00506, 20.00505, 20.00503, 20.00503, 
    20.00505, 20.00508, 20.00507, 20.00509, 20.00509, 20.00512, 20.00511, 
    20.00516, 20.00515, 20.00519, 20.00518, 20.00519, 20.00518, 20.00519, 
    20.00517, 20.00518, 20.00517, 20.00511, 20.00513, 20.00508, 20.00505, 
    20.00504, 20.00502, 20.00503, 20.00503, 20.00505, 20.00506, 20.00508, 
    20.00508, 20.00509, 20.00512, 20.00513, 20.00516, 20.00516, 20.00517, 
    20.00517, 20.00519, 20.00519, 20.00519, 20.00517, 20.00518, 20.00515, 
    20.00516, 20.0051, 20.00507, 20.00506, 20.00505, 20.00503, 20.00504, 
    20.00504, 20.00505, 20.00506, 20.00506, 20.00508, 20.00507, 20.00513, 
    20.00511, 20.00517, 20.00516, 20.00518, 20.00517, 20.00519, 20.00517, 
    20.0052, 20.0052, 20.0052, 20.00521, 20.00517, 20.00519, 20.00506, 
    20.00506, 20.00506, 20.00504, 20.00504, 20.00503, 20.00504, 20.00505, 
    20.00506, 20.00507, 20.00508, 20.00509, 20.00511, 20.00514, 20.00516, 
    20.00517, 20.00517, 20.00517, 20.00516, 20.00516, 20.0052, 20.00518, 
    20.00521, 20.00521, 20.00519, 20.00521, 20.00506, 20.00505, 20.00504, 
    20.00505, 20.00503, 20.00504, 20.00505, 20.00507, 20.00508, 20.00508, 
    20.0051, 20.00511, 20.00513, 20.00516, 20.00518, 20.00517, 20.00517, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00518, 20.00521, 20.0052, 
    20.00521, 20.0052, 20.00505, 20.00506, 20.00506, 20.00507, 20.00506, 
    20.00508, 20.00509, 20.00512, 20.00511, 20.00513, 20.00511, 20.00512, 
    20.00513, 20.00511, 20.00516, 20.00513, 20.00518, 20.00515, 20.00518, 
    20.00518, 20.00518, 20.00519, 20.0052, 20.00522, 20.00522, 20.00523, 
    20.00507, 20.00508, 20.00508, 20.00509, 20.0051, 20.00512, 20.00514, 
    20.00513, 20.00515, 20.00515, 20.00513, 20.00514, 20.00509, 20.0051, 
    20.00509, 20.00507, 20.00513, 20.0051, 20.00516, 20.00514, 20.00519, 
    20.00517, 20.00521, 20.00524, 20.00525, 20.00528, 20.00509, 20.00508, 
    20.00509, 20.00511, 20.00512, 20.00514, 20.00515, 20.00515, 20.00516, 
    20.00517, 20.00515, 20.00517, 20.0051, 20.00514, 20.00508, 20.0051, 
    20.00511, 20.0051, 20.00513, 20.00514, 20.00516, 20.00515, 20.00523, 
    20.0052, 20.00529, 20.00527, 20.00508, 20.00509, 20.00512, 20.0051, 
    20.00515, 20.00516, 20.00516, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00518, 20.00514, 20.00516, 20.00512, 20.00513, 20.00512, 20.00512, 
    20.00513, 20.00515, 20.00515, 20.00516, 20.00517, 20.00515, 20.00524, 
    20.00518, 20.0051, 20.00511, 20.00512, 20.00511, 20.00516, 20.00514, 
    20.00518, 20.00517, 20.00519, 20.00518, 20.00518, 20.00517, 20.00516, 
    20.00514, 20.00512, 20.00511, 20.00511, 20.00513, 20.00515, 20.00518, 
    20.00517, 20.00519, 20.00514, 20.00516, 20.00515, 20.00517, 20.00513, 
    20.00517, 20.00512, 20.00513, 20.00514, 20.00516, 20.00517, 20.00517, 
    20.00517, 20.00515, 20.00515, 20.00514, 20.00513, 20.00513, 20.00512, 
    20.00513, 20.00513, 20.00515, 20.00517, 20.00519, 20.0052, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00526, 20.00517, 20.00521, 20.00514, 
    20.00515, 20.00516, 20.00519, 20.00517, 20.00519, 20.00515, 20.00513, 
    20.00512, 20.00511, 20.00512, 20.00512, 20.00513, 20.00513, 20.00515, 
    20.00514, 20.00518, 20.00519, 20.00523, 20.00526, 20.00528, 20.00529, 
    20.00529, 20.00529,
  20.00479, 20.00481, 20.00481, 20.00483, 20.00482, 20.00483, 20.0048, 
    20.00481, 20.0048, 20.00479, 20.00486, 20.00483, 20.0049, 20.00488, 
    20.00493, 20.0049, 20.00494, 20.00493, 20.00496, 20.00495, 20.00498, 
    20.00496, 20.005, 20.00498, 20.00498, 20.00496, 20.00484, 20.00486, 
    20.00484, 20.00484, 20.00484, 20.00482, 20.00481, 20.00479, 20.00479, 
    20.00481, 20.00484, 20.00483, 20.00486, 20.00485, 20.00488, 20.00487, 
    20.00492, 20.00491, 20.00495, 20.00494, 20.00495, 20.00495, 20.00495, 
    20.00493, 20.00494, 20.00493, 20.00488, 20.00489, 20.00484, 20.00482, 
    20.0048, 20.00478, 20.00479, 20.00479, 20.00481, 20.00482, 20.00484, 
    20.00485, 20.00485, 20.00488, 20.00489, 20.00493, 20.00492, 20.00493, 
    20.00494, 20.00495, 20.00495, 20.00496, 20.00493, 20.00495, 20.00492, 
    20.00493, 20.00486, 20.00483, 20.00482, 20.00481, 20.00479, 20.0048, 
    20.0048, 20.00481, 20.00482, 20.00482, 20.00485, 20.00484, 20.0049, 
    20.00487, 20.00494, 20.00492, 20.00494, 20.00493, 20.00495, 20.00493, 
    20.00496, 20.00497, 20.00496, 20.00498, 20.00493, 20.00495, 20.00482, 
    20.00482, 20.00482, 20.0048, 20.0048, 20.00479, 20.0048, 20.00481, 
    20.00482, 20.00483, 20.00484, 20.00486, 20.00488, 20.0049, 20.00492, 
    20.00494, 20.00493, 20.00493, 20.00493, 20.00492, 20.00496, 20.00494, 
    20.00498, 20.00497, 20.00496, 20.00497, 20.00482, 20.00481, 20.0048, 
    20.00481, 20.00479, 20.0048, 20.00481, 20.00484, 20.00484, 20.00485, 
    20.00486, 20.00487, 20.0049, 20.00492, 20.00494, 20.00494, 20.00494, 
    20.00494, 20.00493, 20.00494, 20.00495, 20.00494, 20.00497, 20.00496, 
    20.00497, 20.00497, 20.00481, 20.00482, 20.00482, 20.00483, 20.00482, 
    20.00484, 20.00485, 20.00489, 20.00487, 20.00489, 20.00488, 20.00488, 
    20.00489, 20.00488, 20.00492, 20.00489, 20.00494, 20.00491, 20.00495, 
    20.00494, 20.00495, 20.00496, 20.00497, 20.00499, 20.00498, 20.005, 
    20.00483, 20.00484, 20.00484, 20.00485, 20.00486, 20.00488, 20.0049, 
    20.00489, 20.00491, 20.00492, 20.00489, 20.00491, 20.00485, 20.00486, 
    20.00485, 20.00484, 20.0049, 20.00486, 20.00492, 20.00491, 20.00496, 
    20.00493, 20.00498, 20.005, 20.00502, 20.00504, 20.00485, 20.00484, 
    20.00485, 20.00487, 20.00489, 20.00491, 20.00491, 20.00491, 20.00492, 
    20.00493, 20.00491, 20.00493, 20.00486, 20.0049, 20.00484, 20.00486, 
    20.00487, 20.00486, 20.00489, 20.0049, 20.00493, 20.00491, 20.005, 
    20.00496, 20.00506, 20.00503, 20.00484, 20.00485, 20.00488, 20.00487, 
    20.00491, 20.00492, 20.00493, 20.00494, 20.00494, 20.00495, 20.00493, 
    20.00495, 20.00491, 20.00492, 20.00488, 20.00489, 20.00488, 20.00488, 
    20.00489, 20.00491, 20.00492, 20.00492, 20.00494, 20.00491, 20.005, 
    20.00494, 20.00486, 20.00488, 20.00488, 20.00487, 20.00492, 20.0049, 
    20.00495, 20.00493, 20.00495, 20.00494, 20.00494, 20.00493, 20.00492, 
    20.0049, 20.00489, 20.00487, 20.00488, 20.00489, 20.00492, 20.00494, 
    20.00493, 20.00495, 20.00491, 20.00492, 20.00492, 20.00494, 20.00489, 
    20.00493, 20.00488, 20.00489, 20.0049, 20.00493, 20.00493, 20.00494, 
    20.00493, 20.00492, 20.00491, 20.0049, 20.0049, 20.00489, 20.00488, 
    20.00489, 20.00489, 20.00492, 20.00494, 20.00496, 20.00496, 20.00499, 
    20.00497, 20.005, 20.00497, 20.00502, 20.00493, 20.00497, 20.0049, 
    20.00491, 20.00492, 20.00495, 20.00494, 20.00496, 20.00491, 20.00489, 
    20.00488, 20.00487, 20.00488, 20.00488, 20.00489, 20.00489, 20.00492, 
    20.0049, 20.00494, 20.00496, 20.005, 20.00502, 20.00505, 20.00506, 
    20.00506, 20.00506,
  20.00426, 20.00427, 20.00427, 20.00429, 20.00428, 20.00429, 20.00426, 
    20.00428, 20.00426, 20.00426, 20.00432, 20.00429, 20.00435, 20.00433, 
    20.00438, 20.00435, 20.00438, 20.00438, 20.0044, 20.00439, 20.00442, 
    20.0044, 20.00444, 20.00442, 20.00442, 20.0044, 20.00429, 20.00431, 
    20.00429, 20.0043, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00427, 20.0043, 20.00429, 20.00431, 20.00431, 20.00434, 20.00433, 
    20.00437, 20.00436, 20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 
    20.00438, 20.00439, 20.00437, 20.00433, 20.00434, 20.0043, 20.00428, 
    20.00426, 20.00425, 20.00425, 20.00425, 20.00427, 20.00428, 20.0043, 
    20.0043, 20.00431, 20.00433, 20.00434, 20.00437, 20.00437, 20.00438, 
    20.00438, 20.0044, 20.00439, 20.0044, 20.00438, 20.00439, 20.00437, 
    20.00437, 20.00431, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00426, 20.00427, 20.00428, 20.00428, 20.0043, 20.00429, 20.00435, 
    20.00432, 20.00438, 20.00437, 20.00439, 20.00438, 20.00439, 20.00438, 
    20.0044, 20.00441, 20.00441, 20.00442, 20.00438, 20.00439, 20.00428, 
    20.00428, 20.00428, 20.00427, 20.00427, 20.00425, 20.00426, 20.00427, 
    20.00428, 20.00429, 20.0043, 20.00431, 20.00433, 20.00435, 20.00437, 
    20.00438, 20.00437, 20.00438, 20.00437, 20.00437, 20.00441, 20.00439, 
    20.00442, 20.00442, 20.0044, 20.00442, 20.00428, 20.00427, 20.00426, 
    20.00427, 20.00425, 20.00426, 20.00427, 20.00429, 20.0043, 20.0043, 
    20.00431, 20.00433, 20.00435, 20.00437, 20.00438, 20.00438, 20.00438, 
    20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 20.00442, 20.00441, 
    20.00442, 20.00441, 20.00428, 20.00428, 20.00428, 20.00429, 20.00428, 
    20.0043, 20.00431, 20.00434, 20.00433, 20.00434, 20.00433, 20.00433, 
    20.00434, 20.00433, 20.00437, 20.00434, 20.00439, 20.00436, 20.00439, 
    20.00438, 20.00439, 20.0044, 20.00441, 20.00443, 20.00442, 20.00444, 
    20.00429, 20.0043, 20.0043, 20.00431, 20.00432, 20.00433, 20.00435, 
    20.00434, 20.00436, 20.00436, 20.00434, 20.00435, 20.00431, 20.00431, 
    20.00431, 20.00429, 20.00435, 20.00432, 20.00437, 20.00435, 20.0044, 
    20.00438, 20.00442, 20.00444, 20.00446, 20.00447, 20.0043, 20.0043, 
    20.00431, 20.00432, 20.00434, 20.00436, 20.00436, 20.00436, 20.00437, 
    20.00438, 20.00436, 20.00438, 20.00432, 20.00435, 20.0043, 20.00431, 
    20.00432, 20.00432, 20.00434, 20.00435, 20.00437, 20.00436, 20.00443, 
    20.0044, 20.00449, 20.00447, 20.0043, 20.0043, 20.00433, 20.00432, 
    20.00436, 20.00437, 20.00437, 20.00438, 20.00438, 20.00439, 20.00438, 
    20.00439, 20.00436, 20.00437, 20.00433, 20.00434, 20.00434, 20.00433, 
    20.00435, 20.00436, 20.00436, 20.00437, 20.00438, 20.00436, 20.00444, 
    20.00439, 20.00431, 20.00433, 20.00433, 20.00433, 20.00437, 20.00435, 
    20.00439, 20.00438, 20.0044, 20.00439, 20.00439, 20.00438, 20.00437, 
    20.00435, 20.00434, 20.00433, 20.00433, 20.00434, 20.00436, 20.00438, 
    20.00438, 20.0044, 20.00435, 20.00437, 20.00437, 20.00438, 20.00434, 
    20.00438, 20.00434, 20.00434, 20.00435, 20.00437, 20.00438, 20.00438, 
    20.00438, 20.00436, 20.00436, 20.00435, 20.00435, 20.00434, 20.00433, 
    20.00434, 20.00434, 20.00436, 20.00438, 20.0044, 20.0044, 20.00443, 
    20.00441, 20.00444, 20.00441, 20.00446, 20.00438, 20.00441, 20.00435, 
    20.00436, 20.00437, 20.0044, 20.00438, 20.0044, 20.00436, 20.00434, 
    20.00434, 20.00433, 20.00434, 20.00434, 20.00434, 20.00434, 20.00436, 
    20.00435, 20.00439, 20.0044, 20.00443, 20.00446, 20.00448, 20.00449, 
    20.00449, 20.00449,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258142, 0.5258148, 0.5258147, 0.5258151, 0.5258149, 0.5258152, 
    0.5258144, 0.5258148, 0.5258145, 0.5258143, 0.525816, 0.5258151, 
    0.5258169, 0.5258163, 0.5258176, 0.5258168, 0.5258178, 0.5258176, 
    0.5258182, 0.525818, 0.5258189, 0.5258183, 0.5258192, 0.5258187, 
    0.5258188, 0.5258183, 0.5258153, 0.5258159, 0.5258153, 0.5258154, 
    0.5258153, 0.5258149, 0.5258147, 0.5258142, 0.5258143, 0.5258147, 
    0.5258154, 0.5258151, 0.5258158, 0.5258158, 0.5258165, 0.5258162, 
    0.5258174, 0.5258171, 0.5258181, 0.5258178, 0.525818, 0.525818, 0.525818, 
    0.5258177, 0.5258179, 0.5258175, 0.5258163, 0.5258166, 0.5258155, 
    0.5258148, 0.5258144, 0.5258141, 0.5258141, 0.5258142, 0.5258147, 
    0.5258151, 0.5258154, 0.5258155, 0.5258158, 0.5258164, 0.5258167, 
    0.5258175, 0.5258173, 0.5258176, 0.5258178, 0.5258182, 0.5258181, 
    0.5258183, 0.5258176, 0.525818, 0.5258173, 0.5258175, 0.5258158, 
    0.5258152, 0.525815, 0.5258147, 0.5258141, 0.5258145, 0.5258144, 
    0.5258148, 0.525815, 0.5258149, 0.5258156, 0.5258153, 0.5258167, 
    0.5258161, 0.5258178, 0.5258174, 0.5258179, 0.5258176, 0.525818, 
    0.5258176, 0.5258183, 0.5258185, 0.5258183, 0.5258188, 0.5258176, 
    0.525818, 0.5258148, 0.5258149, 0.525815, 0.5258146, 0.5258145, 
    0.5258142, 0.5258145, 0.5258147, 0.525815, 0.5258152, 0.5258154, 
    0.5258158, 0.5258163, 0.5258169, 0.5258174, 0.5258178, 0.5258175, 
    0.5258177, 0.5258175, 0.5258174, 0.5258184, 0.5258179, 0.5258187, 
    0.5258186, 0.5258183, 0.5258186, 0.5258149, 0.5258148, 0.5258144, 
    0.5258147, 0.5258142, 0.5258145, 0.5258147, 0.5258153, 0.5258154, 
    0.5258156, 0.5258158, 0.5258162, 0.5258168, 0.5258173, 0.5258178, 
    0.5258178, 0.5258178, 0.5258179, 0.5258176, 0.5258179, 0.525818, 
    0.5258179, 0.5258186, 0.5258184, 0.5258186, 0.5258185, 0.5258148, 
    0.525815, 0.5258149, 0.5258151, 0.525815, 0.5258155, 0.5258157, 
    0.5258165, 0.5258162, 0.5258167, 0.5258163, 0.5258163, 0.5258167, 
    0.5258163, 0.5258173, 0.5258166, 0.5258179, 0.5258172, 0.5258179, 
    0.5258178, 0.525818, 0.5258182, 0.5258185, 0.5258189, 0.5258188, 
    0.5258192, 0.5258152, 0.5258155, 0.5258155, 0.5258157, 0.5258159, 
    0.5258163, 0.525817, 0.5258167, 0.5258172, 0.5258172, 0.5258166, 
    0.525817, 0.5258157, 0.5258159, 0.5258157, 0.5258153, 0.5258168, 
    0.525816, 0.5258174, 0.525817, 0.5258182, 0.5258176, 0.5258188, 
    0.5258193, 0.5258198, 0.5258203, 0.5258157, 0.5258155, 0.5258158, 
    0.5258161, 0.5258166, 0.525817, 0.5258171, 0.5258172, 0.5258174, 
    0.5258176, 0.5258172, 0.5258176, 0.5258159, 0.5258169, 0.5258154, 
    0.5258158, 0.5258161, 0.525816, 0.5258167, 0.5258169, 0.5258175, 
    0.5258172, 0.5258192, 0.5258183, 0.5258207, 0.52582, 0.5258154, 
    0.5258157, 0.5258164, 0.525816, 0.525817, 0.5258173, 0.5258175, 
    0.5258178, 0.5258178, 0.525818, 0.5258177, 0.5258179, 0.525817, 
    0.5258175, 0.5258163, 0.5258166, 0.5258164, 0.5258163, 0.5258167, 
    0.5258172, 0.5258172, 0.5258173, 0.5258178, 0.525817, 0.5258192, 
    0.5258179, 0.5258159, 0.5258163, 0.5258164, 0.5258162, 0.5258173, 
    0.5258169, 0.525818, 0.5258177, 0.5258182, 0.5258179, 0.5258179, 
    0.5258176, 0.5258174, 0.5258169, 0.5258165, 0.5258162, 0.5258163, 
    0.5258166, 0.5258172, 0.5258178, 0.5258177, 0.5258181, 0.525817, 
    0.5258175, 0.5258173, 0.5258178, 0.5258167, 0.5258176, 0.5258165, 
    0.5258166, 0.5258169, 0.5258175, 0.5258176, 0.5258178, 0.5258177, 
    0.5258173, 0.5258172, 0.5258169, 0.5258168, 0.5258166, 0.5258164, 
    0.5258166, 0.5258167, 0.5258173, 0.5258177, 0.5258182, 0.5258183, 
    0.5258189, 0.5258185, 0.5258193, 0.5258186, 0.5258198, 0.5258176, 
    0.5258186, 0.5258169, 0.5258171, 0.5258174, 0.5258182, 0.5258178, 
    0.5258182, 0.5258172, 0.5258166, 0.5258165, 0.5258163, 0.5258165, 
    0.5258165, 0.5258167, 0.5258167, 0.5258173, 0.5258169, 0.5258179, 
    0.5258182, 0.5258192, 0.5258198, 0.5258204, 0.5258207, 0.5258207, 
    0.5258208 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -2.569961e-21, -7.709882e-21, -5.139921e-21, 0, -2.569961e-21, 
    -1.027984e-20, -1.28498e-20, 7.709882e-21, 2.055969e-20, -5.139921e-21, 
    5.139921e-21, -1.798972e-20, 2.569961e-21, -2.055969e-20, -7.709882e-21, 
    1.027984e-20, 7.709882e-21, 1.28498e-20, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    0, 2.569961e-21, 0, 5.139921e-21, -2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -1.798972e-20, -2.826957e-20, -2.569961e-21, 1.28498e-20, 
    -1.003089e-36, -5.139921e-21, 2.055969e-20, 1.28498e-20, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    2.055969e-20, 2.569961e-21, -1.28498e-20, 1.28498e-20, 2.312965e-20, 
    2.569961e-21, -2.569961e-21, 1.541976e-20, -1.798972e-20, 7.709882e-21, 
    1.027984e-20, 1.798972e-20, -1.798972e-20, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 2.569961e-21, -1.28498e-20, 
    7.709882e-21, -1.28498e-20, 1.027984e-20, 7.709882e-21, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, 1.003089e-36, 1.003089e-36, 5.139921e-21, 
    7.709882e-21, 0, -1.798972e-20, 0, -1.28498e-20, 2.569961e-21, 
    -1.027984e-20, -1.28498e-20, 5.139921e-21, -1.027984e-20, -1.798972e-20, 
    2.569961e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, 1.798972e-20, 
    -1.027984e-20, 1.027984e-20, 1.28498e-20, 1.003089e-36, 1.798972e-20, 
    -5.015443e-37, -1.003089e-36, -1.003089e-36, -7.709882e-21, 
    -2.569961e-21, -1.28498e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, -2.055969e-20, 
    2.569961e-21, 2.055969e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    2.569961e-20, -5.139921e-21, -1.28498e-20, -1.027984e-20, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, -1.003089e-36, -1.541976e-20, -1.027984e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, 
    1.003089e-36, -7.709882e-21, -1.28498e-20, 2.569961e-21, -1.798972e-20, 
    -5.139921e-21, -1.28498e-20, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -1.003089e-36, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    1.28498e-20, -2.569961e-21, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, -2.055969e-20, 1.003089e-36, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, -1.541976e-20, 7.709882e-21, 
    0, 1.027984e-20, 1.541976e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 0, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, 5.139921e-21, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, 7.709882e-21, -1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -7.709882e-21, -1.003089e-36, 
    -2.569961e-21, 5.139921e-21, -1.541976e-20, 1.003089e-36, -1.28498e-20, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -1.28498e-20, -1.798972e-20, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -1.798972e-20, 7.709882e-21, 2.569961e-21, 1.027984e-20, -1.003089e-36, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -2.055969e-20, 2.569961e-21, -1.541976e-20, 
    -1.003089e-36, -2.569961e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    1.798972e-20, 1.28498e-20, 0, -2.055969e-20, 0, 1.28498e-20, 
    1.541976e-20, -1.027984e-20, 1.003089e-36, 2.569961e-21, 7.709882e-21, 0, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, 1.28498e-20, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, -2.312965e-20, -1.003089e-36, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -1.28498e-20, 7.709882e-21, 0, 5.139921e-21, 
    1.798972e-20, 5.139921e-21, -2.569961e-21, 1.003089e-36, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, 
    1.003089e-36, -1.027984e-20, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    1.003089e-36, 5.139921e-21, -1.003089e-36, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, 5.139921e-21, 1.003089e-36, 1.541976e-20, 
    -1.003089e-36, -5.139921e-21, -5.139921e-21, 2.312965e-20, -3.083953e-20, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -1.28498e-20, -2.569961e-21, -3.009266e-36, 1.003089e-36, 2.569961e-21, 
    1.28498e-20, -1.003089e-36, 1.027984e-20, -7.709882e-21, 2.569961e-21, 
    -1.28498e-20, -5.139921e-21, -2.569961e-21, 1.027984e-20, -1.003089e-36, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, -2.055969e-20, 2.569961e-21, 
    -2.569961e-21, 1.541976e-20, 1.28498e-20, 1.027984e-20, 2.569961e-21, 
    -1.28498e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -1.798972e-20, 2.569961e-21, 7.709882e-21,
  1.28498e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.28498e-20, -1.027984e-20, 5.139921e-21, -1.798972e-20, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.003089e-36, 7.709882e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -7.709882e-21, 1.027984e-20, 1.541976e-20, -1.003089e-36, 
    -1.28498e-20, 2.569961e-21, -5.139921e-21, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, -1.027984e-20, 2.312965e-20, 1.28498e-20, 
    -7.709882e-21, -2.055969e-20, 1.28498e-20, 5.139921e-21, -1.28498e-20, 
    -1.027984e-20, -1.003089e-36, -5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 0, 2.569961e-21, -1.003089e-36, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 0, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, 0, 5.139921e-21, -2.569961e-21, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -1.28498e-20, -5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, 0, -1.027984e-20, 
    2.569961e-21, 0, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -1.798972e-20, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 0, 
    -7.709882e-21, -5.139921e-21, 1.798972e-20, -7.709882e-21, -2.569961e-21, 
    0, 0, 0, 1.28498e-20, 2.569961e-21, -2.569961e-21, -1.541976e-20, 
    1.003089e-36, 7.709882e-21, 0, 5.139921e-21, 1.541976e-20, 0, 
    -1.003089e-36, -1.798972e-20, 1.28498e-20, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, 
    2.055969e-20, -7.709882e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, 7.709882e-21, 0, 2.055969e-20, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -7.709882e-21, -1.541976e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 0, 
    5.139921e-21, 0, 5.139921e-21, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, -7.709882e-21, 
    1.003089e-36, 0, 2.569961e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, 7.709882e-21, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -1.28498e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 7.709882e-21, -7.709882e-21, -5.139921e-21, 
    0, -5.139921e-21, -1.28498e-20, -1.003089e-36, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.541976e-20, -1.003089e-36, 
    -2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, -1.027984e-20, 
    -2.569961e-21, -1.003089e-36, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 1.28498e-20, -1.28498e-20, 7.709882e-21, 
    1.28498e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.003089e-36, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, 0, 2.569961e-21, 
    -2.569961e-21, 1.28498e-20, 7.709882e-21, 0, 0, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 0, 7.709882e-21, -7.709882e-21, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, 2.569961e-21, 1.541976e-20, -5.139921e-21, -1.28498e-20, 0, 
    1.28498e-20, 0, 5.139921e-21, 2.569961e-21, 2.569961e-21, 1.003089e-36, 
    -2.569961e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 0, 7.709882e-21, 0, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 1.541976e-20, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, 1.003089e-36, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    1.28498e-20, -2.569961e-21, -2.569961e-21, 7.709882e-21, 1.28498e-20, 0, 
    -1.28498e-20, 7.709882e-21, 0, 7.709882e-21, 2.569961e-21, 0, 0, 
    -1.003089e-36, 0,
  1.28498e-20, 7.709882e-21, -7.709882e-21, 1.003089e-36, -1.027984e-20, 
    -1.798972e-20, 5.139921e-21, -5.139921e-21, 0, 7.709882e-21, 
    1.003089e-36, -1.027984e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -1.28498e-20, 0, 1.003089e-36, -1.027984e-20, 1.003089e-36, 
    -1.541976e-20, -7.709882e-21, 2.055969e-20, -2.569961e-21, -5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 0, 7.709882e-21, 1.28498e-20, -2.569961e-21, 
    2.569961e-21, 1.28498e-20, 1.28498e-20, -7.709882e-21, 2.826957e-20, 
    2.569961e-21, -1.541976e-20, 5.139921e-21, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 1.541976e-20, 
    2.569961e-21, -7.709882e-21, 0, -5.139921e-21, -2.569961e-21, 0, 0, 
    -7.709882e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, 0, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, -1.003089e-36, 0, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, -1.003089e-36, 
    -1.28498e-20, -7.709882e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, -1.28498e-20, -1.28498e-20, -5.139921e-21, 
    -1.798972e-20, 5.139921e-21, 1.027984e-20, 0, 2.569961e-21, -1.28498e-20, 
    -1.027984e-20, -2.055969e-20, 0, -7.709882e-21, -1.798972e-20, 0, 
    -1.798972e-20, -7.709882e-21, -7.709882e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 1.027984e-20, 5.139921e-21, 7.709882e-21, 7.709882e-21, 
    7.709882e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, 1.798972e-20, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, 7.709882e-21, 1.798972e-20, 
    -2.569961e-21, 2.569961e-21, 0, 5.139921e-21, 1.003089e-36, 2.569961e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 1.003089e-36, 
    1.027984e-20, -7.709882e-21, 0, -1.798972e-20, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 7.709882e-21, -5.139921e-21, 1.28498e-20, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    1.027984e-20, -2.569961e-21, -2.055969e-20, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, -2.826957e-20, 0, 1.003089e-36, 2.569961e-21, 1.003089e-36, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, 2.569961e-21, 0, 
    -5.139921e-21, 1.027984e-20, -1.798972e-20, 7.709882e-21, 1.027984e-20, 
    1.003089e-36, 2.569961e-21, 2.055969e-20, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -7.709882e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    1.28498e-20, -7.709882e-21, -1.541976e-20, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, -1.003089e-36, 2.569961e-21, 7.709882e-21, -7.709882e-21, 
    -1.541976e-20, 5.139921e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 
    0, -1.027984e-20, 7.709882e-21, 2.055969e-20, -5.139921e-21, 
    -5.139921e-21, 1.003089e-36, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, -2.055969e-20, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 1.027984e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 0, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -1.027984e-20, 1.541976e-20, -5.139921e-21, -2.569961e-21, 
    1.28498e-20, 0, 2.569961e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 1.003089e-36, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -1.027984e-20, -5.139921e-21, -1.28498e-20, -1.798972e-20, 
    1.798972e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, -2.055969e-20, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, 1.798972e-20, 5.139921e-21, 
    -5.139921e-21, 1.003089e-36, 1.003089e-36, 1.541976e-20, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, -2.569961e-21, 
    -1.541976e-20, -1.027984e-20, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 0, -7.709882e-21, -1.28498e-20, 
    1.541976e-20, -7.709882e-21, 1.027984e-20, -1.28498e-20, -1.28498e-20, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, 2.055969e-20, -1.28498e-20, 
    -1.28498e-20, -7.709882e-21, -2.569961e-21, 2.569961e-21, 0, 1.28498e-20, 
    -1.003089e-36, 1.027984e-20, -2.569961e-21, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, 0, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 1.003089e-36, 2.569961e-21, 7.709882e-21, -1.003089e-36, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    1.541976e-20, -5.139921e-21, 1.003089e-36, 5.139921e-21, 0, 1.541976e-20, 
    0, -2.569961e-21, 2.569961e-21, -5.139921e-21, -1.541976e-20, 
    2.569961e-21, 7.709882e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21,
  -1.003089e-36, 2.569961e-21, 7.709882e-21, 1.28498e-20, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, -1.541976e-20, 
    1.027984e-20, -1.28498e-20, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 1.28498e-20, 
    -1.28498e-20, 2.569961e-21, -1.798972e-20, -7.709882e-21, 2.055969e-20, 
    -7.709882e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 2.055969e-20, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 0, 1.28498e-20, 1.003089e-36, 1.027984e-20, 
    -1.28498e-20, -1.027984e-20, 5.139921e-21, 2.569961e-21, -2.569961e-20, 
    7.709882e-21, 1.027984e-20, -2.569961e-21, -1.798972e-20, -2.569961e-21, 
    5.139921e-21, -1.003089e-36, 1.027984e-20, 5.139921e-21, 2.055969e-20, 
    1.28498e-20, -1.027984e-20, 2.569961e-21, 1.798972e-20, 1.027984e-20, 
    1.28498e-20, 7.709882e-21, -1.28498e-20, -1.798972e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, -2.055969e-20, 
    -2.569961e-21, -1.28498e-20, 1.541976e-20, 7.709882e-21, -1.003089e-36, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    1.28498e-20, -1.003089e-36, 1.28498e-20, -1.003089e-36, 5.139921e-21, 0, 
    -1.003089e-36, 5.139921e-21, 2.055969e-20, 0, -1.28498e-20, 
    -7.709882e-21, -1.027984e-20, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    5.139921e-21, 1.003089e-36, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    1.003089e-36, -1.28498e-20, -1.003089e-36, 0, 1.541976e-20, 
    -7.709882e-21, -1.798972e-20, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 2.569961e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.798972e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    0, -7.709882e-21, 1.798972e-20, -1.798972e-20, -1.28498e-20, 
    2.569961e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, 
    1.541976e-20, -5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, -1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 0, 
    -7.709882e-21, -1.798972e-20, 1.28498e-20, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, 1.798972e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 7.709882e-21, 1.798972e-20, 1.027984e-20, 0, 
    7.709882e-21, 1.003089e-36, 7.709882e-21, 1.003089e-36, 1.003089e-36, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    -1.003089e-36, -2.569961e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, 
    2.055969e-20, -5.139921e-21, 1.798972e-20, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, 1.027984e-20, 1.027984e-20, -1.798972e-20, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 2.055969e-20, 
    1.541976e-20, 7.709882e-21, -1.003089e-36, 1.027984e-20, -1.541976e-20, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, -1.541976e-20, 0, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    7.709882e-21, 0, 1.027984e-20, -2.569961e-21, 1.28498e-20, -7.709882e-21, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, 2.569961e-21, 2.055969e-20, 
    -1.28498e-20, 5.139921e-21, 1.027984e-20, -2.569961e-21, -7.709882e-21, 
    2.055969e-20, 1.027984e-20, 2.569961e-21, 2.055969e-20, -5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -1.28498e-20, 1.798972e-20, 7.709882e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 5.139921e-21, -1.541976e-20, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 7.709882e-21, 0, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 0, 
    -1.541976e-20, 0, 1.003089e-36, -5.139921e-21, -1.027984e-20, 
    -7.709882e-21, 0, 5.139921e-21, 2.312965e-20, -1.027984e-20, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 2.055969e-20, -1.28498e-20, 
    1.003089e-36, -7.709882e-21, 5.139921e-21, 1.798972e-20, -1.28498e-20, 
    -2.055969e-20, -1.28498e-20, -1.541976e-20, 2.569961e-21, -1.541976e-20, 
    -1.003089e-36, -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    1.027984e-20, -5.139921e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, -1.541976e-20, -1.541976e-20, 2.569961e-21, -1.027984e-20, 
    1.027984e-20, -1.798972e-20, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 0, -1.541976e-20, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, -1.798972e-20, 
    -1.798972e-20, 1.027984e-20, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 1.541976e-20, 7.709882e-21, -2.569961e-21, 
    -1.003089e-36, -1.28498e-20, 7.709882e-21, -2.569961e-21, -1.003089e-36, 
    1.541976e-20, 5.139921e-21, 1.28498e-20, -1.28498e-20, 5.139921e-21, 
    7.709882e-21,
  -2.569961e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 1.28498e-20, 
    7.709882e-21, -1.003089e-36, 1.28498e-20, -1.003089e-36, -1.003089e-36, 
    -1.798972e-20, 2.569961e-21, -7.709882e-21, 0, 5.139921e-21, 
    -1.541976e-20, 2.569961e-20, 7.709882e-21, 2.569961e-21, 1.798972e-20, 
    2.569961e-21, -1.798972e-20, 2.569961e-21, -1.798972e-20, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, -2.312965e-20, 
    -1.027984e-20, -7.709882e-21, -7.709882e-21, 1.28498e-20, -2.055969e-20, 
    7.709882e-21, 1.003089e-36, 1.027984e-20, 1.003089e-36, -1.003089e-36, 
    1.28498e-20, 2.569961e-20, -2.569961e-21, 0, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 0, -1.027984e-20, 2.569961e-21, 0, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, 1.003089e-36, 1.541976e-20, -2.569961e-21, 
    -5.139921e-21, -2.312965e-20, 2.569961e-21, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 2.312965e-20, 
    0, 7.709882e-21, 1.28498e-20, 5.139921e-21, 1.027984e-20, -2.569961e-21, 
    2.569961e-20, -1.027984e-20, -5.139921e-21, -7.709882e-21, -1.541976e-20, 
    0, 1.027984e-20, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.28498e-20, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, 0, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, 0, 2.312965e-20, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -2.569961e-21, -7.709882e-21, -2.569961e-21, 2.055969e-20, 
    -1.28498e-20, 2.569961e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, 
    -1.28498e-20, -5.139921e-21, -1.027984e-20, -3.083953e-20, 1.28498e-20, 
    2.569961e-21, 7.709882e-21, -5.139921e-21, -1.541976e-20, -1.003089e-36, 
    -7.709882e-21, -1.003089e-36, -1.541976e-20, 1.541976e-20, 7.709882e-21, 
    1.28498e-20, -7.709882e-21, -5.139921e-21, -1.541976e-20, -1.798972e-20, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -2.055969e-20, 1.003089e-36, -7.709882e-21, -1.003089e-36, 2.312965e-20, 
    -2.055969e-20, -2.569961e-20, 2.569961e-21, 5.139921e-21, -1.027984e-20, 
    -1.28498e-20, -1.541976e-20, 3.083953e-20, -1.541976e-20, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, -1.027984e-20, -1.798972e-20, 1.798972e-20, -7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 0, 1.28498e-20, 2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -1.28498e-20, 7.709882e-21, 7.709882e-21, 
    -2.055969e-20, 5.139921e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, -1.541976e-20, -1.28498e-20, 
    -5.139921e-21, 2.055969e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, 7.709882e-21, 
    -1.003089e-36, 7.709882e-21, 2.569961e-21, 0, 1.28498e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 1.28498e-20, 2.569961e-21, 
    -1.027984e-20, -1.003089e-36, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 3.340949e-20, 1.003089e-36, -2.569961e-20, -1.541976e-20, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, 1.28498e-20, -1.28498e-20, 
    2.569961e-21, -7.709882e-21, 1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -5.139921e-21, 5.139921e-21, -2.055969e-20, -7.709882e-21, -1.541976e-20, 
    -1.003089e-36, 1.003089e-36, 5.139921e-21, 1.003089e-36, -5.139921e-21, 
    5.139921e-21, -1.003089e-36, -7.709882e-21, -2.569961e-21, -1.798972e-20, 
    -7.709882e-21, -7.709882e-21, -1.003089e-36, -2.569961e-21, 1.798972e-20, 
    1.027984e-20, -5.139921e-21, -2.312965e-20, -5.139921e-21, -1.541976e-20, 
    1.28498e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, -1.541976e-20, 1.28498e-20, 
    1.027984e-20, 2.569961e-21, -1.798972e-20, -5.139921e-21, 1.027984e-20, 
    3.009266e-36, 1.798972e-20, 1.541976e-20, 2.569961e-21, -1.027984e-20, 
    1.027984e-20, 0, 5.139921e-21, -1.28498e-20, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, 0, -2.569961e-21, -1.28498e-20, 1.027984e-20, 
    -1.541976e-20, 1.28498e-20, 3.083953e-20, 1.798972e-20, 2.569961e-21, 
    7.709882e-21, -1.28498e-20, -1.027984e-20, 1.541976e-20, -2.569961e-21, 
    -1.027984e-20, -5.139921e-21, -1.798972e-20, 5.139921e-21, -5.139921e-21, 
    1.28498e-20, 2.055969e-20, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    2.569961e-21, 0, 5.139921e-21, 1.798972e-20, 1.003089e-36, -2.569961e-21, 
    1.28498e-20, 1.003089e-36, -1.541976e-20, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.798972e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -1.003089e-36, 1.027984e-20, -7.709882e-21, -1.027984e-20, 1.003089e-36, 
    -7.709882e-21,
  6.259378e-29, 6.259384e-29, 6.259382e-29, 6.259388e-29, 6.259385e-29, 
    6.259388e-29, 6.259379e-29, 6.259384e-29, 6.259381e-29, 6.259378e-29, 
    6.259398e-29, 6.259388e-29, 6.259407e-29, 6.259401e-29, 6.259417e-29, 
    6.259407e-29, 6.259419e-29, 6.259416e-29, 6.259423e-29, 6.259421e-29, 
    6.25943e-29, 6.259424e-29, 6.259435e-29, 6.259429e-29, 6.25943e-29, 
    6.259424e-29, 6.25939e-29, 6.259396e-29, 6.25939e-29, 6.25939e-29, 
    6.25939e-29, 6.259385e-29, 6.259382e-29, 6.259377e-29, 6.259378e-29, 
    6.259382e-29, 6.259391e-29, 6.259388e-29, 6.259395e-29, 6.259395e-29, 
    6.259404e-29, 6.2594e-29, 6.259414e-29, 6.25941e-29, 6.259422e-29, 
    6.259419e-29, 6.259421e-29, 6.25942e-29, 6.259421e-29, 6.259417e-29, 
    6.259419e-29, 6.259415e-29, 6.259401e-29, 6.259405e-29, 6.259392e-29, 
    6.259384e-29, 6.259379e-29, 6.259376e-29, 6.259376e-29, 6.259377e-29, 
    6.259382e-29, 6.259387e-29, 6.25939e-29, 6.259393e-29, 6.259395e-29, 
    6.259402e-29, 6.259406e-29, 6.259414e-29, 6.259413e-29, 6.259416e-29, 
    6.259418e-29, 6.259422e-29, 6.259422e-29, 6.259423e-29, 6.259416e-29, 
    6.259421e-29, 6.259412e-29, 6.259414e-29, 6.259396e-29, 6.259388e-29, 
    6.259385e-29, 6.259383e-29, 6.259376e-29, 6.259381e-29, 6.259379e-29, 
    6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259393e-29, 6.25939e-29, 
    6.259407e-29, 6.259399e-29, 6.259418e-29, 6.259413e-29, 6.259419e-29, 
    6.259416e-29, 6.259421e-29, 6.259417e-29, 6.259424e-29, 6.259426e-29, 
    6.259425e-29, 6.259429e-29, 6.259416e-29, 6.259421e-29, 6.259385e-29, 
    6.259385e-29, 6.259386e-29, 6.259381e-29, 6.259381e-29, 6.259377e-29, 
    6.259381e-29, 6.259382e-29, 6.259386e-29, 6.259388e-29, 6.259391e-29, 
    6.259396e-29, 6.259401e-29, 6.259408e-29, 6.259414e-29, 6.259417e-29, 
    6.259415e-29, 6.259417e-29, 6.259415e-29, 6.259414e-29, 6.259425e-29, 
    6.259419e-29, 6.259428e-29, 6.259428e-29, 6.259423e-29, 6.259428e-29, 
    6.259385e-29, 6.259384e-29, 6.259379e-29, 6.259383e-29, 6.259377e-29, 
    6.25938e-29, 6.259382e-29, 6.25939e-29, 6.259391e-29, 6.259393e-29, 
    6.259396e-29, 6.2594e-29, 6.259407e-29, 6.259413e-29, 6.259419e-29, 
    6.259418e-29, 6.259418e-29, 6.259419e-29, 6.259416e-29, 6.25942e-29, 
    6.25942e-29, 6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259428e-29, 
    6.259426e-29, 6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259387e-29, 
    6.259386e-29, 6.259393e-29, 6.259394e-29, 6.259404e-29, 6.2594e-29, 
    6.259406e-29, 6.259401e-29, 6.259402e-29, 6.259406e-29, 6.259401e-29, 
    6.259413e-29, 6.259405e-29, 6.259419e-29, 6.259411e-29, 6.25942e-29, 
    6.259419e-29, 6.259421e-29, 6.259423e-29, 6.259426e-29, 6.259431e-29, 
    6.25943e-29, 6.259434e-29, 6.25939e-29, 6.259392e-29, 6.259392e-29, 
    6.259394e-29, 6.259397e-29, 6.259401e-29, 6.259408e-29, 6.259406e-29, 
    6.259411e-29, 6.259412e-29, 6.259404e-29, 6.259409e-29, 6.259394e-29, 
    6.259396e-29, 6.259395e-29, 6.25939e-29, 6.259407e-29, 6.259398e-29, 
    6.259414e-29, 6.259409e-29, 6.259423e-29, 6.259416e-29, 6.259429e-29, 
    6.259435e-29, 6.25944e-29, 6.259447e-29, 6.259393e-29, 6.259391e-29, 
    6.259395e-29, 6.259399e-29, 6.259404e-29, 6.25941e-29, 6.25941e-29, 
    6.259411e-29, 6.259414e-29, 6.259416e-29, 6.259411e-29, 6.259417e-29, 
    6.259397e-29, 6.259407e-29, 6.259391e-29, 6.259396e-29, 6.259399e-29, 
    6.259398e-29, 6.259405e-29, 6.259407e-29, 6.259415e-29, 6.259411e-29, 
    6.259434e-29, 6.259423e-29, 6.259452e-29, 6.259444e-29, 6.259391e-29, 
    6.259393e-29, 6.259402e-29, 6.259398e-29, 6.25941e-29, 6.259413e-29, 
    6.259415e-29, 6.259418e-29, 6.259419e-29, 6.25942e-29, 6.259417e-29, 
    6.25942e-29, 6.25941e-29, 6.259414e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259401e-29, 6.259406e-29, 6.259411e-29, 6.259411e-29, 
    6.259413e-29, 6.259418e-29, 6.25941e-29, 6.259435e-29, 6.259419e-29, 
    6.259396e-29, 6.259401e-29, 6.259402e-29, 6.2594e-29, 6.259413e-29, 
    6.259408e-29, 6.25942e-29, 6.259417e-29, 6.259422e-29, 6.259419e-29, 
    6.259419e-29, 6.259416e-29, 6.259413e-29, 6.259408e-29, 6.259404e-29, 
    6.2594e-29, 6.259401e-29, 6.259405e-29, 6.259412e-29, 6.259419e-29, 
    6.259417e-29, 6.259422e-29, 6.259409e-29, 6.259414e-29, 6.259412e-29, 
    6.259417e-29, 6.259406e-29, 6.259416e-29, 6.259403e-29, 6.259404e-29, 
    6.259408e-29, 6.259414e-29, 6.259416e-29, 6.259418e-29, 6.259417e-29, 
    6.259412e-29, 6.259411e-29, 6.259408e-29, 6.259407e-29, 6.259404e-29, 
    6.259402e-29, 6.259404e-29, 6.259406e-29, 6.259412e-29, 6.259417e-29, 
    6.259423e-29, 6.259425e-29, 6.259431e-29, 6.259426e-29, 6.259435e-29, 
    6.259427e-29, 6.259441e-29, 6.259416e-29, 6.259427e-29, 6.259408e-29, 
    6.25941e-29, 6.259414e-29, 6.259422e-29, 6.259417e-29, 6.259423e-29, 
    6.259411e-29, 6.259405e-29, 6.259404e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259406e-29, 6.259405e-29, 6.259412e-29, 6.259408e-29, 
    6.259419e-29, 6.259423e-29, 6.259434e-29, 6.259441e-29, 6.259447e-29, 
    6.25945e-29, 6.259452e-29, 6.259452e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.138285e-10, 2.14772e-10, 2.145886e-10, 2.153497e-10, 2.149275e-10, 
    2.154258e-10, 2.140198e-10, 2.148095e-10, 2.143054e-10, 2.139135e-10, 
    2.168265e-10, 2.153836e-10, 2.183257e-10, 2.174053e-10, 2.197175e-10, 
    2.181824e-10, 2.20027e-10, 2.196732e-10, 2.207382e-10, 2.204331e-10, 
    2.217952e-10, 2.20879e-10, 2.225014e-10, 2.215764e-10, 2.217211e-10, 
    2.208487e-10, 2.15674e-10, 2.166469e-10, 2.156164e-10, 2.157551e-10, 
    2.156929e-10, 2.149362e-10, 2.145549e-10, 2.137565e-10, 2.139014e-10, 
    2.144879e-10, 2.158175e-10, 2.153662e-10, 2.165037e-10, 2.16478e-10, 
    2.177445e-10, 2.171735e-10, 2.193023e-10, 2.186972e-10, 2.204458e-10, 
    2.20006e-10, 2.204252e-10, 2.202981e-10, 2.204268e-10, 2.197818e-10, 
    2.200582e-10, 2.194907e-10, 2.172804e-10, 2.179299e-10, 2.159928e-10, 
    2.14828e-10, 2.140545e-10, 2.135056e-10, 2.135832e-10, 2.137311e-10, 
    2.144913e-10, 2.152061e-10, 2.157509e-10, 2.161153e-10, 2.164743e-10, 
    2.175611e-10, 2.181364e-10, 2.194246e-10, 2.191922e-10, 2.19586e-10, 
    2.199623e-10, 2.20594e-10, 2.2049e-10, 2.207683e-10, 2.195756e-10, 
    2.203683e-10, 2.190598e-10, 2.194177e-10, 2.165718e-10, 2.154879e-10, 
    2.150271e-10, 2.146239e-10, 2.136428e-10, 2.143203e-10, 2.140532e-10, 
    2.146887e-10, 2.150924e-10, 2.148927e-10, 2.161252e-10, 2.156461e-10, 
    2.181705e-10, 2.170831e-10, 2.199184e-10, 2.192399e-10, 2.20081e-10, 
    2.196518e-10, 2.203873e-10, 2.197254e-10, 2.208719e-10, 2.211216e-10, 
    2.20951e-10, 2.216064e-10, 2.196887e-10, 2.204251e-10, 2.148871e-10, 
    2.149197e-10, 2.150714e-10, 2.144045e-10, 2.143637e-10, 2.137525e-10, 
    2.142963e-10, 2.145279e-10, 2.151158e-10, 2.154636e-10, 2.157942e-10, 
    2.165211e-10, 2.173329e-10, 2.184682e-10, 2.192839e-10, 2.198307e-10, 
    2.194954e-10, 2.197914e-10, 2.194605e-10, 2.193054e-10, 2.21028e-10, 
    2.200607e-10, 2.215122e-10, 2.214318e-10, 2.20775e-10, 2.214409e-10, 
    2.149426e-10, 2.147552e-10, 2.141045e-10, 2.146137e-10, 2.136859e-10, 
    2.142052e-10, 2.145038e-10, 2.15656e-10, 2.159092e-10, 2.16144e-10, 
    2.166076e-10, 2.172027e-10, 2.182466e-10, 2.191549e-10, 2.199842e-10, 
    2.199234e-10, 2.199448e-10, 2.201301e-10, 2.196712e-10, 2.202054e-10, 
    2.20295e-10, 2.200606e-10, 2.214211e-10, 2.210324e-10, 2.214301e-10, 
    2.211771e-10, 2.148161e-10, 2.151314e-10, 2.14961e-10, 2.152815e-10, 
    2.150557e-10, 2.160595e-10, 2.163605e-10, 2.17769e-10, 2.17191e-10, 
    2.181109e-10, 2.172844e-10, 2.174309e-10, 2.181409e-10, 2.173291e-10, 
    2.191048e-10, 2.179009e-10, 2.201373e-10, 2.189349e-10, 2.202126e-10, 
    2.199806e-10, 2.203648e-10, 2.207088e-10, 2.211416e-10, 2.219403e-10, 
    2.217554e-10, 2.224233e-10, 2.156016e-10, 2.160106e-10, 2.159746e-10, 
    2.164027e-10, 2.167193e-10, 2.174056e-10, 2.185062e-10, 2.180923e-10, 
    2.188522e-10, 2.190048e-10, 2.178503e-10, 2.185591e-10, 2.162844e-10, 
    2.166518e-10, 2.164331e-10, 2.156338e-10, 2.181877e-10, 2.16877e-10, 
    2.192974e-10, 2.185873e-10, 2.206597e-10, 2.19629e-10, 2.216535e-10, 
    2.22519e-10, 2.233337e-10, 2.242857e-10, 2.162339e-10, 2.15956e-10, 
    2.164536e-10, 2.171422e-10, 2.177811e-10, 2.186306e-10, 2.187175e-10, 
    2.188766e-10, 2.192889e-10, 2.196355e-10, 2.189269e-10, 2.197224e-10, 
    2.16737e-10, 2.183014e-10, 2.158509e-10, 2.165887e-10, 2.171016e-10, 
    2.168766e-10, 2.18045e-10, 2.183204e-10, 2.194395e-10, 2.18861e-10, 
    2.223054e-10, 2.207814e-10, 2.250107e-10, 2.238287e-10, 2.158588e-10, 
    2.162329e-10, 2.17535e-10, 2.169155e-10, 2.186873e-10, 2.191234e-10, 
    2.19478e-10, 2.199313e-10, 2.199802e-10, 2.202488e-10, 2.198087e-10, 
    2.202314e-10, 2.186324e-10, 2.193469e-10, 2.173862e-10, 2.178634e-10, 
    2.176439e-10, 2.174031e-10, 2.181463e-10, 2.189381e-10, 2.18955e-10, 
    2.192089e-10, 2.199243e-10, 2.186945e-10, 2.22502e-10, 2.201504e-10, 
    2.166409e-10, 2.173614e-10, 2.174644e-10, 2.171853e-10, 2.190797e-10, 
    2.183933e-10, 2.202422e-10, 2.197425e-10, 2.205613e-10, 2.201544e-10, 
    2.200946e-10, 2.19572e-10, 2.192467e-10, 2.184247e-10, 2.17756e-10, 
    2.172258e-10, 2.173491e-10, 2.179315e-10, 2.189865e-10, 2.199846e-10, 
    2.19766e-10, 2.204991e-10, 2.185588e-10, 2.193724e-10, 2.190579e-10, 
    2.198779e-10, 2.180813e-10, 2.19611e-10, 2.176903e-10, 2.178587e-10, 
    2.183796e-10, 2.194275e-10, 2.196594e-10, 2.19907e-10, 2.197542e-10, 
    2.190133e-10, 2.188919e-10, 2.18367e-10, 2.18222e-10, 2.178221e-10, 
    2.174909e-10, 2.177935e-10, 2.181112e-10, 2.190136e-10, 2.198269e-10, 
    2.207137e-10, 2.209307e-10, 2.219667e-10, 2.211233e-10, 2.225151e-10, 
    2.213317e-10, 2.233803e-10, 2.196997e-10, 2.21297e-10, 2.184034e-10, 
    2.187151e-10, 2.192789e-10, 2.205721e-10, 2.19874e-10, 2.206905e-10, 
    2.188872e-10, 2.179516e-10, 2.177096e-10, 2.17258e-10, 2.177199e-10, 
    2.176824e-10, 2.181244e-10, 2.179823e-10, 2.190436e-10, 2.184735e-10, 
    2.200931e-10, 2.206841e-10, 2.223533e-10, 2.233766e-10, 2.244184e-10, 
    2.248784e-10, 2.250184e-10, 2.250769e-10 ;

 SOIL2N_TO_SOIL3N =
  1.527347e-11, 1.534086e-11, 1.532776e-11, 1.538212e-11, 1.535197e-11, 
    1.538756e-11, 1.528713e-11, 1.534354e-11, 1.530753e-11, 1.527954e-11, 
    1.548761e-11, 1.538454e-11, 1.559469e-11, 1.552895e-11, 1.56941e-11, 
    1.558446e-11, 1.571621e-11, 1.569095e-11, 1.576701e-11, 1.574522e-11, 
    1.584251e-11, 1.577707e-11, 1.589295e-11, 1.582688e-11, 1.583722e-11, 
    1.577491e-11, 1.540529e-11, 1.547478e-11, 1.540117e-11, 1.541108e-11, 
    1.540663e-11, 1.535259e-11, 1.532535e-11, 1.526832e-11, 1.527867e-11, 
    1.532056e-11, 1.541553e-11, 1.53833e-11, 1.546455e-11, 1.546272e-11, 
    1.555318e-11, 1.551239e-11, 1.566445e-11, 1.562123e-11, 1.574613e-11, 
    1.571472e-11, 1.574465e-11, 1.573558e-11, 1.574477e-11, 1.56987e-11, 
    1.571844e-11, 1.567791e-11, 1.552003e-11, 1.556642e-11, 1.542805e-11, 
    1.534486e-11, 1.52896e-11, 1.52504e-11, 1.525594e-11, 1.526651e-11, 
    1.532081e-11, 1.537187e-11, 1.541078e-11, 1.54368e-11, 1.546245e-11, 
    1.554008e-11, 1.558117e-11, 1.567319e-11, 1.565659e-11, 1.568472e-11, 
    1.571159e-11, 1.575672e-11, 1.574929e-11, 1.576917e-11, 1.568397e-11, 
    1.574059e-11, 1.564713e-11, 1.567269e-11, 1.546941e-11, 1.539199e-11, 
    1.535908e-11, 1.533028e-11, 1.52602e-11, 1.530859e-11, 1.528952e-11, 
    1.533491e-11, 1.536374e-11, 1.534948e-11, 1.543752e-11, 1.540329e-11, 
    1.558361e-11, 1.550594e-11, 1.570846e-11, 1.565999e-11, 1.572007e-11, 
    1.568942e-11, 1.574195e-11, 1.569467e-11, 1.577657e-11, 1.57944e-11, 
    1.578221e-11, 1.582903e-11, 1.569205e-11, 1.574465e-11, 1.534908e-11, 
    1.535141e-11, 1.536225e-11, 1.53146e-11, 1.531169e-11, 1.526803e-11, 
    1.530688e-11, 1.532342e-11, 1.536542e-11, 1.539026e-11, 1.541387e-11, 
    1.546579e-11, 1.552378e-11, 1.560487e-11, 1.566314e-11, 1.570219e-11, 
    1.567824e-11, 1.569939e-11, 1.567575e-11, 1.566467e-11, 1.578772e-11, 
    1.571862e-11, 1.58223e-11, 1.581656e-11, 1.576964e-11, 1.581721e-11, 
    1.535304e-11, 1.533965e-11, 1.529318e-11, 1.532955e-11, 1.526328e-11, 
    1.530037e-11, 1.53217e-11, 1.5404e-11, 1.542209e-11, 1.543886e-11, 
    1.547197e-11, 1.551448e-11, 1.558904e-11, 1.565392e-11, 1.571316e-11, 
    1.570882e-11, 1.571034e-11, 1.572358e-11, 1.56908e-11, 1.572896e-11, 
    1.573536e-11, 1.571862e-11, 1.581579e-11, 1.578803e-11, 1.581644e-11, 
    1.579836e-11, 1.534401e-11, 1.536653e-11, 1.535436e-11, 1.537725e-11, 
    1.536112e-11, 1.543283e-11, 1.545432e-11, 1.555493e-11, 1.551364e-11, 
    1.557935e-11, 1.552032e-11, 1.553078e-11, 1.558149e-11, 1.552351e-11, 
    1.565034e-11, 1.556435e-11, 1.572409e-11, 1.56382e-11, 1.572947e-11, 
    1.57129e-11, 1.574034e-11, 1.576491e-11, 1.579583e-11, 1.585288e-11, 
    1.583967e-11, 1.588738e-11, 1.540011e-11, 1.542933e-11, 1.542676e-11, 
    1.545734e-11, 1.547995e-11, 1.552897e-11, 1.560759e-11, 1.557802e-11, 
    1.56323e-11, 1.56432e-11, 1.556074e-11, 1.561136e-11, 1.544889e-11, 
    1.547513e-11, 1.545951e-11, 1.540242e-11, 1.558483e-11, 1.549121e-11, 
    1.56641e-11, 1.561338e-11, 1.576141e-11, 1.568779e-11, 1.58324e-11, 
    1.589421e-11, 1.595241e-11, 1.602041e-11, 1.544528e-11, 1.542542e-11, 
    1.546097e-11, 1.551015e-11, 1.555579e-11, 1.561647e-11, 1.562268e-11, 
    1.563405e-11, 1.566349e-11, 1.568825e-11, 1.563764e-11, 1.569445e-11, 
    1.548122e-11, 1.559296e-11, 1.541792e-11, 1.547062e-11, 1.550726e-11, 
    1.549119e-11, 1.557465e-11, 1.559432e-11, 1.567425e-11, 1.563293e-11, 
    1.587896e-11, 1.57701e-11, 1.607219e-11, 1.598776e-11, 1.541849e-11, 
    1.544521e-11, 1.553821e-11, 1.549396e-11, 1.562052e-11, 1.565167e-11, 
    1.5677e-11, 1.570938e-11, 1.571287e-11, 1.573205e-11, 1.570062e-11, 
    1.573081e-11, 1.56166e-11, 1.566764e-11, 1.552758e-11, 1.556167e-11, 
    1.554599e-11, 1.552879e-11, 1.558188e-11, 1.563843e-11, 1.563965e-11, 
    1.565778e-11, 1.570888e-11, 1.562103e-11, 1.5893e-11, 1.572503e-11, 
    1.547435e-11, 1.552582e-11, 1.553317e-11, 1.551323e-11, 1.564855e-11, 
    1.559952e-11, 1.573159e-11, 1.569589e-11, 1.575438e-11, 1.572532e-11, 
    1.572104e-11, 1.568371e-11, 1.566048e-11, 1.560177e-11, 1.5554e-11, 
    1.551613e-11, 1.552493e-11, 1.556654e-11, 1.564189e-11, 1.571319e-11, 
    1.569757e-11, 1.574993e-11, 1.561135e-11, 1.566946e-11, 1.564699e-11, 
    1.570556e-11, 1.557724e-11, 1.56865e-11, 1.554931e-11, 1.556134e-11, 
    1.559855e-11, 1.567339e-11, 1.568996e-11, 1.570764e-11, 1.569673e-11, 
    1.564381e-11, 1.563514e-11, 1.559764e-11, 1.558729e-11, 1.555872e-11, 
    1.553506e-11, 1.555668e-11, 1.557937e-11, 1.564383e-11, 1.570192e-11, 
    1.576526e-11, 1.578077e-11, 1.585477e-11, 1.579452e-11, 1.589393e-11, 
    1.580941e-11, 1.595573e-11, 1.569284e-11, 1.580693e-11, 1.560024e-11, 
    1.562251e-11, 1.566278e-11, 1.575515e-11, 1.570529e-11, 1.576361e-11, 
    1.56348e-11, 1.556797e-11, 1.555069e-11, 1.551843e-11, 1.555142e-11, 
    1.554874e-11, 1.558031e-11, 1.557017e-11, 1.564597e-11, 1.560525e-11, 
    1.572093e-11, 1.576315e-11, 1.588238e-11, 1.595547e-11, 1.602989e-11, 
    1.606274e-11, 1.607274e-11, 1.607692e-11 ;

 SOIL2N_vr =
  1.818719, 1.818721, 1.81872, 1.818722, 1.818721, 1.818722, 1.81872, 
    1.818721, 1.81872, 1.818719, 1.818724, 1.818722, 1.818726, 1.818725, 
    1.818728, 1.818726, 1.818729, 1.818728, 1.81873, 1.81873, 1.818732, 
    1.81873, 1.818733, 1.818731, 1.818732, 1.81873, 1.818722, 1.818724, 
    1.818722, 1.818722, 1.818722, 1.818721, 1.81872, 1.818719, 1.818719, 
    1.81872, 1.818722, 1.818722, 1.818723, 1.818723, 1.818725, 1.818725, 
    1.818728, 1.818727, 1.81873, 1.818729, 1.81873, 1.818729, 1.81873, 
    1.818729, 1.818729, 1.818728, 1.818725, 1.818726, 1.818723, 1.818721, 
    1.81872, 1.818719, 1.818719, 1.818719, 1.81872, 1.818721, 1.818722, 
    1.818723, 1.818723, 1.818725, 1.818726, 1.818728, 1.818728, 1.818728, 
    1.818729, 1.81873, 1.81873, 1.81873, 1.818728, 1.818729, 1.818727, 
    1.818728, 1.818724, 1.818722, 1.818721, 1.818721, 1.818719, 1.81872, 
    1.81872, 1.818721, 1.818721, 1.818721, 1.818723, 1.818722, 1.818726, 
    1.818724, 1.818729, 1.818728, 1.818729, 1.818728, 1.81873, 1.818728, 
    1.81873, 1.818731, 1.81873, 1.818731, 1.818728, 1.81873, 1.818721, 
    1.818721, 1.818721, 1.81872, 1.81872, 1.818719, 1.81872, 1.81872, 
    1.818721, 1.818722, 1.818722, 1.818723, 1.818725, 1.818727, 1.818728, 
    1.818729, 1.818728, 1.818729, 1.818728, 1.818728, 1.81873, 1.818729, 
    1.818731, 1.818731, 1.81873, 1.818731, 1.818721, 1.818721, 1.81872, 
    1.818721, 1.818719, 1.81872, 1.81872, 1.818722, 1.818722, 1.818723, 
    1.818724, 1.818725, 1.818726, 1.818728, 1.818729, 1.818729, 1.818729, 
    1.818729, 1.818728, 1.818729, 1.818729, 1.818729, 1.818731, 1.81873, 
    1.818731, 1.818731, 1.818721, 1.818721, 1.818721, 1.818722, 1.818721, 
    1.818723, 1.818723, 1.818725, 1.818725, 1.818726, 1.818725, 1.818725, 
    1.818726, 1.818725, 1.818727, 1.818726, 1.818729, 1.818727, 1.818729, 
    1.818729, 1.818729, 1.81873, 1.818731, 1.818732, 1.818732, 1.818733, 
    1.818722, 1.818723, 1.818723, 1.818723, 1.818724, 1.818725, 1.818727, 
    1.818726, 1.818727, 1.818727, 1.818726, 1.818727, 1.818723, 1.818724, 
    1.818723, 1.818722, 1.818726, 1.818724, 1.818728, 1.818727, 1.81873, 
    1.818728, 1.818731, 1.818733, 1.818734, 1.818735, 1.818723, 1.818723, 
    1.818723, 1.818725, 1.818725, 1.818727, 1.818727, 1.818727, 1.818728, 
    1.818728, 1.818727, 1.818728, 1.818724, 1.818726, 1.818722, 1.818724, 
    1.818724, 1.818724, 1.818726, 1.818726, 1.818728, 1.818727, 1.818732, 
    1.81873, 1.818737, 1.818735, 1.818722, 1.818723, 1.818725, 1.818724, 
    1.818727, 1.818727, 1.818728, 1.818729, 1.818729, 1.818729, 1.818729, 
    1.818729, 1.818727, 1.818728, 1.818725, 1.818726, 1.818725, 1.818725, 
    1.818726, 1.818727, 1.818727, 1.818728, 1.818729, 1.818727, 1.818733, 
    1.818729, 1.818724, 1.818725, 1.818725, 1.818725, 1.818727, 1.818726, 
    1.818729, 1.818728, 1.81873, 1.818729, 1.818729, 1.818728, 1.818728, 
    1.818726, 1.818725, 1.818725, 1.818725, 1.818726, 1.818727, 1.818729, 
    1.818729, 1.81873, 1.818727, 1.818728, 1.818727, 1.818729, 1.818726, 
    1.818728, 1.818725, 1.818726, 1.818726, 1.818728, 1.818728, 1.818729, 
    1.818728, 1.818727, 1.818727, 1.818726, 1.818726, 1.818725, 1.818725, 
    1.818725, 1.818726, 1.818727, 1.818729, 1.81873, 1.81873, 1.818732, 
    1.818731, 1.818733, 1.818731, 1.818734, 1.818728, 1.818731, 1.818726, 
    1.818727, 1.818728, 1.81873, 1.818729, 1.81873, 1.818727, 1.818726, 
    1.818725, 1.818725, 1.818725, 1.818725, 1.818726, 1.818726, 1.818727, 
    1.818727, 1.818729, 1.81873, 1.818733, 1.818734, 1.818736, 1.818736, 
    1.818737, 1.818737,
  1.818668, 1.818669, 1.818669, 1.818671, 1.81867, 1.818671, 1.818668, 
    1.81867, 1.818668, 1.818668, 1.818673, 1.818671, 1.818676, 1.818675, 
    1.818679, 1.818676, 1.81868, 1.818679, 1.818681, 1.818681, 1.818683, 
    1.818681, 1.818685, 1.818683, 1.818683, 1.818681, 1.818671, 1.818673, 
    1.818671, 1.818671, 1.818671, 1.81867, 1.818669, 1.818667, 1.818668, 
    1.818669, 1.818671, 1.818671, 1.818673, 1.818673, 1.818675, 1.818674, 
    1.818678, 1.818677, 1.818681, 1.81868, 1.818681, 1.81868, 1.818681, 
    1.818679, 1.81868, 1.818679, 1.818674, 1.818676, 1.818672, 1.81867, 
    1.818668, 1.818667, 1.818667, 1.818667, 1.818669, 1.81867, 1.818671, 
    1.818672, 1.818673, 1.818675, 1.818676, 1.818679, 1.818678, 1.818679, 
    1.81868, 1.818681, 1.818681, 1.818681, 1.818679, 1.81868, 1.818678, 
    1.818678, 1.818673, 1.818671, 1.81867, 1.818669, 1.818667, 1.818669, 
    1.818668, 1.818669, 1.81867, 1.81867, 1.818672, 1.818671, 1.818676, 
    1.818674, 1.81868, 1.818678, 1.81868, 1.818679, 1.81868, 1.818679, 
    1.818681, 1.818682, 1.818682, 1.818683, 1.818679, 1.818681, 1.81867, 
    1.81867, 1.81867, 1.818669, 1.818669, 1.818667, 1.818668, 1.818669, 
    1.81867, 1.818671, 1.818671, 1.818673, 1.818674, 1.818677, 1.818678, 
    1.818679, 1.818679, 1.818679, 1.818679, 1.818678, 1.818682, 1.81868, 
    1.818683, 1.818682, 1.818681, 1.818683, 1.81867, 1.818669, 1.818668, 
    1.818669, 1.818667, 1.818668, 1.818669, 1.818671, 1.818672, 1.818672, 
    1.818673, 1.818674, 1.818676, 1.818678, 1.81868, 1.81868, 1.81868, 
    1.81868, 1.818679, 1.81868, 1.81868, 1.81868, 1.818682, 1.818682, 
    1.818682, 1.818682, 1.81867, 1.81867, 1.81867, 1.818671, 1.81867, 
    1.818672, 1.818673, 1.818675, 1.818674, 1.818676, 1.818674, 1.818675, 
    1.818676, 1.818674, 1.818678, 1.818676, 1.81868, 1.818678, 1.81868, 
    1.81868, 1.81868, 1.818681, 1.818682, 1.818684, 1.818683, 1.818684, 
    1.818671, 1.818672, 1.818672, 1.818673, 1.818673, 1.818675, 1.818677, 
    1.818676, 1.818677, 1.818678, 1.818676, 1.818677, 1.818672, 1.818673, 
    1.818673, 1.818671, 1.818676, 1.818674, 1.818678, 1.818677, 1.818681, 
    1.818679, 1.818683, 1.818685, 1.818686, 1.818688, 1.818672, 1.818672, 
    1.818673, 1.818674, 1.818675, 1.818677, 1.818677, 1.818678, 1.818678, 
    1.818679, 1.818678, 1.818679, 1.818673, 1.818676, 1.818672, 1.818673, 
    1.818674, 1.818674, 1.818676, 1.818676, 1.818679, 1.818677, 1.818684, 
    1.818681, 1.818689, 1.818687, 1.818672, 1.818672, 1.818675, 1.818674, 
    1.818677, 1.818678, 1.818679, 1.81868, 1.81868, 1.81868, 1.818679, 
    1.81868, 1.818677, 1.818678, 1.818675, 1.818676, 1.818675, 1.818675, 
    1.818676, 1.818678, 1.818678, 1.818678, 1.81868, 1.818677, 1.818685, 
    1.81868, 1.818673, 1.818675, 1.818675, 1.818674, 1.818678, 1.818677, 
    1.81868, 1.818679, 1.818681, 1.81868, 1.81868, 1.818679, 1.818678, 
    1.818677, 1.818675, 1.818674, 1.818675, 1.818676, 1.818678, 1.81868, 
    1.818679, 1.818681, 1.818677, 1.818678, 1.818678, 1.818679, 1.818676, 
    1.818679, 1.818675, 1.818676, 1.818676, 1.818679, 1.818679, 1.81868, 
    1.818679, 1.818678, 1.818678, 1.818676, 1.818676, 1.818675, 1.818675, 
    1.818675, 1.818676, 1.818678, 1.818679, 1.818681, 1.818681, 1.818684, 
    1.818682, 1.818685, 1.818682, 1.818686, 1.818679, 1.818682, 1.818677, 
    1.818677, 1.818678, 1.818681, 1.818679, 1.818681, 1.818678, 1.818676, 
    1.818675, 1.818674, 1.818675, 1.818675, 1.818676, 1.818676, 1.818678, 
    1.818677, 1.81868, 1.818681, 1.818684, 1.818686, 1.818688, 1.818689, 
    1.818689, 1.81869,
  1.818639, 1.818641, 1.818641, 1.818642, 1.818642, 1.818643, 1.81864, 
    1.818641, 1.81864, 1.818639, 1.818646, 1.818642, 1.818649, 1.818647, 
    1.818652, 1.818648, 1.818653, 1.818652, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818656, 1.818656, 1.818654, 1.818643, 1.818645, 
    1.818643, 1.818643, 1.818643, 1.818642, 1.818641, 1.818639, 1.818639, 
    1.818641, 1.818643, 1.818642, 1.818645, 1.818645, 1.818648, 1.818646, 
    1.818651, 1.81865, 1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 
    1.818652, 1.818653, 1.818651, 1.818647, 1.818648, 1.818644, 1.818641, 
    1.81864, 1.818638, 1.818639, 1.818639, 1.818641, 1.818642, 1.818643, 
    1.818644, 1.818645, 1.818647, 1.818648, 1.818651, 1.818651, 1.818652, 
    1.818652, 1.818654, 1.818653, 1.818654, 1.818651, 1.818653, 1.81865, 
    1.818651, 1.818645, 1.818643, 1.818642, 1.818641, 1.818639, 1.81864, 
    1.81864, 1.818641, 1.818642, 1.818641, 1.818644, 1.818643, 1.818648, 
    1.818646, 1.818652, 1.818651, 1.818653, 1.818652, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818654, 1.818656, 1.818652, 1.818653, 1.818641, 
    1.818642, 1.818642, 1.81864, 1.81864, 1.818639, 1.81864, 1.818641, 
    1.818642, 1.818643, 1.818643, 1.818645, 1.818647, 1.818649, 1.818651, 
    1.818652, 1.818651, 1.818652, 1.818651, 1.818651, 1.818655, 1.818653, 
    1.818656, 1.818655, 1.818654, 1.818655, 1.818642, 1.818641, 1.81864, 
    1.818641, 1.818639, 1.81864, 1.818641, 1.818643, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818649, 1.818651, 1.818652, 1.818652, 1.818652, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 1.818655, 1.818655, 
    1.818655, 1.818655, 1.818641, 1.818642, 1.818642, 1.818642, 1.818642, 
    1.818644, 1.818645, 1.818648, 1.818646, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.818647, 1.81865, 1.818648, 1.818653, 1.81865, 1.818653, 
    1.818652, 1.818653, 1.818654, 1.818655, 1.818657, 1.818656, 1.818658, 
    1.818643, 1.818644, 1.818644, 1.818645, 1.818645, 1.818647, 1.818649, 
    1.818648, 1.81865, 1.81865, 1.818648, 1.818649, 1.818644, 1.818645, 
    1.818645, 1.818643, 1.818648, 1.818646, 1.818651, 1.818649, 1.818654, 
    1.818652, 1.818656, 1.818658, 1.81866, 1.818662, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818648, 1.818649, 1.81865, 1.81865, 1.818651, 
    1.818652, 1.81865, 1.818652, 1.818645, 1.818649, 1.818643, 1.818645, 
    1.818646, 1.818646, 1.818648, 1.818649, 1.818651, 1.81865, 1.818657, 
    1.818654, 1.818663, 1.818661, 1.818644, 1.818644, 1.818647, 1.818646, 
    1.81865, 1.81865, 1.818651, 1.818652, 1.818652, 1.818653, 1.818652, 
    1.818653, 1.818649, 1.818651, 1.818647, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.81865, 1.81865, 1.818651, 1.818652, 1.81865, 1.818658, 
    1.818653, 1.818645, 1.818647, 1.818647, 1.818646, 1.81865, 1.818649, 
    1.818653, 1.818652, 1.818654, 1.818653, 1.818653, 1.818651, 1.818651, 
    1.818649, 1.818648, 1.818646, 1.818647, 1.818648, 1.81865, 1.818652, 
    1.818652, 1.818653, 1.818649, 1.818651, 1.81865, 1.818652, 1.818648, 
    1.818652, 1.818648, 1.818648, 1.818649, 1.818651, 1.818652, 1.818652, 
    1.818652, 1.81865, 1.81865, 1.818649, 1.818649, 1.818648, 1.818647, 
    1.818648, 1.818648, 1.81865, 1.818652, 1.818654, 1.818654, 1.818657, 
    1.818655, 1.818658, 1.818655, 1.81866, 1.818652, 1.818655, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818652, 1.818654, 1.81865, 1.818648, 
    1.818648, 1.818647, 1.818648, 1.818647, 1.818648, 1.818648, 1.81865, 
    1.818649, 1.818653, 1.818654, 1.818657, 1.81866, 1.818662, 1.818663, 
    1.818663, 1.818663,
  1.818617, 1.818619, 1.818619, 1.818621, 1.81862, 1.818621, 1.818618, 
    1.818619, 1.818618, 1.818618, 1.818624, 1.818621, 1.818627, 1.818625, 
    1.81863, 1.818627, 1.818631, 1.81863, 1.818632, 1.818632, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818635, 1.818633, 1.818621, 1.818624, 
    1.818621, 1.818622, 1.818622, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818619, 1.818622, 1.818621, 1.818623, 1.818623, 1.818626, 1.818625, 
    1.818629, 1.818628, 1.818632, 1.818631, 1.818632, 1.818632, 1.818632, 
    1.81863, 1.818631, 1.81863, 1.818625, 1.818626, 1.818622, 1.81862, 
    1.818618, 1.818617, 1.818617, 1.818617, 1.818619, 1.81862, 1.818622, 
    1.818622, 1.818623, 1.818626, 1.818627, 1.81863, 1.818629, 1.81863, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.81863, 1.818632, 1.818629, 
    1.81863, 1.818623, 1.818621, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818618, 1.818619, 1.81862, 1.81862, 1.818622, 1.818621, 1.818627, 
    1.818624, 1.818631, 1.818629, 1.818631, 1.81863, 1.818632, 1.81863, 
    1.818633, 1.818633, 1.818633, 1.818634, 1.81863, 1.818632, 1.81862, 
    1.81862, 1.81862, 1.818619, 1.818619, 1.818617, 1.818618, 1.818619, 
    1.81862, 1.818621, 1.818622, 1.818623, 1.818625, 1.818628, 1.818629, 
    1.818631, 1.81863, 1.81863, 1.81863, 1.818629, 1.818633, 1.818631, 
    1.818634, 1.818634, 1.818633, 1.818634, 1.81862, 1.818619, 1.818618, 
    1.818619, 1.818617, 1.818618, 1.818619, 1.818621, 1.818622, 1.818622, 
    1.818623, 1.818625, 1.818627, 1.818629, 1.818631, 1.818631, 1.818631, 
    1.818631, 1.81863, 1.818631, 1.818632, 1.818631, 1.818634, 1.818633, 
    1.818634, 1.818633, 1.818619, 1.81862, 1.81862, 1.818621, 1.81862, 
    1.818622, 1.818623, 1.818626, 1.818625, 1.818627, 1.818625, 1.818625, 
    1.818627, 1.818625, 1.818629, 1.818626, 1.818631, 1.818629, 1.818631, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.818635, 1.818635, 1.818636, 
    1.818621, 1.818622, 1.818622, 1.818623, 1.818624, 1.818625, 1.818628, 
    1.818627, 1.818628, 1.818629, 1.818626, 1.818628, 1.818623, 1.818624, 
    1.818623, 1.818621, 1.818627, 1.818624, 1.818629, 1.818628, 1.818632, 
    1.81863, 1.818635, 1.818636, 1.818638, 1.81864, 1.818623, 1.818622, 
    1.818623, 1.818625, 1.818626, 1.818628, 1.818628, 1.818628, 1.818629, 
    1.81863, 1.818629, 1.81863, 1.818624, 1.818627, 1.818622, 1.818623, 
    1.818624, 1.818624, 1.818627, 1.818627, 1.81863, 1.818628, 1.818636, 
    1.818633, 1.818642, 1.818639, 1.818622, 1.818623, 1.818625, 1.818624, 
    1.818628, 1.818629, 1.81863, 1.818631, 1.818631, 1.818631, 1.81863, 
    1.818631, 1.818628, 1.81863, 1.818625, 1.818626, 1.818626, 1.818625, 
    1.818627, 1.818629, 1.818629, 1.818629, 1.818631, 1.818628, 1.818636, 
    1.818631, 1.818624, 1.818625, 1.818625, 1.818625, 1.818629, 1.818627, 
    1.818631, 1.81863, 1.818632, 1.818631, 1.818631, 1.81863, 1.818629, 
    1.818627, 1.818626, 1.818625, 1.818625, 1.818626, 1.818629, 1.818631, 
    1.81863, 1.818632, 1.818628, 1.81863, 1.818629, 1.818631, 1.818627, 
    1.81863, 1.818626, 1.818626, 1.818627, 1.81863, 1.81863, 1.818631, 
    1.81863, 1.818629, 1.818628, 1.818627, 1.818627, 1.818626, 1.818625, 
    1.818626, 1.818627, 1.818629, 1.81863, 1.818632, 1.818633, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818638, 1.81863, 1.818634, 1.818627, 
    1.818628, 1.818629, 1.818632, 1.818631, 1.818632, 1.818628, 1.818626, 
    1.818626, 1.818625, 1.818626, 1.818626, 1.818627, 1.818627, 1.818629, 
    1.818628, 1.818631, 1.818632, 1.818636, 1.818638, 1.818641, 1.818642, 
    1.818642, 1.818642,
  1.818569, 1.81857, 1.81857, 1.818572, 1.818571, 1.818572, 1.818569, 
    1.81857, 1.81857, 1.818569, 1.818574, 1.818572, 1.818577, 1.818576, 
    1.81858, 1.818577, 1.818581, 1.81858, 1.818582, 1.818581, 1.818584, 
    1.818582, 1.818585, 1.818583, 1.818584, 1.818582, 1.818572, 1.818574, 
    1.818572, 1.818572, 1.818572, 1.818571, 1.81857, 1.818568, 1.818569, 
    1.81857, 1.818572, 1.818572, 1.818574, 1.818574, 1.818576, 1.818575, 
    1.818579, 1.818578, 1.818581, 1.818581, 1.818581, 1.818581, 1.818581, 
    1.81858, 1.818581, 1.818579, 1.818575, 1.818576, 1.818573, 1.81857, 
    1.818569, 1.818568, 1.818568, 1.818568, 1.81857, 1.818571, 1.818572, 
    1.818573, 1.818574, 1.818576, 1.818577, 1.818579, 1.818579, 1.81858, 
    1.81858, 1.818582, 1.818581, 1.818582, 1.81858, 1.818581, 1.818579, 
    1.818579, 1.818574, 1.818572, 1.818571, 1.81857, 1.818568, 1.81857, 
    1.818569, 1.81857, 1.818571, 1.818571, 1.818573, 1.818572, 1.818577, 
    1.818575, 1.81858, 1.818579, 1.818581, 1.81858, 1.818581, 1.81858, 
    1.818582, 1.818583, 1.818582, 1.818583, 1.81858, 1.818581, 1.818571, 
    1.818571, 1.818571, 1.81857, 1.81857, 1.818568, 1.81857, 1.81857, 
    1.818571, 1.818572, 1.818572, 1.818574, 1.818575, 1.818578, 1.818579, 
    1.81858, 1.818579, 1.81858, 1.818579, 1.818579, 1.818582, 1.818581, 
    1.818583, 1.818583, 1.818582, 1.818583, 1.818571, 1.81857, 1.818569, 
    1.81857, 1.818568, 1.818569, 1.81857, 1.818572, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818577, 1.818579, 1.81858, 1.81858, 1.81858, 
    1.818581, 1.81858, 1.818581, 1.818581, 1.818581, 1.818583, 1.818582, 
    1.818583, 1.818583, 1.81857, 1.818571, 1.818571, 1.818571, 1.818571, 
    1.818573, 1.818573, 1.818576, 1.818575, 1.818577, 1.818575, 1.818576, 
    1.818577, 1.818575, 1.818579, 1.818576, 1.818581, 1.818578, 1.818581, 
    1.81858, 1.818581, 1.818582, 1.818583, 1.818584, 1.818584, 1.818585, 
    1.818572, 1.818573, 1.818573, 1.818574, 1.818574, 1.818576, 1.818578, 
    1.818577, 1.818578, 1.818579, 1.818576, 1.818578, 1.818573, 1.818574, 
    1.818574, 1.818572, 1.818577, 1.818574, 1.818579, 1.818578, 1.818582, 
    1.81858, 1.818584, 1.818585, 1.818587, 1.818589, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818576, 1.818578, 1.818578, 1.818578, 1.818579, 
    1.81858, 1.818578, 1.81858, 1.818574, 1.818577, 1.818573, 1.818574, 
    1.818575, 1.818574, 1.818577, 1.818577, 1.818579, 1.818578, 1.818585, 
    1.818582, 1.81859, 1.818588, 1.818573, 1.818573, 1.818576, 1.818575, 
    1.818578, 1.818579, 1.818579, 1.81858, 1.81858, 1.818581, 1.81858, 
    1.818581, 1.818578, 1.818579, 1.818576, 1.818576, 1.818576, 1.818576, 
    1.818577, 1.818578, 1.818578, 1.818579, 1.81858, 1.818578, 1.818585, 
    1.818581, 1.818574, 1.818575, 1.818576, 1.818575, 1.818579, 1.818577, 
    1.818581, 1.81858, 1.818582, 1.818581, 1.818581, 1.81858, 1.818579, 
    1.818577, 1.818576, 1.818575, 1.818575, 1.818576, 1.818578, 1.81858, 
    1.81858, 1.818581, 1.818578, 1.818579, 1.818579, 1.81858, 1.818577, 
    1.81858, 1.818576, 1.818576, 1.818577, 1.818579, 1.81858, 1.81858, 
    1.81858, 1.818579, 1.818578, 1.818577, 1.818577, 1.818576, 1.818576, 
    1.818576, 1.818577, 1.818579, 1.81858, 1.818582, 1.818582, 1.818584, 
    1.818583, 1.818585, 1.818583, 1.818587, 1.81858, 1.818583, 1.818577, 
    1.818578, 1.818579, 1.818582, 1.81858, 1.818582, 1.818578, 1.818577, 
    1.818576, 1.818575, 1.818576, 1.818576, 1.818577, 1.818577, 1.818579, 
    1.818578, 1.818581, 1.818582, 1.818585, 1.818587, 1.818589, 1.81859, 
    1.81859, 1.81859,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.293663e-09, 1.299371e-09, 1.298261e-09, 1.302865e-09, 1.300312e-09, 
    1.303326e-09, 1.29482e-09, 1.299597e-09, 1.296548e-09, 1.294177e-09, 
    1.3118e-09, 1.303071e-09, 1.32087e-09, 1.315302e-09, 1.329291e-09, 
    1.320004e-09, 1.331163e-09, 1.329023e-09, 1.335466e-09, 1.33362e-09, 
    1.341861e-09, 1.336318e-09, 1.346133e-09, 1.340537e-09, 1.341412e-09, 
    1.336135e-09, 1.304828e-09, 1.310714e-09, 1.304479e-09, 1.305318e-09, 
    1.304942e-09, 1.300364e-09, 1.298057e-09, 1.293227e-09, 1.294104e-09, 
    1.297652e-09, 1.305696e-09, 1.302965e-09, 1.309847e-09, 1.309692e-09, 
    1.317354e-09, 1.3139e-09, 1.326779e-09, 1.323118e-09, 1.333697e-09, 
    1.331037e-09, 1.333572e-09, 1.332803e-09, 1.333582e-09, 1.32968e-09, 
    1.331352e-09, 1.327919e-09, 1.314546e-09, 1.318476e-09, 1.306756e-09, 
    1.299709e-09, 1.29503e-09, 1.291709e-09, 1.292178e-09, 1.293073e-09, 
    1.297672e-09, 1.301997e-09, 1.305293e-09, 1.307497e-09, 1.30967e-09, 
    1.316245e-09, 1.319725e-09, 1.327519e-09, 1.326113e-09, 1.328495e-09, 
    1.330772e-09, 1.334594e-09, 1.333965e-09, 1.335649e-09, 1.328433e-09, 
    1.333228e-09, 1.325312e-09, 1.327477e-09, 1.310259e-09, 1.303702e-09, 
    1.300914e-09, 1.298475e-09, 1.292539e-09, 1.296638e-09, 1.295022e-09, 
    1.298866e-09, 1.301309e-09, 1.300101e-09, 1.307558e-09, 1.304659e-09, 
    1.319932e-09, 1.313353e-09, 1.330506e-09, 1.326401e-09, 1.33149e-09, 
    1.328894e-09, 1.333343e-09, 1.329339e-09, 1.336275e-09, 1.337786e-09, 
    1.336753e-09, 1.340719e-09, 1.329117e-09, 1.333572e-09, 1.300067e-09, 
    1.300264e-09, 1.301182e-09, 1.297147e-09, 1.2969e-09, 1.293203e-09, 
    1.296493e-09, 1.297894e-09, 1.301451e-09, 1.303555e-09, 1.305555e-09, 
    1.309952e-09, 1.314864e-09, 1.321733e-09, 1.326668e-09, 1.329976e-09, 
    1.327947e-09, 1.329738e-09, 1.327736e-09, 1.326798e-09, 1.33722e-09, 
    1.331367e-09, 1.340149e-09, 1.339663e-09, 1.335689e-09, 1.339717e-09, 
    1.300403e-09, 1.299269e-09, 1.295332e-09, 1.298413e-09, 1.2928e-09, 
    1.295942e-09, 1.297748e-09, 1.304719e-09, 1.306251e-09, 1.307671e-09, 
    1.310476e-09, 1.314076e-09, 1.320392e-09, 1.325887e-09, 1.330904e-09, 
    1.330537e-09, 1.330666e-09, 1.331787e-09, 1.329011e-09, 1.332243e-09, 
    1.332785e-09, 1.331367e-09, 1.339598e-09, 1.337246e-09, 1.339652e-09, 
    1.338121e-09, 1.299637e-09, 1.301545e-09, 1.300514e-09, 1.302453e-09, 
    1.301087e-09, 1.30716e-09, 1.308981e-09, 1.317502e-09, 1.314005e-09, 
    1.319571e-09, 1.314571e-09, 1.315457e-09, 1.319752e-09, 1.314841e-09, 
    1.325584e-09, 1.3183e-09, 1.33183e-09, 1.324556e-09, 1.332286e-09, 
    1.330883e-09, 1.333207e-09, 1.335288e-09, 1.337907e-09, 1.342739e-09, 
    1.34162e-09, 1.345661e-09, 1.30439e-09, 1.306864e-09, 1.306647e-09, 
    1.309236e-09, 1.311152e-09, 1.315304e-09, 1.321963e-09, 1.319459e-09, 
    1.324056e-09, 1.324979e-09, 1.317994e-09, 1.322283e-09, 1.308521e-09, 
    1.310744e-09, 1.30942e-09, 1.304585e-09, 1.320035e-09, 1.312106e-09, 
    1.326749e-09, 1.322453e-09, 1.334991e-09, 1.328755e-09, 1.341004e-09, 
    1.34624e-09, 1.351169e-09, 1.356928e-09, 1.308215e-09, 1.306534e-09, 
    1.309544e-09, 1.31371e-09, 1.317576e-09, 1.322715e-09, 1.323241e-09, 
    1.324204e-09, 1.326698e-09, 1.328795e-09, 1.324508e-09, 1.32932e-09, 
    1.311259e-09, 1.320724e-09, 1.305898e-09, 1.310362e-09, 1.313465e-09, 
    1.312104e-09, 1.319172e-09, 1.320839e-09, 1.327609e-09, 1.324109e-09, 
    1.344947e-09, 1.335728e-09, 1.361315e-09, 1.354163e-09, 1.305946e-09, 
    1.308209e-09, 1.316087e-09, 1.312339e-09, 1.323058e-09, 1.325697e-09, 
    1.327842e-09, 1.330584e-09, 1.33088e-09, 1.332505e-09, 1.329843e-09, 
    1.3324e-09, 1.322726e-09, 1.327049e-09, 1.315186e-09, 1.318073e-09, 
    1.316745e-09, 1.315288e-09, 1.319785e-09, 1.324575e-09, 1.324678e-09, 
    1.326214e-09, 1.330542e-09, 1.323102e-09, 1.346137e-09, 1.33191e-09, 
    1.310677e-09, 1.315037e-09, 1.31566e-09, 1.313971e-09, 1.325432e-09, 
    1.321279e-09, 1.332465e-09, 1.329442e-09, 1.334396e-09, 1.331934e-09, 
    1.331572e-09, 1.328411e-09, 1.326442e-09, 1.32147e-09, 1.317424e-09, 
    1.314216e-09, 1.314962e-09, 1.318486e-09, 1.324868e-09, 1.330907e-09, 
    1.329584e-09, 1.334019e-09, 1.322281e-09, 1.327203e-09, 1.3253e-09, 
    1.330261e-09, 1.319392e-09, 1.328647e-09, 1.317026e-09, 1.318045e-09, 
    1.321197e-09, 1.327536e-09, 1.32894e-09, 1.330437e-09, 1.329513e-09, 
    1.325031e-09, 1.324296e-09, 1.32112e-09, 1.320243e-09, 1.317824e-09, 
    1.31582e-09, 1.31765e-09, 1.319573e-09, 1.325033e-09, 1.329953e-09, 
    1.335318e-09, 1.336631e-09, 1.342899e-09, 1.337796e-09, 1.346216e-09, 
    1.339057e-09, 1.351451e-09, 1.329183e-09, 1.338847e-09, 1.32134e-09, 
    1.323226e-09, 1.326637e-09, 1.334461e-09, 1.330238e-09, 1.335178e-09, 
    1.324268e-09, 1.318607e-09, 1.317143e-09, 1.314411e-09, 1.317206e-09, 
    1.316978e-09, 1.319652e-09, 1.318793e-09, 1.325214e-09, 1.321765e-09, 
    1.331563e-09, 1.335139e-09, 1.345237e-09, 1.351429e-09, 1.357731e-09, 
    1.360514e-09, 1.361361e-09, 1.361715e-09 ;

 SOIL2_HR_S3 =
  9.240448e-11, 9.281221e-11, 9.273295e-11, 9.306182e-11, 9.287939e-11, 
    9.309473e-11, 9.248715e-11, 9.282839e-11, 9.261055e-11, 9.244119e-11, 
    9.370003e-11, 9.307649e-11, 9.434788e-11, 9.395015e-11, 9.494933e-11, 
    9.428597e-11, 9.50831e-11, 9.493022e-11, 9.539042e-11, 9.525858e-11, 
    9.584719e-11, 9.545127e-11, 9.615236e-11, 9.575266e-11, 9.581517e-11, 
    9.543821e-11, 9.320199e-11, 9.362239e-11, 9.317708e-11, 9.323702e-11, 
    9.321013e-11, 9.288315e-11, 9.271837e-11, 9.237333e-11, 9.243597e-11, 
    9.26894e-11, 9.326398e-11, 9.306895e-11, 9.356053e-11, 9.354943e-11, 
    9.409674e-11, 9.384996e-11, 9.476993e-11, 9.450845e-11, 9.526408e-11, 
    9.507404e-11, 9.525515e-11, 9.520024e-11, 9.525587e-11, 9.497715e-11, 
    9.509656e-11, 9.485132e-11, 9.389618e-11, 9.417687e-11, 9.333972e-11, 
    9.283638e-11, 9.250211e-11, 9.22649e-11, 9.229844e-11, 9.236236e-11, 
    9.269088e-11, 9.299979e-11, 9.32352e-11, 9.339267e-11, 9.354784e-11, 
    9.401747e-11, 9.42661e-11, 9.482279e-11, 9.472234e-11, 9.489252e-11, 
    9.505514e-11, 9.532813e-11, 9.52832e-11, 9.540347e-11, 9.488805e-11, 
    9.523059e-11, 9.466512e-11, 9.481978e-11, 9.358995e-11, 9.312157e-11, 
    9.292243e-11, 9.274818e-11, 9.232422e-11, 9.261699e-11, 9.250158e-11, 
    9.277618e-11, 9.295065e-11, 9.286436e-11, 9.339698e-11, 9.318991e-11, 
    9.428083e-11, 9.381092e-11, 9.503617e-11, 9.474296e-11, 9.510645e-11, 
    9.492097e-11, 9.523878e-11, 9.495275e-11, 9.544823e-11, 9.555613e-11, 
    9.548239e-11, 9.576563e-11, 9.49369e-11, 9.525514e-11, 9.286194e-11, 
    9.287602e-11, 9.294158e-11, 9.265335e-11, 9.263572e-11, 9.237161e-11, 
    9.260662e-11, 9.27067e-11, 9.296078e-11, 9.311105e-11, 9.325392e-11, 
    9.356804e-11, 9.391886e-11, 9.440947e-11, 9.476197e-11, 9.499826e-11, 
    9.485337e-11, 9.498129e-11, 9.483829e-11, 9.477127e-11, 9.551569e-11, 
    9.509768e-11, 9.572489e-11, 9.569019e-11, 9.540633e-11, 9.56941e-11, 
    9.28859e-11, 9.280491e-11, 9.252371e-11, 9.274378e-11, 9.234285e-11, 
    9.256725e-11, 9.269629e-11, 9.319422e-11, 9.330364e-11, 9.340508e-11, 
    9.360545e-11, 9.386259e-11, 9.43137e-11, 9.470624e-11, 9.50646e-11, 
    9.503834e-11, 9.504759e-11, 9.512763e-11, 9.492934e-11, 9.516019e-11, 
    9.519893e-11, 9.509763e-11, 9.568554e-11, 9.551758e-11, 9.568945e-11, 
    9.558009e-11, 9.283124e-11, 9.296752e-11, 9.289387e-11, 9.303235e-11, 
    9.293479e-11, 9.336858e-11, 9.349865e-11, 9.410731e-11, 9.385753e-11, 
    9.425508e-11, 9.389792e-11, 9.39612e-11, 9.426802e-11, 9.391722e-11, 
    9.468458e-11, 9.41643e-11, 9.513074e-11, 9.461114e-11, 9.516331e-11, 
    9.506305e-11, 9.522905e-11, 9.537773e-11, 9.556478e-11, 9.590991e-11, 
    9.583e-11, 9.611864e-11, 9.317069e-11, 9.334745e-11, 9.33319e-11, 
    9.351689e-11, 9.36537e-11, 9.395026e-11, 9.44259e-11, 9.424705e-11, 
    9.457542e-11, 9.464134e-11, 9.414246e-11, 9.444875e-11, 9.346576e-11, 
    9.362455e-11, 9.353001e-11, 9.318463e-11, 9.428824e-11, 9.372184e-11, 
    9.476779e-11, 9.446093e-11, 9.535653e-11, 9.491111e-11, 9.5786e-11, 
    9.616e-11, 9.651208e-11, 9.692346e-11, 9.344393e-11, 9.332382e-11, 
    9.353889e-11, 9.383644e-11, 9.411256e-11, 9.447964e-11, 9.451721e-11, 
    9.458598e-11, 9.476412e-11, 9.49139e-11, 9.460771e-11, 9.495145e-11, 
    9.366136e-11, 9.433741e-11, 9.327841e-11, 9.359726e-11, 9.38189e-11, 
    9.372169e-11, 9.422661e-11, 9.434561e-11, 9.482921e-11, 9.457922e-11, 
    9.606768e-11, 9.540911e-11, 9.723675e-11, 9.672596e-11, 9.328185e-11, 
    9.344352e-11, 9.400618e-11, 9.373847e-11, 9.450415e-11, 9.469264e-11, 
    9.484587e-11, 9.504172e-11, 9.506288e-11, 9.517893e-11, 9.498876e-11, 
    9.517143e-11, 9.448042e-11, 9.478921e-11, 9.394189e-11, 9.414811e-11, 
    9.405324e-11, 9.394917e-11, 9.427036e-11, 9.461253e-11, 9.461985e-11, 
    9.472957e-11, 9.503872e-11, 9.450726e-11, 9.615264e-11, 9.513643e-11, 
    9.361981e-11, 9.39312e-11, 9.39757e-11, 9.385508e-11, 9.467373e-11, 
    9.43771e-11, 9.517611e-11, 9.496016e-11, 9.531399e-11, 9.513817e-11, 
    9.511229e-11, 9.488647e-11, 9.474588e-11, 9.439069e-11, 9.410171e-11, 
    9.387257e-11, 9.392585e-11, 9.417755e-11, 9.463346e-11, 9.506479e-11, 
    9.49703e-11, 9.52871e-11, 9.444864e-11, 9.48002e-11, 9.466431e-11, 
    9.501865e-11, 9.424229e-11, 9.490333e-11, 9.407332e-11, 9.414609e-11, 
    9.437121e-11, 9.482403e-11, 9.492425e-11, 9.503122e-11, 9.496522e-11, 
    9.464504e-11, 9.459259e-11, 9.436574e-11, 9.430309e-11, 9.413025e-11, 
    9.398714e-11, 9.411789e-11, 9.425519e-11, 9.464518e-11, 9.499664e-11, 
    9.537984e-11, 9.547363e-11, 9.592133e-11, 9.555685e-11, 9.61583e-11, 
    9.564691e-11, 9.65322e-11, 9.494167e-11, 9.563191e-11, 9.438145e-11, 
    9.451617e-11, 9.47598e-11, 9.531868e-11, 9.501698e-11, 9.536982e-11, 
    9.459054e-11, 9.418624e-11, 9.408165e-11, 9.38865e-11, 9.408611e-11, 
    9.406988e-11, 9.42609e-11, 9.419951e-11, 9.465813e-11, 9.441178e-11, 
    9.511164e-11, 9.536704e-11, 9.608839e-11, 9.65306e-11, 9.698082e-11, 
    9.717958e-11, 9.724007e-11, 9.726536e-11 ;

 SOIL3C =
  5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611 ;

 SOIL3C_TO_SOIL1C =
  2.55107e-11, 2.562324e-11, 2.560136e-11, 2.569213e-11, 2.564178e-11, 
    2.570122e-11, 2.553352e-11, 2.56277e-11, 2.556758e-11, 2.552083e-11, 
    2.586829e-11, 2.569618e-11, 2.604711e-11, 2.593733e-11, 2.621312e-11, 
    2.603002e-11, 2.625004e-11, 2.620784e-11, 2.633486e-11, 2.629848e-11, 
    2.646094e-11, 2.635166e-11, 2.654517e-11, 2.643485e-11, 2.64521e-11, 
    2.634806e-11, 2.573082e-11, 2.584686e-11, 2.572395e-11, 2.574049e-11, 
    2.573307e-11, 2.564282e-11, 2.559734e-11, 2.55021e-11, 2.551939e-11, 
    2.558934e-11, 2.574794e-11, 2.56941e-11, 2.582979e-11, 2.582672e-11, 
    2.597779e-11, 2.590968e-11, 2.61636e-11, 2.609143e-11, 2.629999e-11, 
    2.624754e-11, 2.629753e-11, 2.628237e-11, 2.629773e-11, 2.62208e-11, 
    2.625376e-11, 2.618607e-11, 2.592243e-11, 2.599991e-11, 2.576884e-11, 
    2.562991e-11, 2.553764e-11, 2.547217e-11, 2.548143e-11, 2.549907e-11, 
    2.558975e-11, 2.567501e-11, 2.573999e-11, 2.578346e-11, 2.582628e-11, 
    2.595591e-11, 2.602454e-11, 2.617819e-11, 2.615047e-11, 2.619744e-11, 
    2.624232e-11, 2.631767e-11, 2.630527e-11, 2.633847e-11, 2.61962e-11, 
    2.629075e-11, 2.613467e-11, 2.617736e-11, 2.583791e-11, 2.570863e-11, 
    2.565366e-11, 2.560557e-11, 2.548855e-11, 2.556936e-11, 2.55375e-11, 
    2.561329e-11, 2.566145e-11, 2.563763e-11, 2.578465e-11, 2.572749e-11, 
    2.60286e-11, 2.58989e-11, 2.623709e-11, 2.615616e-11, 2.625648e-11, 
    2.620529e-11, 2.629301e-11, 2.621406e-11, 2.635082e-11, 2.63806e-11, 
    2.636025e-11, 2.643843e-11, 2.620969e-11, 2.629753e-11, 2.563697e-11, 
    2.564085e-11, 2.565895e-11, 2.557939e-11, 2.557453e-11, 2.550163e-11, 
    2.556649e-11, 2.559412e-11, 2.566425e-11, 2.570572e-11, 2.574516e-11, 
    2.583186e-11, 2.592869e-11, 2.606411e-11, 2.61614e-11, 2.622662e-11, 
    2.618663e-11, 2.622194e-11, 2.618247e-11, 2.616397e-11, 2.636944e-11, 
    2.625406e-11, 2.642719e-11, 2.641761e-11, 2.633926e-11, 2.641868e-11, 
    2.564358e-11, 2.562122e-11, 2.554361e-11, 2.560435e-11, 2.549369e-11, 
    2.555563e-11, 2.559124e-11, 2.572868e-11, 2.575888e-11, 2.578688e-11, 
    2.584219e-11, 2.591316e-11, 2.603768e-11, 2.614602e-11, 2.624493e-11, 
    2.623769e-11, 2.624024e-11, 2.626233e-11, 2.62076e-11, 2.627132e-11, 
    2.628201e-11, 2.625405e-11, 2.641632e-11, 2.636996e-11, 2.64174e-11, 
    2.638722e-11, 2.562849e-11, 2.566611e-11, 2.564578e-11, 2.5684e-11, 
    2.565707e-11, 2.577681e-11, 2.581271e-11, 2.598071e-11, 2.591176e-11, 
    2.602149e-11, 2.592291e-11, 2.594038e-11, 2.602507e-11, 2.592824e-11, 
    2.614004e-11, 2.599644e-11, 2.626319e-11, 2.611977e-11, 2.627218e-11, 
    2.624451e-11, 2.629033e-11, 2.633136e-11, 2.638299e-11, 2.647825e-11, 
    2.645619e-11, 2.653587e-11, 2.572218e-11, 2.577097e-11, 2.576668e-11, 
    2.581774e-11, 2.585551e-11, 2.593736e-11, 2.606865e-11, 2.601928e-11, 
    2.610991e-11, 2.612811e-11, 2.599041e-11, 2.607495e-11, 2.580363e-11, 
    2.584746e-11, 2.582136e-11, 2.572603e-11, 2.603065e-11, 2.587431e-11, 
    2.616301e-11, 2.607831e-11, 2.632551e-11, 2.620257e-11, 2.644405e-11, 
    2.654728e-11, 2.664446e-11, 2.6758e-11, 2.57976e-11, 2.576445e-11, 
    2.582382e-11, 2.590594e-11, 2.598216e-11, 2.608348e-11, 2.609385e-11, 
    2.611283e-11, 2.6162e-11, 2.620334e-11, 2.611883e-11, 2.62137e-11, 
    2.585762e-11, 2.604422e-11, 2.575192e-11, 2.583993e-11, 2.59011e-11, 
    2.587427e-11, 2.601364e-11, 2.604648e-11, 2.617996e-11, 2.611096e-11, 
    2.65218e-11, 2.634002e-11, 2.684448e-11, 2.670349e-11, 2.575287e-11, 
    2.579749e-11, 2.59528e-11, 2.58789e-11, 2.609024e-11, 2.614227e-11, 
    2.618456e-11, 2.623862e-11, 2.624446e-11, 2.627649e-11, 2.6224e-11, 
    2.627442e-11, 2.608369e-11, 2.616892e-11, 2.593505e-11, 2.599197e-11, 
    2.596578e-11, 2.593706e-11, 2.602571e-11, 2.612015e-11, 2.612218e-11, 
    2.615246e-11, 2.623779e-11, 2.60911e-11, 2.654525e-11, 2.626476e-11, 
    2.584615e-11, 2.59321e-11, 2.594438e-11, 2.591109e-11, 2.613705e-11, 
    2.605517e-11, 2.627571e-11, 2.621611e-11, 2.631377e-11, 2.626524e-11, 
    2.62581e-11, 2.619577e-11, 2.615696e-11, 2.605893e-11, 2.597916e-11, 
    2.591592e-11, 2.593062e-11, 2.60001e-11, 2.612593e-11, 2.624499e-11, 
    2.621891e-11, 2.630635e-11, 2.607492e-11, 2.617196e-11, 2.613445e-11, 
    2.623225e-11, 2.601796e-11, 2.620042e-11, 2.597133e-11, 2.599141e-11, 
    2.605355e-11, 2.617853e-11, 2.62062e-11, 2.623572e-11, 2.62175e-11, 
    2.612913e-11, 2.611465e-11, 2.605204e-11, 2.603475e-11, 2.598704e-11, 
    2.594754e-11, 2.598363e-11, 2.602153e-11, 2.612917e-11, 2.622618e-11, 
    2.633194e-11, 2.635783e-11, 2.648141e-11, 2.63808e-11, 2.654681e-11, 
    2.640566e-11, 2.665001e-11, 2.6211e-11, 2.640152e-11, 2.605638e-11, 
    2.609356e-11, 2.616081e-11, 2.631506e-11, 2.623179e-11, 2.632918e-11, 
    2.611409e-11, 2.600249e-11, 2.597363e-11, 2.591976e-11, 2.597486e-11, 
    2.597038e-11, 2.60231e-11, 2.600616e-11, 2.613274e-11, 2.606475e-11, 
    2.625792e-11, 2.632841e-11, 2.652751e-11, 2.664957e-11, 2.677383e-11, 
    2.68287e-11, 2.684539e-11, 2.685237e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  -2.569961e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 0, 
    2.569961e-21, 2.055969e-20, 3.009266e-36, -1.28498e-20, -2.569961e-21, 
    -1.28498e-20, -1.28498e-20, 1.541976e-20, 1.541976e-20, -7.709882e-21, 
    -2.569961e-20, 7.709882e-21, 2.569961e-21, 2.569961e-21, -1.28498e-20, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 1.28498e-20, 0, 2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 1.28498e-20, -7.709882e-21, -1.027984e-20, 
    -7.709882e-21, -1.027984e-20, 7.709882e-21, -7.709882e-21, -1.541976e-20, 
    -1.027984e-20, 2.569961e-21, -1.541976e-20, -7.709882e-21, 1.027984e-20, 
    1.003089e-36, 1.003089e-36, -5.139921e-21, -1.027984e-20, 1.28498e-20, 
    -1.798972e-20, 1.28498e-20, -7.709882e-21, -5.139921e-21, 1.003089e-36, 
    -1.003089e-36, -2.569961e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 1.003089e-36, 1.798972e-20, -1.541976e-20, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -1.798972e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, -1.541976e-20, -2.569961e-21, 
    -1.541976e-20, 7.709882e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    1.027984e-20, 2.569961e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, -1.28498e-20, 7.709882e-21, 1.28498e-20, -1.027984e-20, 
    7.709882e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, -7.709882e-21, 
    -2.569961e-21, 0, -7.709882e-21, 5.139921e-21, 0, 7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 1.003089e-36, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, 2.312965e-20, -7.709882e-21, -1.003089e-36, 
    -1.027984e-20, -2.055969e-20, 7.709882e-21, -1.28498e-20, -1.798972e-20, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, 0, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -1.541976e-20, -2.569961e-21, 
    1.003089e-36, -1.541976e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -1.541976e-20, -2.569961e-21, 7.709882e-21, -2.569961e-21, -1.003089e-36, 
    1.28498e-20, 5.139921e-21, 1.541976e-20, 1.003089e-36, 5.139921e-21, 
    -2.055969e-20, 1.28498e-20, 5.139921e-21, -5.139921e-21, 2.055969e-20, 
    2.569961e-21, -2.055969e-20, 7.709882e-21, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, 2.569961e-21, -1.027984e-20, 2.569961e-21, -1.003089e-36, 
    -1.027984e-20, -1.541976e-20, 1.003089e-36, 0, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -1.541976e-20, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, -1.28498e-20, 1.798972e-20, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -1.28498e-20, 1.28498e-20, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    1.541976e-20, -2.569961e-21, 2.569961e-21, 0, -1.541976e-20, 
    2.055969e-20, 2.312965e-20, 1.541976e-20, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, 0, 5.139921e-21, -1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, -2.312965e-20, 2.569961e-21, 2.569961e-21, 
    1.798972e-20, 7.709882e-21, -5.139921e-21, -1.28498e-20, -1.28498e-20, 0, 
    -1.027984e-20, 7.709882e-21, 2.055969e-20, 2.312965e-20, -7.709882e-21, 
    -1.798972e-20, 1.541976e-20, 2.569961e-21, -7.709882e-21, 1.28498e-20, 
    -2.569961e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.541976e-20, -1.28498e-20, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, 1.027984e-20, 7.709882e-21, 
    -1.798972e-20, 1.003089e-36, -5.139921e-21, -2.569961e-21, 0, 
    2.055969e-20, 7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 1.541976e-20, -3.083953e-20, -2.569961e-21, 1.541976e-20, 
    -7.709882e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, 7.709882e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, 
    1.541976e-20, 7.709882e-21, -7.709882e-21, 5.139921e-21, 2.312965e-20, 
    -1.798972e-20, -2.055969e-20, -2.569961e-21, 7.709882e-21, -2.312965e-20, 
    -1.798972e-20, -7.709882e-21, -7.709882e-21, 0, 5.139921e-21, 
    -1.541976e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 1.28498e-20, 1.28498e-20, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, 1.003089e-36, 7.709882e-21, 1.027984e-20, -1.003089e-36, 
    -1.798972e-20, 0, -2.569961e-21, -5.139921e-21, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, -1.798972e-20, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, 1.027984e-20, -7.709882e-21, 
    -1.003089e-36, -1.027984e-20, -5.139921e-21, 1.003089e-36, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -1.798972e-20, 1.541976e-20, 2.569961e-21, 
    -1.003089e-36,
  0, -2.569961e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, 0, 2.569961e-21, -5.139921e-21, 0, 2.569961e-21, 
    -2.569961e-21, 0, 1.027984e-20, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 0, -7.709882e-21, -2.569961e-21, 0, -1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, 0, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.798972e-20, 2.055969e-20, 0, 
    -5.139921e-21, -7.709882e-21, 0, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 7.709882e-21, -2.569961e-21, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, -1.027984e-20, 0, 2.569961e-21, -2.569961e-21, 
    -1.541976e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 0, 5.139921e-21, 0, 1.28498e-20, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    0, -7.709882e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, -1.027984e-20, 2.569961e-21, -1.798972e-20, 0, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    0, 1.027984e-20, 5.139921e-21, -7.709882e-21, 5.139921e-21, 7.709882e-21, 
    -1.003089e-36, 7.709882e-21, -1.541976e-20, -1.798972e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, 7.709882e-21, 0, 
    1.027984e-20, 5.139921e-21, -7.709882e-21, 5.139921e-21, -7.709882e-21, 
    0, -5.139921e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 
    1.28498e-20, -5.139921e-21, 1.28498e-20, -2.569961e-21, 2.569961e-21, 
    1.003089e-36, -7.709882e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, 1.28498e-20, 1.027984e-20, -1.003089e-36, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 1.28498e-20, -7.709882e-21, -5.139921e-21, 
    0, -1.541976e-20, 1.541976e-20, -7.709882e-21, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -1.003089e-36, 0, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 0, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, 1.003089e-36, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    1.28498e-20, 7.709882e-21, 1.027984e-20, -7.709882e-21, 0, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, -5.139921e-21, -1.28498e-20, 
    0, 5.139921e-21, -1.541976e-20, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, -1.541976e-20, -2.569961e-21, -1.28498e-20, 1.798972e-20, 
    5.139921e-21, -1.541976e-20, -7.709882e-21, 1.798972e-20, -1.28498e-20, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 0, 
    -2.569961e-21, 1.027984e-20, 1.541976e-20, -1.027984e-20, -5.139921e-21, 
    -1.28498e-20, -1.027984e-20, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -1.003089e-36, -2.569961e-21, 1.003089e-36, 
    1.798972e-20, 5.139921e-21, -5.139921e-21, 0, 0, -5.139921e-21, 
    7.709882e-21, 1.027984e-20, 2.569961e-21, 0, -2.569961e-21, 1.28498e-20, 
    7.709882e-21, -5.139921e-21, 1.28498e-20, 1.541976e-20, 2.569961e-21, 
    1.027984e-20, -7.709882e-21, 2.569961e-21, 0, 0, 0, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 0, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, 0, -5.139921e-21, 1.28498e-20, 2.569961e-21, 
    5.139921e-21, -2.055969e-20, 7.709882e-21, -1.798972e-20, 0, 
    -1.541976e-20, 0, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -1.003089e-36, 1.027984e-20, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, 0, 0, 7.709882e-21, 
    -1.28498e-20, 0, 2.569961e-21, 0, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 0, -7.709882e-21, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, -7.709882e-21, -1.003089e-36, -2.569961e-21, 
    -1.28498e-20, 7.709882e-21, -5.139921e-21, 1.28498e-20, -7.709882e-21, 0, 
    -1.003089e-36, 0, 0, -5.139921e-21, 5.139921e-21, -2.569961e-21,
  1.541976e-20, 2.569961e-21, 5.139921e-21, 0, 0, 1.28498e-20, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, -1.027984e-20, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, -1.003089e-36, 0, 
    -1.027984e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -1.798972e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 2.826957e-20, -1.541976e-20, -1.798972e-20, 1.003089e-36, 
    0, 1.28498e-20, 2.569961e-21, 5.139921e-21, 0, -2.312965e-20, 
    7.709882e-21, -2.569961e-21, 1.003089e-36, 1.027984e-20, 2.569961e-21, 
    1.027984e-20, 1.027984e-20, 7.709882e-21, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 0, 2.569961e-21, 7.709882e-21, 
    -1.027984e-20, -1.027984e-20, 0, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -1.28498e-20, -1.28498e-20, -1.027984e-20, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, 7.709882e-21, -1.027984e-20, 1.28498e-20, -1.798972e-20, 
    1.027984e-20, -1.027984e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -5.139921e-21, 0, 1.003089e-36, 
    -2.569961e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -1.541976e-20, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 0, 
    1.541976e-20, 1.541976e-20, -7.709882e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-20, 1.027984e-20, -1.003089e-36, -2.569961e-21, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -1.541976e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    0, 0, 1.28498e-20, 0, -1.541976e-20, -7.709882e-21, 5.139921e-21, 
    -1.003089e-36, 7.709882e-21, -2.569961e-21, 1.027984e-20, 0, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -1.28498e-20, -5.139921e-21, 0, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 2.312965e-20, -1.541976e-20, -2.569961e-21, 
    -5.139921e-21, -1.798972e-20, 1.28498e-20, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, 
    2.569961e-21, 1.027984e-20, 0, 7.709882e-21, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, -1.28498e-20, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, 1.027984e-20, 0, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, 0, -7.709882e-21, 
    -1.027984e-20, 1.027984e-20, -1.027984e-20, -2.569961e-21, 0, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.28498e-20, 1.541976e-20, 0, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    -1.541976e-20, -7.709882e-21, -7.709882e-21, -1.003089e-36, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, 2.055969e-20, 1.003089e-36, 1.541976e-20, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -2.312965e-20, 1.027984e-20, 0, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 0, -1.003089e-36, -5.139921e-21, 7.709882e-21, 
    1.003089e-36, 7.709882e-21, -1.027984e-20, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    0, -2.569961e-21, -1.003089e-36, -7.709882e-21, 5.139921e-21, 0, 
    1.541976e-20, -7.709882e-21, -1.798972e-20, 0, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, 7.709882e-21, -1.541976e-20, 
    -1.027984e-20, -5.139921e-21, -2.569961e-21, 0, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, 0, 5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, 0, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, 1.003089e-36, 5.139921e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, -2.055969e-20, 5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -7.709882e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, 0, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, -2.569961e-21, -1.798972e-20, -5.139921e-21, 
    1.003089e-36, 0, -1.027984e-20, -1.027984e-20, -7.709882e-21, 
    1.027984e-20, 0, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 0, -2.569961e-21, 5.139921e-21, 0, 
    -5.139921e-21, -1.003089e-36, 5.139921e-21,
  0, 1.28498e-20, 2.569961e-21, -5.139921e-21, 1.027984e-20, 0, 2.569961e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 1.28498e-20, 
    -1.027984e-20, 7.709882e-21, 0, 1.28498e-20, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.003089e-36, 1.541976e-20, 7.709882e-21, 1.003089e-36, 
    7.709882e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    -1.28498e-20, -1.003089e-36, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, -2.055969e-20, 
    -1.003089e-36, -1.027984e-20, 1.28498e-20, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, -1.798972e-20, 0, -1.027984e-20, 
    -1.003089e-36, -5.139921e-21, 1.798972e-20, -1.541976e-20, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, 7.709882e-21, -1.003089e-36, -1.28498e-20, 
    -1.027984e-20, 1.541976e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    1.798972e-20, -5.139921e-21, 1.28498e-20, 0, 1.541976e-20, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 2.569961e-20, 
    1.027984e-20, 1.027984e-20, -2.569961e-21, 2.569961e-21, 0, 1.027984e-20, 
    1.798972e-20, 2.569961e-21, -1.027984e-20, -1.003089e-36, 5.139921e-21, 
    -1.027984e-20, -1.003089e-36, 1.541976e-20, -1.027984e-20, 1.28498e-20, 
    -7.709882e-21, -1.28498e-20, 1.027984e-20, 2.569961e-21, -1.541976e-20, 
    1.28498e-20, 7.709882e-21, 5.139921e-21, -1.003089e-36, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, -1.003089e-36, 
    0, 2.569961e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.798972e-20, -2.569961e-21, 7.709882e-21, -2.055969e-20, -7.709882e-21, 
    -1.541976e-20, 1.003089e-36, -1.798972e-20, 0, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, 1.003089e-36, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    0, -5.139921e-21, 5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 
    1.28498e-20, 7.709882e-21, 2.312965e-20, 1.003089e-36, 5.139921e-21, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -2.055969e-20, 1.28498e-20, 1.003089e-36, 1.28498e-20, 
    2.569961e-21, -1.003089e-36, -1.027984e-20, -2.569961e-21, -2.312965e-20, 
    1.003089e-36, -5.139921e-21, 7.709882e-21, 1.28498e-20, -1.798972e-20, 
    -1.28498e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -2.826957e-20, -7.709882e-21, -5.139921e-21, 0, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 1.28498e-20, -1.541976e-20, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, -1.003089e-36, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    1.003089e-36, -2.569961e-21, 1.027984e-20, 1.003089e-36, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.798972e-20, 1.003089e-36, -1.28498e-20, 5.139921e-21, 
    2.569961e-21, 1.541976e-20, 1.003089e-36, -1.027984e-20, 1.28498e-20, 
    7.709882e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, 1.027984e-20, 
    -2.569961e-20, -2.569961e-21, 1.28498e-20, 5.139921e-21, -1.798972e-20, 
    -1.28498e-20, 5.139921e-21, 5.139921e-21, 2.569961e-21, -1.798972e-20, 
    1.798972e-20, 2.569961e-21, 1.003089e-36, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 7.709882e-21, 1.28498e-20, -7.709882e-21, 7.709882e-21, 
    1.027984e-20, -5.139921e-21, -7.709882e-21, -1.798972e-20, 2.569961e-21, 
    -1.798972e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    1.798972e-20, -2.569961e-21, 1.541976e-20, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 1.28498e-20, 5.139921e-21, 1.027984e-20, -1.541976e-20, 
    1.28498e-20, 5.139921e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, 1.003089e-36, 0, -7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 5.139921e-21, -1.027984e-20, 1.28498e-20, 
    1.027984e-20, -2.569961e-21, -1.798972e-20, 1.28498e-20, 1.003089e-36, 
    -7.709882e-21, -5.139921e-21, -1.027984e-20, 1.798972e-20, -2.569961e-21, 
    1.28498e-20, -1.027984e-20, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    -1.28498e-20, -5.139921e-21, 5.139921e-21, 1.28498e-20, -5.139921e-21, 
    1.28498e-20, 5.139921e-21, 0, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21,
  7.709882e-21, 7.709882e-21, 1.003089e-36, 1.28498e-20, -5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -1.798972e-20, -1.541976e-20, 
    -1.027984e-20, -1.798972e-20, 7.709882e-21, 1.798972e-20, 2.055969e-20, 
    1.28498e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, -1.798972e-20, 
    -1.027984e-20, 0, 0, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, -1.003089e-36, 2.569961e-21, 1.28498e-20, 1.003089e-36, 
    5.139921e-21, -1.541976e-20, -2.569961e-21, 1.027984e-20, 1.541976e-20, 
    5.139921e-21, 1.541976e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, -1.798972e-20, 5.139921e-21, -1.28498e-20, 
    -5.139921e-21, -1.027984e-20, 1.541976e-20, -1.027984e-20, 2.569961e-21, 
    -1.28498e-20, 7.709882e-21, 7.709882e-21, -2.569961e-21, -1.003089e-36, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, -1.541976e-20, 2.569961e-21, 
    -2.569961e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 1.28498e-20, 1.003089e-36, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, -1.003089e-36, -7.709882e-21, 0, 
    -1.003089e-36, 7.709882e-21, -1.28498e-20, -1.541976e-20, 1.003089e-36, 
    -5.139921e-21, -5.139921e-21, -5.015443e-37, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, -2.826957e-20, 0, -2.569961e-20, 1.027984e-20, 
    2.569961e-21, -1.28498e-20, 5.139921e-21, 7.709882e-21, -1.28498e-20, 
    2.569961e-21, 2.312965e-20, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 0, 1.28498e-20, 5.139921e-21, 
    -2.569961e-21, -1.798972e-20, -1.003089e-36, 0, -1.541976e-20, 
    -1.798972e-20, 1.003089e-36, 1.28498e-20, -1.798972e-20, -1.027984e-20, 
    -7.709882e-21, 1.541976e-20, 1.003089e-36, 5.139921e-21, 2.569961e-21, 
    -2.569961e-20, -1.003089e-36, 7.709882e-21, -7.709882e-21, 0, 
    5.139921e-21, -7.709882e-21, 1.28498e-20, 2.569961e-21, 1.541976e-20, 
    2.569961e-21, 2.569961e-21, 2.569961e-20, 2.569961e-21, 1.541976e-20, 
    1.541976e-20, -1.541976e-20, -1.541976e-20, -2.312965e-20, 2.569961e-21, 
    -2.569961e-20, 1.798972e-20, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 2.312965e-20, 5.139921e-21, -1.28498e-20, 5.139921e-21, 
    7.709882e-21, -1.027984e-20, 1.027984e-20, 7.709882e-21, 2.569961e-21, 
    1.798972e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 1.28498e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, -1.28498e-20, 
    1.798972e-20, -7.709882e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 1.28498e-20, 1.28498e-20, 7.709882e-21, 2.569961e-21, 
    1.541976e-20, 1.027984e-20, 1.003089e-36, -7.709882e-21, 1.027984e-20, 
    7.709882e-21, 1.28498e-20, -1.28498e-20, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 1.798972e-20, -1.003089e-36, -2.569961e-21, 1.28498e-20, 
    -1.027984e-20, 1.28498e-20, -1.003089e-36, -5.139921e-21, -2.055969e-20, 
    -1.027984e-20, 7.709882e-21, -1.003089e-36, 7.709882e-21, 7.709882e-21, 
    1.027984e-20, 2.569961e-21, 0, -1.28498e-20, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 1.541976e-20, -2.569961e-21, 2.055969e-20, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, -1.003089e-36, 7.709882e-21, 
    1.541976e-20, -1.541976e-20, 2.569961e-21, 1.027984e-20, -1.027984e-20, 
    -3.340949e-20, -1.003089e-36, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    1.28498e-20, 5.139921e-21, 1.003089e-36, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 1.28498e-20, -1.28498e-20, 2.569961e-21, 2.055969e-20, 
    -2.569961e-21, 1.798972e-20, 1.003089e-36, -7.709882e-21, 1.027984e-20, 
    -1.28498e-20, 2.569961e-21, -1.541976e-20, -1.28498e-20, -1.541976e-20, 
    2.569961e-21, 5.139921e-21, 2.569961e-20, 2.312965e-20, 5.139921e-21, 
    2.569961e-21, 2.055969e-20, -2.569961e-21, 1.003089e-36, 1.003089e-36, 
    -2.312965e-20, -2.569961e-21, -1.541976e-20, -1.003089e-36, 
    -2.569961e-21, -1.28498e-20, 2.569961e-21, -1.28498e-20, -7.709882e-21, 
    5.139921e-21, -1.28498e-20, -2.569961e-20, 5.139921e-21, -1.541976e-20, 
    0, -1.541976e-20, 2.569961e-21, 1.28498e-20, -7.709882e-21, 
    -2.312965e-20, 7.709882e-21, 1.28498e-20, 1.027984e-20, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, 1.798972e-20, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 1.541976e-20, -7.709882e-21, -7.709882e-21, 
    -2.312965e-20, 0, -2.569961e-21, 5.139921e-21, 1.003089e-36, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 1.541976e-20, 1.28498e-20, -2.569961e-21, -1.027984e-20, 
    1.541976e-20, -1.541976e-20, 5.139921e-21, 1.027984e-20, 0, 
    -1.027984e-20, -1.027984e-20, 1.798972e-20, -1.027984e-20,
  6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.153676e-12, 5.176412e-12, 5.171992e-12, 5.19033e-12, 5.180158e-12, 
    5.192165e-12, 5.158286e-12, 5.177314e-12, 5.165167e-12, 5.155724e-12, 
    5.225918e-12, 5.191148e-12, 5.262042e-12, 5.239865e-12, 5.29558e-12, 
    5.25859e-12, 5.303038e-12, 5.294514e-12, 5.320175e-12, 5.312823e-12, 
    5.345644e-12, 5.323568e-12, 5.362661e-12, 5.340373e-12, 5.343859e-12, 
    5.322839e-12, 5.198146e-12, 5.221588e-12, 5.196757e-12, 5.2001e-12, 
    5.1986e-12, 5.180368e-12, 5.171179e-12, 5.151939e-12, 5.155433e-12, 
    5.169564e-12, 5.201603e-12, 5.190728e-12, 5.218139e-12, 5.21752e-12, 
    5.248038e-12, 5.234278e-12, 5.285576e-12, 5.270996e-12, 5.31313e-12, 
    5.302533e-12, 5.312632e-12, 5.30957e-12, 5.312672e-12, 5.297131e-12, 
    5.303789e-12, 5.290114e-12, 5.236855e-12, 5.252506e-12, 5.205827e-12, 
    5.177759e-12, 5.159121e-12, 5.145894e-12, 5.147763e-12, 5.151328e-12, 
    5.169646e-12, 5.186871e-12, 5.199998e-12, 5.208779e-12, 5.217431e-12, 
    5.243618e-12, 5.257482e-12, 5.288524e-12, 5.282923e-12, 5.292412e-12, 
    5.301479e-12, 5.316701e-12, 5.314196e-12, 5.320902e-12, 5.292163e-12, 
    5.311262e-12, 5.279732e-12, 5.288355e-12, 5.219779e-12, 5.193662e-12, 
    5.182558e-12, 5.172842e-12, 5.149201e-12, 5.165526e-12, 5.159091e-12, 
    5.174403e-12, 5.184132e-12, 5.17932e-12, 5.209019e-12, 5.197473e-12, 
    5.258304e-12, 5.232101e-12, 5.300422e-12, 5.284072e-12, 5.30434e-12, 
    5.293998e-12, 5.311719e-12, 5.29577e-12, 5.323398e-12, 5.329414e-12, 
    5.325303e-12, 5.341097e-12, 5.294886e-12, 5.312632e-12, 5.179185e-12, 
    5.17997e-12, 5.183626e-12, 5.167554e-12, 5.166571e-12, 5.151843e-12, 
    5.164948e-12, 5.170529e-12, 5.184696e-12, 5.193076e-12, 5.201042e-12, 
    5.218557e-12, 5.238119e-12, 5.265476e-12, 5.285132e-12, 5.298307e-12, 
    5.290229e-12, 5.297361e-12, 5.289388e-12, 5.285651e-12, 5.32716e-12, 
    5.303851e-12, 5.338825e-12, 5.33689e-12, 5.321062e-12, 5.337108e-12, 
    5.180521e-12, 5.176005e-12, 5.160325e-12, 5.172596e-12, 5.15024e-12, 
    5.162753e-12, 5.169948e-12, 5.197713e-12, 5.203814e-12, 5.209471e-12, 
    5.220644e-12, 5.234982e-12, 5.260137e-12, 5.282024e-12, 5.302007e-12, 
    5.300543e-12, 5.301058e-12, 5.305522e-12, 5.294465e-12, 5.307337e-12, 
    5.309497e-12, 5.303849e-12, 5.336631e-12, 5.327265e-12, 5.336849e-12, 
    5.330751e-12, 5.177473e-12, 5.185072e-12, 5.180965e-12, 5.188687e-12, 
    5.183247e-12, 5.207436e-12, 5.214689e-12, 5.248628e-12, 5.2347e-12, 
    5.256868e-12, 5.236952e-12, 5.24048e-12, 5.257589e-12, 5.238028e-12, 
    5.280817e-12, 5.251806e-12, 5.305695e-12, 5.276722e-12, 5.307511e-12, 
    5.30192e-12, 5.311177e-12, 5.319467e-12, 5.329897e-12, 5.349142e-12, 
    5.344686e-12, 5.360781e-12, 5.196401e-12, 5.206257e-12, 5.20539e-12, 
    5.215705e-12, 5.223334e-12, 5.239871e-12, 5.266393e-12, 5.256419e-12, 
    5.27473e-12, 5.278406e-12, 5.250588e-12, 5.267667e-12, 5.212854e-12, 
    5.221709e-12, 5.216437e-12, 5.197178e-12, 5.258717e-12, 5.227133e-12, 
    5.285457e-12, 5.268346e-12, 5.318285e-12, 5.293448e-12, 5.342232e-12, 
    5.363087e-12, 5.382719e-12, 5.405658e-12, 5.211637e-12, 5.20494e-12, 
    5.216932e-12, 5.233524e-12, 5.248921e-12, 5.269389e-12, 5.271484e-12, 
    5.275319e-12, 5.285252e-12, 5.293604e-12, 5.276531e-12, 5.295697e-12, 
    5.223761e-12, 5.261458e-12, 5.202408e-12, 5.220187e-12, 5.232546e-12, 
    5.227125e-12, 5.25528e-12, 5.261915e-12, 5.288881e-12, 5.274942e-12, 
    5.357939e-12, 5.321217e-12, 5.423127e-12, 5.394645e-12, 5.2026e-12, 
    5.211615e-12, 5.242989e-12, 5.228061e-12, 5.270756e-12, 5.281266e-12, 
    5.28981e-12, 5.300732e-12, 5.301911e-12, 5.308382e-12, 5.297778e-12, 
    5.307964e-12, 5.269433e-12, 5.286651e-12, 5.239404e-12, 5.250903e-12, 
    5.245613e-12, 5.23981e-12, 5.257719e-12, 5.276799e-12, 5.277208e-12, 
    5.283326e-12, 5.300564e-12, 5.27093e-12, 5.362676e-12, 5.306012e-12, 
    5.221445e-12, 5.238808e-12, 5.241289e-12, 5.234563e-12, 5.280212e-12, 
    5.263671e-12, 5.308225e-12, 5.296183e-12, 5.315913e-12, 5.306109e-12, 
    5.304666e-12, 5.292075e-12, 5.284235e-12, 5.26443e-12, 5.248315e-12, 
    5.235539e-12, 5.23851e-12, 5.252545e-12, 5.277966e-12, 5.302018e-12, 
    5.296749e-12, 5.314414e-12, 5.26766e-12, 5.287264e-12, 5.279686e-12, 
    5.299444e-12, 5.256154e-12, 5.293014e-12, 5.246732e-12, 5.25079e-12, 
    5.263343e-12, 5.288592e-12, 5.294181e-12, 5.300146e-12, 5.296465e-12, 
    5.278612e-12, 5.275687e-12, 5.263038e-12, 5.259545e-12, 5.249907e-12, 
    5.241927e-12, 5.249218e-12, 5.256874e-12, 5.27862e-12, 5.298217e-12, 
    5.319585e-12, 5.324814e-12, 5.349779e-12, 5.329455e-12, 5.362992e-12, 
    5.334477e-12, 5.383841e-12, 5.295152e-12, 5.333641e-12, 5.263914e-12, 
    5.271426e-12, 5.285012e-12, 5.316174e-12, 5.299352e-12, 5.319026e-12, 
    5.275573e-12, 5.253028e-12, 5.247197e-12, 5.236315e-12, 5.247446e-12, 
    5.246541e-12, 5.257192e-12, 5.253769e-12, 5.279342e-12, 5.265605e-12, 
    5.30463e-12, 5.318871e-12, 5.359093e-12, 5.383752e-12, 5.408856e-12, 
    5.419938e-12, 5.423312e-12, 5.424722e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.117974e-11, 3.131729e-11, 3.129055e-11, 3.14015e-11, 3.133995e-11, 
    3.14126e-11, 3.120763e-11, 3.132275e-11, 3.124926e-11, 3.119213e-11, 
    3.16168e-11, 3.140645e-11, 3.183535e-11, 3.170118e-11, 3.203825e-11, 
    3.181447e-11, 3.208338e-11, 3.203181e-11, 3.218706e-11, 3.214258e-11, 
    3.234115e-11, 3.220759e-11, 3.24441e-11, 3.230926e-11, 3.233035e-11, 
    3.220318e-11, 3.144878e-11, 3.159061e-11, 3.144038e-11, 3.14606e-11, 
    3.145153e-11, 3.134122e-11, 3.128563e-11, 3.116923e-11, 3.119037e-11, 
    3.127586e-11, 3.14697e-11, 3.14039e-11, 3.156974e-11, 3.1566e-11, 
    3.175063e-11, 3.166738e-11, 3.197773e-11, 3.188953e-11, 3.214444e-11, 
    3.208033e-11, 3.214142e-11, 3.21229e-11, 3.214166e-11, 3.204764e-11, 
    3.208793e-11, 3.200519e-11, 3.168297e-11, 3.177766e-11, 3.149525e-11, 
    3.132544e-11, 3.121268e-11, 3.113266e-11, 3.114397e-11, 3.116553e-11, 
    3.127636e-11, 3.138057e-11, 3.145999e-11, 3.151311e-11, 3.156546e-11, 
    3.172389e-11, 3.180777e-11, 3.199557e-11, 3.196168e-11, 3.201909e-11, 
    3.207395e-11, 3.216604e-11, 3.215089e-11, 3.219146e-11, 3.201758e-11, 
    3.213314e-11, 3.194238e-11, 3.199455e-11, 3.157967e-11, 3.142165e-11, 
    3.135447e-11, 3.129569e-11, 3.115267e-11, 3.125144e-11, 3.12125e-11, 
    3.130514e-11, 3.1364e-11, 3.133489e-11, 3.151457e-11, 3.144471e-11, 
    3.181274e-11, 3.165421e-11, 3.206755e-11, 3.196864e-11, 3.209126e-11, 
    3.202869e-11, 3.21359e-11, 3.203941e-11, 3.220656e-11, 3.224296e-11, 
    3.221809e-11, 3.231363e-11, 3.203406e-11, 3.214142e-11, 3.133407e-11, 
    3.133882e-11, 3.136094e-11, 3.12637e-11, 3.125775e-11, 3.116865e-11, 
    3.124793e-11, 3.12817e-11, 3.136741e-11, 3.141811e-11, 3.146631e-11, 
    3.157227e-11, 3.169062e-11, 3.185613e-11, 3.197505e-11, 3.205476e-11, 
    3.200588e-11, 3.204903e-11, 3.200079e-11, 3.197819e-11, 3.222932e-11, 
    3.20883e-11, 3.229989e-11, 3.228819e-11, 3.219242e-11, 3.22895e-11, 
    3.134215e-11, 3.131483e-11, 3.121996e-11, 3.12942e-11, 3.115895e-11, 
    3.123465e-11, 3.127818e-11, 3.144616e-11, 3.148308e-11, 3.15173e-11, 
    3.158489e-11, 3.167164e-11, 3.182382e-11, 3.195625e-11, 3.207714e-11, 
    3.206828e-11, 3.20714e-11, 3.209841e-11, 3.203151e-11, 3.210939e-11, 
    3.212246e-11, 3.208829e-11, 3.228662e-11, 3.222995e-11, 3.228794e-11, 
    3.225104e-11, 3.132371e-11, 3.136968e-11, 3.134484e-11, 3.139156e-11, 
    3.135864e-11, 3.150499e-11, 3.154887e-11, 3.17542e-11, 3.166993e-11, 
    3.180405e-11, 3.168356e-11, 3.170491e-11, 3.180841e-11, 3.169007e-11, 
    3.194894e-11, 3.177342e-11, 3.209946e-11, 3.192417e-11, 3.211044e-11, 
    3.207662e-11, 3.213262e-11, 3.218277e-11, 3.224588e-11, 3.236231e-11, 
    3.233535e-11, 3.243272e-11, 3.143823e-11, 3.149786e-11, 3.149261e-11, 
    3.155502e-11, 3.160117e-11, 3.170122e-11, 3.186168e-11, 3.180134e-11, 
    3.191212e-11, 3.193436e-11, 3.176606e-11, 3.186939e-11, 3.153777e-11, 
    3.159134e-11, 3.155945e-11, 3.144293e-11, 3.181523e-11, 3.162416e-11, 
    3.197701e-11, 3.187349e-11, 3.217562e-11, 3.202536e-11, 3.232051e-11, 
    3.244667e-11, 3.256545e-11, 3.270423e-11, 3.15304e-11, 3.148989e-11, 
    3.156244e-11, 3.166282e-11, 3.175597e-11, 3.18798e-11, 3.189248e-11, 
    3.191568e-11, 3.197578e-11, 3.202631e-11, 3.192301e-11, 3.203897e-11, 
    3.160375e-11, 3.183183e-11, 3.147456e-11, 3.158213e-11, 3.16569e-11, 
    3.162411e-11, 3.179444e-11, 3.183459e-11, 3.199773e-11, 3.19134e-11, 
    3.241553e-11, 3.219336e-11, 3.280992e-11, 3.26376e-11, 3.147573e-11, 
    3.153027e-11, 3.172008e-11, 3.162977e-11, 3.188808e-11, 3.195166e-11, 
    3.200335e-11, 3.206943e-11, 3.207656e-11, 3.211571e-11, 3.205156e-11, 
    3.211318e-11, 3.188007e-11, 3.198424e-11, 3.169839e-11, 3.176796e-11, 
    3.173596e-11, 3.170085e-11, 3.18092e-11, 3.192463e-11, 3.192711e-11, 
    3.196412e-11, 3.206841e-11, 3.188912e-11, 3.244419e-11, 3.210137e-11, 
    3.158974e-11, 3.169479e-11, 3.17098e-11, 3.16691e-11, 3.194528e-11, 
    3.184521e-11, 3.211476e-11, 3.204191e-11, 3.216127e-11, 3.210196e-11, 
    3.209323e-11, 3.201705e-11, 3.196962e-11, 3.18498e-11, 3.175231e-11, 
    3.167501e-11, 3.169298e-11, 3.17779e-11, 3.19317e-11, 3.207721e-11, 
    3.204533e-11, 3.21522e-11, 3.186934e-11, 3.198795e-11, 3.194211e-11, 
    3.206164e-11, 3.179973e-11, 3.202274e-11, 3.174273e-11, 3.176728e-11, 
    3.184322e-11, 3.199599e-11, 3.20298e-11, 3.206588e-11, 3.204361e-11, 
    3.19356e-11, 3.191791e-11, 3.184138e-11, 3.182025e-11, 3.176194e-11, 
    3.171366e-11, 3.175777e-11, 3.180409e-11, 3.193565e-11, 3.205421e-11, 
    3.218349e-11, 3.221513e-11, 3.236616e-11, 3.22432e-11, 3.24461e-11, 
    3.227359e-11, 3.257224e-11, 3.203567e-11, 3.226852e-11, 3.184668e-11, 
    3.189213e-11, 3.197432e-11, 3.216286e-11, 3.206108e-11, 3.218011e-11, 
    3.191722e-11, 3.178082e-11, 3.174554e-11, 3.167971e-11, 3.174705e-11, 
    3.174157e-11, 3.180601e-11, 3.17853e-11, 3.194002e-11, 3.185691e-11, 
    3.209301e-11, 3.217917e-11, 3.242252e-11, 3.25717e-11, 3.272358e-11, 
    3.279063e-11, 3.281104e-11, 3.281957e-11 ;

 SOILC =
  17.34481, 17.34479, 17.3448, 17.34479, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.34481, 17.34476, 17.34479, 17.34474, 17.34476, 
    17.34472, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34471, 17.34472, 17.34471, 17.34473, 17.34472, 17.34473, 
    17.34473, 17.34477, 17.34478, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.3448, 17.3448, 17.34479, 17.34479, 17.34477, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34472, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.3448, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.3447, 17.34471, 17.34479, 17.34479, 17.34479, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34475, 17.34476, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34476, 17.34473, 17.34475, 17.34472, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 17.3447, 17.34469, 
    17.34478, 17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 
    17.34475, 17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 
    17.34477, 17.34478, 17.34475, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34473, 17.3447, 17.34469, 17.34468, 17.34466, 17.34477, 17.34478, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34474, 17.34473, 
    17.34473, 17.34474, 17.34472, 17.34477, 17.34475, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 
    17.34471, 17.34465, 17.34467, 17.34478, 17.34477, 17.34476, 17.34476, 
    17.34474, 17.34473, 17.34473, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34474, 17.34473, 17.34476, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 
    17.34472, 17.34477, 17.34476, 17.34476, 17.34476, 17.34473, 17.34474, 
    17.34472, 17.34472, 17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34474, 17.34473, 17.34473, 17.34472, 17.34475, 
    17.34473, 17.34475, 17.34475, 17.34474, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34469, 17.3447, 17.34468, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34474, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34475, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 SOILC_HR =
  6.195739e-08, 6.223058e-08, 6.217748e-08, 6.239782e-08, 6.22756e-08, 
    6.241988e-08, 6.201279e-08, 6.224143e-08, 6.209547e-08, 6.198199e-08, 
    6.282544e-08, 6.240766e-08, 6.325951e-08, 6.299303e-08, 6.36625e-08, 
    6.321804e-08, 6.375213e-08, 6.364969e-08, 6.395803e-08, 6.38697e-08, 
    6.426407e-08, 6.39988e-08, 6.446854e-08, 6.420073e-08, 6.424262e-08, 
    6.399005e-08, 6.249174e-08, 6.277342e-08, 6.247505e-08, 6.251522e-08, 
    6.24972e-08, 6.227812e-08, 6.216771e-08, 6.193653e-08, 6.19785e-08, 
    6.21483e-08, 6.253328e-08, 6.240261e-08, 6.273198e-08, 6.272454e-08, 
    6.309124e-08, 6.29259e-08, 6.354229e-08, 6.33671e-08, 6.387339e-08, 
    6.374605e-08, 6.38674e-08, 6.38306e-08, 6.386788e-08, 6.368114e-08, 
    6.376114e-08, 6.359683e-08, 6.295686e-08, 6.314493e-08, 6.258403e-08, 
    6.224678e-08, 6.202281e-08, 6.186388e-08, 6.188635e-08, 6.192918e-08, 
    6.21493e-08, 6.235626e-08, 6.2514e-08, 6.261951e-08, 6.272347e-08, 
    6.303814e-08, 6.320472e-08, 6.357771e-08, 6.351041e-08, 6.362443e-08, 
    6.373339e-08, 6.39163e-08, 6.388619e-08, 6.396677e-08, 6.362144e-08, 
    6.385094e-08, 6.347207e-08, 6.357569e-08, 6.275169e-08, 6.243786e-08, 
    6.230444e-08, 6.218769e-08, 6.190362e-08, 6.209979e-08, 6.202245e-08, 
    6.220644e-08, 6.232334e-08, 6.226553e-08, 6.262239e-08, 6.248365e-08, 
    6.321459e-08, 6.289974e-08, 6.372068e-08, 6.352423e-08, 6.376777e-08, 
    6.36435e-08, 6.385643e-08, 6.366479e-08, 6.399677e-08, 6.406906e-08, 
    6.401966e-08, 6.420943e-08, 6.365416e-08, 6.38674e-08, 6.226391e-08, 
    6.227334e-08, 6.231727e-08, 6.212414e-08, 6.211233e-08, 6.193537e-08, 
    6.209284e-08, 6.215989e-08, 6.233013e-08, 6.243081e-08, 6.252654e-08, 
    6.273701e-08, 6.297206e-08, 6.330077e-08, 6.353696e-08, 6.369527e-08, 
    6.35982e-08, 6.368391e-08, 6.35881e-08, 6.354319e-08, 6.404196e-08, 
    6.376189e-08, 6.418213e-08, 6.415888e-08, 6.396869e-08, 6.41615e-08, 
    6.227996e-08, 6.222569e-08, 6.203729e-08, 6.218473e-08, 6.19161e-08, 
    6.206646e-08, 6.215291e-08, 6.248654e-08, 6.255986e-08, 6.262782e-08, 
    6.276207e-08, 6.293436e-08, 6.323661e-08, 6.349962e-08, 6.373973e-08, 
    6.372213e-08, 6.372833e-08, 6.378196e-08, 6.36491e-08, 6.380377e-08, 
    6.382973e-08, 6.376186e-08, 6.415576e-08, 6.404323e-08, 6.415839e-08, 
    6.408511e-08, 6.224334e-08, 6.233464e-08, 6.22853e-08, 6.237808e-08, 
    6.231271e-08, 6.260337e-08, 6.269052e-08, 6.309833e-08, 6.293097e-08, 
    6.319734e-08, 6.295803e-08, 6.300043e-08, 6.320601e-08, 6.297097e-08, 
    6.348511e-08, 6.313651e-08, 6.378404e-08, 6.343591e-08, 6.380586e-08, 
    6.373869e-08, 6.384992e-08, 6.394953e-08, 6.407485e-08, 6.43061e-08, 
    6.425255e-08, 6.444595e-08, 6.247078e-08, 6.25892e-08, 6.257878e-08, 
    6.270273e-08, 6.27944e-08, 6.29931e-08, 6.331179e-08, 6.319195e-08, 
    6.341197e-08, 6.345614e-08, 6.312188e-08, 6.33271e-08, 6.266848e-08, 
    6.277487e-08, 6.271153e-08, 6.248011e-08, 6.321955e-08, 6.284005e-08, 
    6.354086e-08, 6.333526e-08, 6.393532e-08, 6.363688e-08, 6.422307e-08, 
    6.447366e-08, 6.470955e-08, 6.498519e-08, 6.265385e-08, 6.257338e-08, 
    6.271748e-08, 6.291684e-08, 6.310184e-08, 6.33478e-08, 6.337297e-08, 
    6.341904e-08, 6.35384e-08, 6.363876e-08, 6.34336e-08, 6.366392e-08, 
    6.279953e-08, 6.32525e-08, 6.254295e-08, 6.275658e-08, 6.290509e-08, 
    6.283995e-08, 6.317826e-08, 6.325799e-08, 6.358201e-08, 6.341452e-08, 
    6.44118e-08, 6.397055e-08, 6.51951e-08, 6.485286e-08, 6.254526e-08, 
    6.265358e-08, 6.303058e-08, 6.28512e-08, 6.336422e-08, 6.34905e-08, 
    6.359317e-08, 6.37244e-08, 6.373858e-08, 6.381633e-08, 6.368892e-08, 
    6.38113e-08, 6.334832e-08, 6.355521e-08, 6.298749e-08, 6.312566e-08, 
    6.30621e-08, 6.299238e-08, 6.320757e-08, 6.343683e-08, 6.344175e-08, 
    6.351525e-08, 6.372239e-08, 6.33663e-08, 6.446873e-08, 6.378785e-08, 
    6.27717e-08, 6.298033e-08, 6.301015e-08, 6.292932e-08, 6.347784e-08, 
    6.327909e-08, 6.381444e-08, 6.366975e-08, 6.390682e-08, 6.378902e-08, 
    6.377169e-08, 6.362038e-08, 6.352618e-08, 6.32882e-08, 6.309457e-08, 
    6.294105e-08, 6.297675e-08, 6.314539e-08, 6.345086e-08, 6.373985e-08, 
    6.367654e-08, 6.388881e-08, 6.332702e-08, 6.356257e-08, 6.347153e-08, 
    6.370894e-08, 6.318876e-08, 6.363167e-08, 6.307555e-08, 6.312431e-08, 
    6.327515e-08, 6.357854e-08, 6.364569e-08, 6.371736e-08, 6.367314e-08, 
    6.345861e-08, 6.342348e-08, 6.327148e-08, 6.322951e-08, 6.31137e-08, 
    6.301781e-08, 6.310542e-08, 6.319741e-08, 6.345871e-08, 6.369419e-08, 
    6.395094e-08, 6.401378e-08, 6.431375e-08, 6.406955e-08, 6.447252e-08, 
    6.412989e-08, 6.472303e-08, 6.365737e-08, 6.411983e-08, 6.328201e-08, 
    6.337227e-08, 6.353551e-08, 6.390996e-08, 6.370782e-08, 6.394423e-08, 
    6.34221e-08, 6.315121e-08, 6.308114e-08, 6.295038e-08, 6.308413e-08, 
    6.307325e-08, 6.320123e-08, 6.316011e-08, 6.346739e-08, 6.330233e-08, 
    6.377125e-08, 6.394237e-08, 6.442568e-08, 6.472197e-08, 6.502361e-08, 
    6.515678e-08, 6.519732e-08, 6.521426e-08 ;

 SOILC_LOSS =
  6.195739e-08, 6.223058e-08, 6.217748e-08, 6.239782e-08, 6.22756e-08, 
    6.241988e-08, 6.201279e-08, 6.224143e-08, 6.209547e-08, 6.198199e-08, 
    6.282544e-08, 6.240766e-08, 6.325951e-08, 6.299303e-08, 6.36625e-08, 
    6.321804e-08, 6.375213e-08, 6.364969e-08, 6.395803e-08, 6.38697e-08, 
    6.426407e-08, 6.39988e-08, 6.446854e-08, 6.420073e-08, 6.424262e-08, 
    6.399005e-08, 6.249174e-08, 6.277342e-08, 6.247505e-08, 6.251522e-08, 
    6.24972e-08, 6.227812e-08, 6.216771e-08, 6.193653e-08, 6.19785e-08, 
    6.21483e-08, 6.253328e-08, 6.240261e-08, 6.273198e-08, 6.272454e-08, 
    6.309124e-08, 6.29259e-08, 6.354229e-08, 6.33671e-08, 6.387339e-08, 
    6.374605e-08, 6.38674e-08, 6.38306e-08, 6.386788e-08, 6.368114e-08, 
    6.376114e-08, 6.359683e-08, 6.295686e-08, 6.314493e-08, 6.258403e-08, 
    6.224678e-08, 6.202281e-08, 6.186388e-08, 6.188635e-08, 6.192918e-08, 
    6.21493e-08, 6.235626e-08, 6.2514e-08, 6.261951e-08, 6.272347e-08, 
    6.303814e-08, 6.320472e-08, 6.357771e-08, 6.351041e-08, 6.362443e-08, 
    6.373339e-08, 6.39163e-08, 6.388619e-08, 6.396677e-08, 6.362144e-08, 
    6.385094e-08, 6.347207e-08, 6.357569e-08, 6.275169e-08, 6.243786e-08, 
    6.230444e-08, 6.218769e-08, 6.190362e-08, 6.209979e-08, 6.202245e-08, 
    6.220644e-08, 6.232334e-08, 6.226553e-08, 6.262239e-08, 6.248365e-08, 
    6.321459e-08, 6.289974e-08, 6.372068e-08, 6.352423e-08, 6.376777e-08, 
    6.36435e-08, 6.385643e-08, 6.366479e-08, 6.399677e-08, 6.406906e-08, 
    6.401966e-08, 6.420943e-08, 6.365416e-08, 6.38674e-08, 6.226391e-08, 
    6.227334e-08, 6.231727e-08, 6.212414e-08, 6.211233e-08, 6.193537e-08, 
    6.209284e-08, 6.215989e-08, 6.233013e-08, 6.243081e-08, 6.252654e-08, 
    6.273701e-08, 6.297206e-08, 6.330077e-08, 6.353696e-08, 6.369527e-08, 
    6.35982e-08, 6.368391e-08, 6.35881e-08, 6.354319e-08, 6.404196e-08, 
    6.376189e-08, 6.418213e-08, 6.415888e-08, 6.396869e-08, 6.41615e-08, 
    6.227996e-08, 6.222569e-08, 6.203729e-08, 6.218473e-08, 6.19161e-08, 
    6.206646e-08, 6.215291e-08, 6.248654e-08, 6.255986e-08, 6.262782e-08, 
    6.276207e-08, 6.293436e-08, 6.323661e-08, 6.349962e-08, 6.373973e-08, 
    6.372213e-08, 6.372833e-08, 6.378196e-08, 6.36491e-08, 6.380377e-08, 
    6.382973e-08, 6.376186e-08, 6.415576e-08, 6.404323e-08, 6.415839e-08, 
    6.408511e-08, 6.224334e-08, 6.233464e-08, 6.22853e-08, 6.237808e-08, 
    6.231271e-08, 6.260337e-08, 6.269052e-08, 6.309833e-08, 6.293097e-08, 
    6.319734e-08, 6.295803e-08, 6.300043e-08, 6.320601e-08, 6.297097e-08, 
    6.348511e-08, 6.313651e-08, 6.378404e-08, 6.343591e-08, 6.380586e-08, 
    6.373869e-08, 6.384992e-08, 6.394953e-08, 6.407485e-08, 6.43061e-08, 
    6.425255e-08, 6.444595e-08, 6.247078e-08, 6.25892e-08, 6.257878e-08, 
    6.270273e-08, 6.27944e-08, 6.29931e-08, 6.331179e-08, 6.319195e-08, 
    6.341197e-08, 6.345614e-08, 6.312188e-08, 6.33271e-08, 6.266848e-08, 
    6.277487e-08, 6.271153e-08, 6.248011e-08, 6.321955e-08, 6.284005e-08, 
    6.354086e-08, 6.333526e-08, 6.393532e-08, 6.363688e-08, 6.422307e-08, 
    6.447366e-08, 6.470955e-08, 6.498519e-08, 6.265385e-08, 6.257338e-08, 
    6.271748e-08, 6.291684e-08, 6.310184e-08, 6.33478e-08, 6.337297e-08, 
    6.341904e-08, 6.35384e-08, 6.363876e-08, 6.34336e-08, 6.366392e-08, 
    6.279953e-08, 6.32525e-08, 6.254295e-08, 6.275658e-08, 6.290509e-08, 
    6.283995e-08, 6.317826e-08, 6.325799e-08, 6.358201e-08, 6.341452e-08, 
    6.44118e-08, 6.397055e-08, 6.51951e-08, 6.485286e-08, 6.254526e-08, 
    6.265358e-08, 6.303058e-08, 6.28512e-08, 6.336422e-08, 6.34905e-08, 
    6.359317e-08, 6.37244e-08, 6.373858e-08, 6.381633e-08, 6.368892e-08, 
    6.38113e-08, 6.334832e-08, 6.355521e-08, 6.298749e-08, 6.312566e-08, 
    6.30621e-08, 6.299238e-08, 6.320757e-08, 6.343683e-08, 6.344175e-08, 
    6.351525e-08, 6.372239e-08, 6.33663e-08, 6.446873e-08, 6.378785e-08, 
    6.27717e-08, 6.298033e-08, 6.301015e-08, 6.292932e-08, 6.347784e-08, 
    6.327909e-08, 6.381444e-08, 6.366975e-08, 6.390682e-08, 6.378902e-08, 
    6.377169e-08, 6.362038e-08, 6.352618e-08, 6.32882e-08, 6.309457e-08, 
    6.294105e-08, 6.297675e-08, 6.314539e-08, 6.345086e-08, 6.373985e-08, 
    6.367654e-08, 6.388881e-08, 6.332702e-08, 6.356257e-08, 6.347153e-08, 
    6.370894e-08, 6.318876e-08, 6.363167e-08, 6.307555e-08, 6.312431e-08, 
    6.327515e-08, 6.357854e-08, 6.364569e-08, 6.371736e-08, 6.367314e-08, 
    6.345861e-08, 6.342348e-08, 6.327148e-08, 6.322951e-08, 6.31137e-08, 
    6.301781e-08, 6.310542e-08, 6.319741e-08, 6.345871e-08, 6.369419e-08, 
    6.395094e-08, 6.401378e-08, 6.431375e-08, 6.406955e-08, 6.447252e-08, 
    6.412989e-08, 6.472303e-08, 6.365737e-08, 6.411983e-08, 6.328201e-08, 
    6.337227e-08, 6.353551e-08, 6.390996e-08, 6.370782e-08, 6.394423e-08, 
    6.34221e-08, 6.315121e-08, 6.308114e-08, 6.295038e-08, 6.308413e-08, 
    6.307325e-08, 6.320123e-08, 6.316011e-08, 6.346739e-08, 6.330233e-08, 
    6.377125e-08, 6.394237e-08, 6.442568e-08, 6.472197e-08, 6.502361e-08, 
    6.515678e-08, 6.519732e-08, 6.521426e-08 ;

 SOILICE =
  96.3256, 96.77938, 96.69106, 97.05782, 96.85425, 97.09457, 96.41747, 
    96.79745, 96.55476, 96.36636, 97.77205, 97.0742, 98.49985, 98.05251, 
    99.17845, 98.43019, 99.32972, 99.15676, 99.67771, 99.52831, 100.1965, 
    99.74671, 100.5438, 100.0889, 100.16, 99.7319, 97.21435, 97.68502, 
    97.18652, 97.25353, 97.22344, 96.85847, 96.67489, 96.29093, 96.36056, 
    96.64258, 97.28368, 97.06573, 97.61546, 97.60303, 98.21721, 97.94, 
    98.97568, 98.68066, 99.53454, 99.3194, 99.52444, 99.46223, 99.52525, 
    99.20983, 99.3449, 99.0676, 97.9919, 98.30733, 97.36835, 96.80642, 
    96.43413, 96.17051, 96.20775, 96.27878, 96.64423, 96.98854, 97.25144, 
    97.42754, 97.60124, 98.12828, 98.40778, 99.03542, 98.92194, 99.1142, 
    99.29801, 99.60712, 99.5562, 99.69254, 99.10909, 99.49664, 98.85733, 
    99.03196, 97.64868, 97.12449, 96.90236, 96.70804, 96.2364, 96.56196, 
    96.43355, 96.73918, 96.93372, 96.83747, 97.43236, 97.20083, 98.42437, 
    97.89623, 99.27656, 98.94521, 99.35607, 99.14629, 99.50591, 99.18221, 
    99.74329, 99.86573, 99.78205, 100.1036, 99.1643, 99.52445, 96.83479, 
    96.85048, 96.9236, 96.60244, 96.5828, 96.28903, 96.55038, 96.66182, 
    96.94499, 97.11275, 97.27238, 97.62389, 98.0174, 98.56918, 98.96667, 
    99.23367, 99.06989, 99.21447, 99.05286, 98.97716, 99.81985, 99.34617, 
    100.0573, 100.0179, 99.69579, 100.0224, 96.8615, 96.77119, 96.45815, 
    96.70309, 96.25707, 96.5066, 96.65026, 97.20571, 97.32796, 97.44145, 
    97.66579, 97.95419, 98.46132, 98.90379, 99.3087, 99.279, 99.28945, 
    99.38005, 99.15575, 99.4169, 99.46078, 99.34609, 100.0126, 99.82194, 
    100.0171, 99.89288, 96.80054, 96.95253, 96.87038, 97.02489, 96.91604, 
    97.40068, 97.54626, 98.22916, 97.94851, 98.39535, 97.99384, 98.06492, 
    98.41003, 98.0155, 98.8794, 98.29328, 99.38358, 98.7966, 99.42043, 
    99.30695, 99.49486, 99.66335, 99.87551, 100.2677, 100.1768, 100.5053, 
    97.17935, 97.377, 97.35955, 97.56659, 97.71989, 98.0526, 98.58766, 
    98.38624, 98.75616, 98.83054, 98.26859, 98.61343, 97.50938, 97.68729, 
    97.58131, 97.19495, 98.43269, 97.79634, 98.97326, 98.62711, 99.63932, 
    99.13521, 100.1268, 100.5525, 100.954, 101.4245, 97.48492, 97.35052, 
    97.59122, 97.9249, 98.23499, 98.64821, 98.69052, 98.76808, 98.96909, 
    99.1383, 98.79264, 99.18074, 97.72865, 98.48801, 97.29977, 97.65672, 
    97.90519, 97.79611, 98.36323, 98.49718, 99.04266, 98.76044, 100.4474, 
    99.69901, 101.7834, 101.1985, 97.3036, 97.48444, 98.11548, 97.81493, 
    98.67581, 98.88841, 99.06141, 99.28287, 99.30677, 99.43813, 99.22292, 
    99.42961, 98.64909, 98.99744, 98.04318, 98.27496, 98.16828, 98.05137, 
    98.41247, 98.79809, 98.80628, 98.93014, 99.27974, 98.67931, 100.5443, 
    99.39025, 97.68188, 98.0313, 98.08119, 97.94572, 98.86709, 98.53266, 
    99.43492, 99.19059, 99.59109, 99.39196, 99.36269, 99.1073, 98.94852, 
    98.548, 98.2228, 97.96535, 98.02518, 98.3081, 98.82169, 99.30896, 
    99.20211, 99.56062, 98.61324, 99.00988, 98.85649, 99.25674, 98.38091, 
    99.12662, 98.19085, 98.27267, 98.52603, 99.03686, 99.14999, 99.27098, 
    99.1963, 98.83474, 98.77555, 98.51986, 98.44936, 98.25485, 98.09402, 
    98.24097, 98.39545, 98.83487, 99.23187, 99.66576, 99.77208, 100.2809, 
    99.86666, 100.5508, 99.96911, 100.9772, 99.16985, 99.95191, 98.53755, 
    98.68935, 98.9643, 99.59651, 99.25485, 99.65446, 98.77323, 98.3179, 
    98.20022, 97.981, 98.20524, 98.18699, 98.40181, 98.33274, 98.84948, 
    98.57171, 99.36197, 99.65128, 100.4709, 100.9753, 101.4901, 101.7178, 
    101.7872, 101.8162,
  95.28641, 95.75723, 95.66557, 96.0462, 95.8349, 96.08433, 95.3817, 
    95.77599, 95.52415, 95.32867, 96.78765, 96.06319, 97.54329, 97.07873, 
    98.24815, 97.47096, 98.4053, 98.22558, 98.76684, 98.61159, 99.30606, 
    98.83854, 99.66703, 99.19423, 99.26815, 98.82316, 96.20862, 96.6973, 
    96.17973, 96.24931, 96.21806, 95.83929, 95.64884, 95.25041, 95.32265, 
    95.61528, 96.2806, 96.05437, 96.62495, 96.61205, 97.24973, 96.9619, 
    98.03746, 97.73101, 98.61806, 98.39454, 98.60757, 98.54294, 98.60841, 
    98.28072, 98.42104, 98.13294, 97.01579, 97.34334, 96.36848, 95.78535, 
    95.39899, 95.12549, 95.16413, 95.23783, 95.617, 95.97426, 96.2471, 
    96.42989, 96.61019, 97.15747, 97.44768, 98.09955, 97.98163, 98.18138, 
    98.37231, 98.6935, 98.64058, 98.78226, 98.17604, 98.57872, 97.91451, 
    98.09592, 96.65959, 96.11536, 95.8849, 95.6832, 95.19385, 95.53163, 
    95.39839, 95.7155, 95.91737, 95.81748, 96.43489, 96.19458, 97.4649, 
    96.91647, 98.35004, 98.00581, 98.43263, 98.21468, 98.58834, 98.25201, 
    98.83499, 98.96225, 98.87528, 99.20949, 98.2334, 98.6076, 95.8147, 
    95.83099, 95.90686, 95.57363, 95.55325, 95.24845, 95.5196, 95.63525, 
    95.92905, 96.10317, 96.26884, 96.63373, 97.04229, 97.61526, 98.02811, 
    98.30546, 98.13531, 98.28552, 98.11763, 98.03899, 98.91458, 98.42237, 
    99.16138, 99.12038, 98.78564, 99.125, 95.84242, 95.74871, 95.4239, 
    95.67804, 95.21529, 95.47418, 95.62327, 96.19968, 96.32652, 96.44434, 
    96.67722, 96.97662, 97.50324, 97.96281, 98.38342, 98.35255, 98.36342, 
    98.45756, 98.22453, 98.49584, 98.54146, 98.42227, 99.1149, 98.91672, 
    99.11951, 98.99044, 95.77916, 95.93689, 95.85164, 96.012, 95.89903, 
    96.40205, 96.55318, 97.26219, 96.97074, 97.43474, 97.01778, 97.09161, 
    97.45004, 97.04027, 97.9375, 97.32879, 98.46122, 97.85152, 98.4995, 
    98.38159, 98.57683, 98.75192, 98.9724, 99.38008, 99.28557, 99.62703, 
    96.17229, 96.37745, 96.35931, 96.57423, 96.73338, 97.0788, 97.63445, 
    97.42525, 97.80943, 97.8867, 97.30306, 97.66122, 96.51485, 96.69958, 
    96.58952, 96.18851, 97.47353, 96.81278, 98.03496, 97.67541, 98.72696, 
    98.20322, 99.23358, 99.67619, 100.0811, 100.5555, 96.48946, 96.34994, 
    96.59979, 96.94625, 97.2682, 97.69733, 97.74126, 97.82182, 98.03061, 
    98.20639, 97.84737, 98.25048, 96.74258, 97.53098, 96.29728, 96.66785, 
    96.92577, 96.81252, 97.40134, 97.54046, 98.10706, 97.81387, 99.5669, 
    98.78902, 100.9174, 100.3277, 96.30124, 96.48895, 97.14411, 96.83204, 
    97.72598, 97.94682, 98.1265, 98.3566, 98.38142, 98.51791, 98.2943, 
    98.50905, 97.69824, 98.06007, 97.06901, 97.3097, 97.19891, 97.07751, 
    97.45248, 97.85303, 97.8615, 97.99017, 98.3535, 97.72961, 99.66777, 
    98.4683, 96.69391, 97.05673, 97.10849, 96.96782, 97.92467, 97.57732, 
    98.51456, 98.2607, 98.67683, 98.46992, 98.43951, 98.17419, 98.00925, 
    97.59325, 97.25555, 96.9882, 97.05032, 97.34412, 97.87754, 98.38371, 
    98.27271, 98.64516, 97.661, 98.07301, 97.91367, 98.32944, 97.41972, 
    98.1944, 97.22234, 97.30731, 97.57043, 98.10107, 98.21854, 98.34425, 
    98.26665, 97.89108, 97.82959, 97.56401, 97.49081, 97.2888, 97.1218, 
    97.2744, 97.43484, 97.8912, 98.30363, 98.75443, 98.8649, 99.39381, 
    98.96328, 99.67449, 99.06985, 100.1047, 98.23924, 99.05189, 97.58238, 
    97.74003, 98.02569, 98.68252, 98.32748, 98.74272, 97.82717, 97.35432, 
    97.23208, 97.00446, 97.23728, 97.21833, 97.44141, 97.36968, 97.90637, 
    97.61786, 98.43878, 98.73941, 99.59125, 100.1026, 100.6216, 100.8512, 
    100.9212, 100.9505,
  129.4638, 130.152, 130.018, 130.5745, 130.2655, 130.6302, 129.603, 
    130.1794, 129.8112, 129.5255, 131.659, 130.5993, 132.765, 132.085, 
    133.7973, 132.6591, 134.0275, 133.7642, 134.5573, 134.3298, 135.3478, 
    134.6624, 135.8772, 135.1838, 135.2922, 134.6399, 130.812, 131.5268, 
    130.7698, 130.8715, 130.8258, 130.2719, 129.9935, 129.4112, 129.5167, 
    129.9445, 130.9173, 130.5864, 131.421, 131.4021, 132.3353, 131.914, 
    133.4887, 133.0399, 134.3393, 134.0118, 134.3239, 134.2292, 134.3252, 
    133.845, 134.0506, 133.6286, 131.9929, 132.4723, 131.0458, 130.1931, 
    129.6283, 129.2286, 129.2851, 129.3928, 129.947, 130.4693, 130.8683, 
    131.1357, 131.3994, 132.2002, 132.625, 133.5796, 133.4069, 133.6995, 
    133.9792, 134.4498, 134.3723, 134.5799, 133.6917, 134.2816, 133.3086, 
    133.5743, 131.4716, 130.6756, 130.3386, 130.0437, 129.3285, 129.8222, 
    129.6274, 130.091, 130.3861, 130.2401, 131.143, 130.7915, 132.6502, 
    131.8475, 133.9466, 133.4423, 134.0676, 133.7483, 134.2957, 133.803, 
    134.6572, 134.8438, 134.7163, 135.2062, 133.7757, 134.324, 130.236, 
    130.2598, 130.3707, 129.8836, 129.8538, 129.4083, 129.8046, 129.9736, 
    130.4032, 130.6578, 130.9001, 131.4338, 132.0316, 132.8704, 133.475, 
    133.8813, 133.632, 133.8521, 133.6061, 133.4909, 134.7739, 134.0526, 
    135.1357, 135.0756, 134.5849, 135.0823, 130.2765, 130.1395, 129.6647, 
    130.0362, 129.3598, 129.7382, 129.9561, 130.7989, 130.9845, 131.1568, 
    131.4975, 131.9356, 132.7064, 133.3793, 133.9955, 133.9503, 133.9662, 
    134.1041, 133.7627, 134.1602, 134.227, 134.0524, 135.0675, 134.777, 
    135.0743, 134.8851, 130.184, 130.4146, 130.29, 130.5245, 130.3593, 
    131.0949, 131.316, 132.3535, 131.927, 132.6061, 131.9958, 132.1038, 
    132.6285, 132.0287, 133.3423, 132.451, 134.1095, 133.2164, 134.1656, 
    133.9928, 134.2789, 134.5355, 134.8586, 135.4563, 135.3177, 135.8185, 
    130.7589, 131.0589, 131.0324, 131.3468, 131.5796, 132.0851, 132.8985, 
    132.5922, 133.1547, 133.2679, 132.4133, 132.9377, 131.2599, 131.5302, 
    131.3692, 130.7826, 132.6629, 131.6958, 133.485, 132.9585, 134.4989, 
    133.7315, 135.2415, 135.8906, 136.5028, 137.221, 131.2228, 131.0187, 
    131.3842, 131.8911, 132.3623, 132.9906, 133.0549, 133.1729, 133.4787, 
    133.7361, 133.2103, 133.8007, 131.5931, 132.747, 130.9417, 131.4837, 
    131.8611, 131.6954, 132.5572, 132.7609, 133.5906, 133.1612, 135.7303, 
    134.5898, 137.7691, 136.8759, 130.9475, 131.222, 132.1807, 131.724, 
    133.0325, 133.3559, 133.6191, 133.9562, 133.9926, 134.1925, 133.8649, 
    134.1796, 132.9919, 133.5218, 132.0708, 132.4231, 132.2609, 132.0832, 
    132.6321, 133.2186, 133.231, 133.4194, 133.9516, 133.0378, 135.8782, 
    134.1198, 131.5219, 132.0528, 132.1286, 131.9227, 133.3235, 132.8148, 
    134.1876, 133.8157, 134.4254, 134.1222, 134.0777, 133.689, 133.4474, 
    132.8382, 132.3438, 131.9525, 132.0434, 132.4734, 133.2545, 133.9959, 
    133.8333, 134.379, 132.9374, 133.5408, 133.3074, 133.9164, 132.5841, 
    133.7185, 132.2952, 132.4196, 132.8048, 133.5818, 133.7539, 133.9381, 
    133.8244, 133.2743, 133.1842, 132.7954, 132.6882, 132.3925, 132.148, 
    132.3714, 132.6062, 133.2745, 133.8786, 134.5392, 134.7011, 135.4765, 
    134.8452, 135.8881, 135.0014, 136.5384, 133.7842, 134.9751, 132.8223, 
    133.0531, 133.4714, 134.4337, 133.9135, 134.522, 133.1807, 132.4884, 
    132.3094, 131.9763, 132.3171, 132.2893, 132.6159, 132.5109, 133.2967, 
    132.8742, 134.0766, 134.5171, 135.766, 136.5353, 137.321, 137.6688, 
    137.7748, 137.8191,
  194.4207, 195.5341, 195.3173, 196.2009, 195.7176, 196.2882, 194.646, 
    195.5785, 194.9828, 194.5206, 197.8987, 196.2398, 199.632, 198.5661, 
    201.2515, 199.466, 201.6129, 201.1996, 202.4449, 202.0876, 203.687, 
    202.61, 204.5194, 203.4293, 203.5996, 202.5746, 196.5726, 197.6916, 
    196.5065, 196.6658, 196.5943, 195.7276, 195.2776, 194.3356, 194.5064, 
    195.1983, 196.7374, 196.2197, 197.5261, 197.4965, 198.9584, 198.2983, 
    200.7672, 200.0632, 202.1025, 201.5882, 202.0783, 201.9296, 202.0803, 
    201.3264, 201.6492, 200.9867, 198.4218, 199.1732, 196.9386, 195.6006, 
    194.6868, 194.0404, 194.1317, 194.3058, 195.2024, 196.0364, 196.6608, 
    197.0793, 197.4922, 198.7466, 199.4126, 200.9099, 200.6389, 201.098, 
    201.5371, 202.2761, 202.1543, 202.4804, 201.0858, 202.0119, 200.4847, 
    200.9016, 197.6052, 196.3592, 195.8318, 195.359, 194.2019, 195.0005, 
    194.6854, 195.4354, 195.9062, 195.6768, 197.0907, 196.5405, 199.4521, 
    198.1941, 201.4859, 200.6945, 201.6758, 201.1746, 202.0341, 201.2604, 
    202.6018, 202.8949, 202.6946, 203.4645, 201.2176, 202.0784, 195.6702, 
    195.7086, 195.8822, 195.0998, 195.0516, 194.331, 194.972, 195.2455, 
    195.933, 196.3313, 196.7105, 197.5461, 198.4826, 199.7973, 200.7457, 
    201.3833, 200.9922, 201.3375, 200.9515, 200.7707, 202.7851, 201.6522, 
    203.3536, 203.2592, 202.4882, 203.2698, 195.7348, 195.514, 194.7457, 
    195.3468, 194.2526, 194.8646, 195.2172, 196.5521, 196.8426, 197.1123, 
    197.6458, 198.332, 199.5401, 200.5956, 201.5626, 201.4917, 201.5166, 
    201.7332, 201.1972, 201.8213, 201.9262, 201.652, 203.2465, 202.79, 
    203.2572, 202.9598, 195.5861, 195.9509, 195.7559, 196.1227, 195.8643, 
    197.0155, 197.3616, 198.9869, 198.3185, 199.3829, 198.4264, 198.5957, 
    199.418, 198.478, 200.5374, 199.1397, 201.7416, 200.3399, 201.8297, 
    201.5585, 202.0076, 202.4106, 202.9182, 203.8576, 203.6398, 204.4271, 
    196.4895, 196.9591, 196.9176, 197.4099, 197.7745, 198.5663, 199.8414, 
    199.3612, 200.2433, 200.4208, 199.0808, 199.9028, 197.2738, 197.697, 
    197.4449, 196.5266, 199.4719, 197.9564, 200.7614, 199.9355, 202.3531, 
    201.1482, 203.52, 204.5405, 205.5038, 206.6344, 197.2157, 196.8962, 
    197.4684, 198.2623, 199.0008, 199.9858, 200.0867, 200.2717, 200.7515, 
    201.1555, 200.3304, 201.2569, 197.7954, 199.6038, 196.7756, 197.6243, 
    198.2154, 197.9558, 199.3063, 199.6256, 200.9271, 200.2535, 204.2883, 
    202.4959, 207.4979, 206.0911, 196.7847, 197.2145, 198.7161, 198.0006, 
    200.0516, 200.5589, 200.9719, 201.5009, 201.558, 201.872, 201.3577, 
    201.8516, 199.9879, 200.8192, 198.5439, 199.096, 198.8418, 198.5634, 
    199.4237, 200.3434, 200.3629, 200.6585, 201.4936, 200.06, 204.5209, 
    201.7577, 197.684, 198.5157, 198.6344, 198.3119, 200.508, 199.7102, 
    201.8643, 201.2804, 202.2377, 201.7616, 201.6917, 201.0815, 200.7024, 
    199.7468, 198.9717, 198.3586, 198.501, 199.175, 200.3997, 201.5633, 
    201.308, 202.1649, 199.9024, 200.8489, 200.4827, 201.4385, 199.3484, 
    201.1278, 198.8956, 199.0905, 199.6944, 200.9133, 201.1835, 201.4725, 
    201.2941, 200.4308, 200.2896, 199.6797, 199.5116, 199.048, 198.6649, 
    199.015, 199.3831, 200.4311, 201.3791, 202.4164, 202.6707, 203.8892, 
    202.8971, 204.5364, 203.1425, 205.5596, 201.231, 203.1012, 199.7219, 
    200.0839, 200.7401, 202.2508, 201.434, 202.3893, 200.284, 199.1983, 
    198.9179, 198.3959, 198.9299, 198.8864, 199.3983, 199.2337, 200.466, 
    199.8033, 201.69, 202.3817, 204.3446, 205.5549, 206.792, 207.34, 207.507, 
    207.5768,
  318.5596, 320.359, 320.0084, 321.4653, 320.6563, 321.6114, 318.9236, 
    320.4308, 319.4678, 318.7211, 324.3105, 321.5304, 327.1914, 325.4309, 
    329.8244, 326.9217, 330.4126, 329.7401, 331.7679, 331.1857, 333.7932, 
    332.037, 335.1525, 333.3729, 333.6507, 331.9792, 322.0879, 323.9633, 
    321.9771, 322.2439, 322.1241, 320.6731, 319.9443, 318.4223, 318.6981, 
    319.8161, 322.3638, 321.4967, 323.6858, 323.6362, 326.0896, 324.9813, 
    329.0365, 327.8919, 331.21, 330.3725, 331.1706, 330.9284, 331.1738, 
    329.9464, 330.4717, 329.3936, 325.1886, 326.4462, 322.701, 320.4664, 
    318.9896, 317.9456, 318.093, 318.3742, 319.8226, 321.1898, 322.2355, 
    322.9368, 323.6291, 325.7338, 326.8349, 329.2686, 328.8279, 329.5746, 
    330.2893, 331.4928, 331.2944, 331.8257, 329.5547, 331.0624, 328.5771, 
    329.2551, 323.8183, 321.7304, 320.8474, 320.0758, 318.2064, 319.4963, 
    318.9873, 320.1995, 320.972, 320.5897, 322.956, 322.0341, 326.8991, 
    324.8064, 330.2058, 328.9183, 330.5152, 329.6993, 331.0985, 329.839, 
    332.0236, 332.5013, 332.1748, 333.4303, 329.7693, 331.1707, 320.579, 
    320.6413, 320.9318, 319.6569, 319.579, 318.4148, 319.4504, 319.8925, 
    321.0168, 321.6837, 322.3189, 323.7195, 325.2905, 327.4599, 329.0016, 
    330.039, 329.4025, 329.9644, 329.3363, 329.0423, 332.3222, 330.4767, 
    333.2495, 333.0954, 331.8384, 333.1128, 320.6851, 320.3265, 319.0847, 
    320.0562, 318.2883, 319.2768, 319.8466, 322.0535, 322.5401, 322.9922, 
    323.8866, 325.0379, 327.0422, 328.7575, 330.3309, 330.2153, 330.256, 
    330.6085, 329.7361, 330.7519, 330.9228, 330.4763, 333.0748, 332.3304, 
    333.0921, 332.6072, 320.443, 321.0468, 320.7204, 321.3344, 320.9018, 
    322.8298, 323.4099, 326.1374, 325.0153, 326.7868, 325.1964, 325.4805, 
    326.8436, 325.2829, 328.6628, 326.3919, 330.6222, 328.3416, 330.7657, 
    330.324, 331.0554, 331.7119, 332.5394, 334.0719, 333.7164, 335.0018, 
    321.9487, 322.7354, 322.666, 323.491, 324.1024, 325.4312, 327.5315, 
    326.7516, 328.1847, 328.4732, 326.2952, 327.6313, 323.2629, 323.9723, 
    323.5496, 322.0107, 326.9313, 324.4075, 329.0272, 327.6844, 331.6182, 
    329.6563, 333.5209, 335.1869, 336.7615, 338.6118, 323.1654, 322.63, 
    323.5891, 324.9209, 326.1607, 327.7661, 327.9302, 328.2309, 329.011, 
    329.6683, 328.3262, 329.8333, 324.1374, 327.1456, 322.4279, 323.8504, 
    324.8422, 324.4066, 326.6625, 327.1811, 329.2967, 328.2013, 334.7751, 
    331.8509, 340.0269, 337.7224, 322.4431, 323.1635, 325.6826, 324.4817, 
    327.8731, 328.6978, 329.3695, 330.2304, 330.3233, 330.8346, 329.9973, 
    330.8014, 327.7696, 329.1211, 325.3936, 326.3207, 325.8938, 325.4263, 
    326.8531, 328.3473, 328.3791, 328.8597, 330.2182, 327.8867, 335.1547, 
    330.6482, 323.9507, 325.346, 325.5455, 325.0041, 328.615, 327.3185, 
    330.8221, 329.8715, 331.4303, 330.6548, 330.5409, 329.5478, 328.9311, 
    327.3778, 326.1119, 325.0826, 325.3216, 326.4492, 328.4389, 330.3319, 
    329.9163, 331.3116, 327.6306, 329.1694, 328.5739, 330.1287, 326.7309, 
    329.6229, 325.9841, 326.3115, 327.2928, 329.2741, 329.7137, 330.1841, 
    329.8937, 328.4895, 328.2599, 327.2689, 326.9958, 326.2402, 325.5968, 
    326.1847, 326.7872, 328.49, 330.0321, 331.7213, 332.1359, 334.1233, 
    332.5049, 335.1801, 332.9048, 336.8528, 329.7909, 332.8377, 327.3374, 
    327.9256, 328.9924, 331.4514, 330.1214, 331.6772, 328.2509, 326.4871, 
    326.0216, 325.1451, 326.0417, 325.9686, 326.8118, 326.5445, 328.5467, 
    327.4697, 330.5381, 331.6649, 334.8669, 336.845, 338.87, 339.768, 
    340.0417, 340.1562,
  524.3479, 527.6205, 526.9822, 529.6362, 528.1619, 529.9026, 525.0092, 
    527.751, 525.9987, 524.6413, 534.8335, 529.7549, 540.1708, 536.8854, 
    545.1854, 539.6581, 546.3083, 545.0246, 548.8989, 547.7855, 552.7794, 
    549.4138, 555.39, 551.9731, 552.506, 549.3032, 530.7719, 534.1981, 
    530.5698, 531.0565, 530.838, 528.1924, 526.8655, 524.0986, 524.5995, 
    526.6322, 531.2755, 529.6935, 533.6908, 533.6002, 538.0932, 536.0616, 
    543.6831, 541.5033, 547.8319, 546.2318, 547.7567, 547.2936, 547.7627, 
    545.4183, 546.4212, 544.3638, 536.4415, 538.755, 531.8911, 527.8159, 
    525.1292, 523.2268, 523.5005, 524.0112, 526.6442, 529.134, 531.0413, 
    532.3218, 533.5871, 537.4407, 539.4933, 544.1254, 543.2855, 544.709, 
    546.0729, 548.3726, 547.9932, 549.0095, 544.6712, 547.5497, 542.8079, 
    544.0998, 533.933, 530.1197, 528.5099, 527.1049, 523.7064, 526.0505, 
    525.125, 527.33, 528.7371, 528.0405, 532.3568, 530.6737, 539.6154, 
    535.7413, 545.9136, 543.4578, 546.5042, 544.947, 547.6187, 545.2134, 
    549.3882, 550.3027, 549.6776, 552.0833, 545.0805, 547.7568, 528.0211, 
    528.1346, 528.6638, 526.3425, 526.2009, 524.0849, 525.9671, 526.7712, 
    528.8187, 530.0345, 531.1934, 533.7523, 536.6282, 540.6814, 543.6165, 
    545.5952, 544.3807, 545.4528, 544.2546, 543.6941, 549.9599, 546.4307, 
    551.7365, 551.4412, 549.0337, 551.4744, 528.2143, 527.5613, 525.3022, 
    527.0692, 523.855, 525.6514, 526.6877, 530.7091, 531.5974, 532.423, 
    534.058, 536.1654, 539.8872, 543.1513, 546.1523, 545.9317, 546.0093, 
    546.6825, 545.0172, 546.9565, 547.2829, 546.4301, 551.4016, 549.9755, 
    551.4349, 550.5057, 527.7734, 528.8732, 528.2786, 529.3975, 528.609, 
    532.1262, 533.1863, 538.1809, 536.1239, 539.4019, 536.4556, 536.9763, 
    539.5098, 536.6143, 542.9709, 538.6517, 546.7087, 542.3591, 546.9827, 
    546.1393, 547.5364, 548.7917, 550.3759, 553.3142, 552.632, 555.1005, 
    530.5178, 531.954, 531.8271, 533.3345, 534.4528, 536.8861, 540.8177, 
    539.335, 542.0605, 542.6099, 538.4704, 541.0076, 532.9176, 534.2147, 
    533.4418, 530.631, 539.6765, 535.011, 543.6653, 541.1085, 548.6126, 
    544.8648, 552.257, 555.4561, 558.4692, 561.9199, 532.7395, 531.7614, 
    533.514, 535.951, 538.2238, 541.264, 541.5761, 542.1486, 543.6344, 
    544.8878, 542.3299, 545.2025, 534.5166, 540.0837, 531.3924, 533.9917, 
    535.8069, 535.0095, 539.1658, 540.1512, 544.179, 542.0921, 554.6646, 
    549.0577, 564.5654, 560.2599, 531.4202, 532.736, 537.3469, 535.1469, 
    541.4676, 543.0377, 544.3179, 545.9604, 546.1379, 547.1144, 545.5154, 
    547.051, 541.2705, 543.8442, 536.8171, 538.5172, 537.7342, 536.8771, 
    539.5278, 542.3701, 542.4307, 543.3462, 545.937, 541.4933, 555.3942, 
    546.7582, 534.1754, 536.7299, 537.0956, 536.1035, 542.88, 540.4125, 
    547.0905, 545.2755, 548.2532, 546.771, 546.5534, 544.658, 543.4822, 
    540.5254, 538.1343, 536.2472, 536.6852, 538.7606, 542.5445, 546.1542, 
    545.361, 548.0261, 541.0062, 543.9363, 542.8016, 545.7664, 539.2957, 
    544.801, 537.8998, 538.5004, 540.3636, 544.136, 544.9744, 545.8721, 
    545.3179, 542.6409, 542.2037, 540.3182, 539.7992, 538.3696, 537.1896, 
    538.2676, 539.4027, 542.6418, 545.5818, 548.8097, 549.6031, 553.4128, 
    550.3096, 555.4429, 551.0756, 558.6389, 545.1215, 550.947, 540.4485, 
    541.5674, 543.5989, 548.2935, 545.7524, 548.7254, 542.1866, 538.8326, 
    537.9686, 536.3618, 538.0054, 537.8714, 539.4495, 538.9418, 542.7498, 
    540.7001, 546.548, 548.7018, 554.8412, 558.6246, 562.4023, 564.081, 
    564.5932, 564.8076,
  947.2584, 954.1312, 952.7881, 958.382, 955.2715, 958.9449, 948.6445, 
    954.4061, 950.7208, 947.8732, 969.2601, 958.6328, 980.2999, 973.493, 
    990.7613, 979.2354, 993.116, 990.4244, 998.5654, 996.2203, 1006.774, 
    999.6513, 1012.327, 1005.064, 1006.194, 999.4181, 960.7829, 967.9522, 
    960.3553, 961.3853, 960.9227, 955.3359, 952.5425, 946.7362, 947.7856, 
    952.0521, 961.849, 958.5031, 966.9091, 966.7227, 975.9911, 971.792, 
    987.618, 983.0713, 996.3179, 992.9552, 996.1596, 995.1858, 996.1723, 
    991.2491, 993.3529, 989.0411, 972.576, 977.3621, 963.1533, 954.5427, 
    948.896, 944.9249, 945.4846, 946.5532, 952.0771, 957.3218, 961.3531, 
    964.0666, 966.6959, 974.6409, 978.8933, 988.5426, 986.7875, 989.7637, 
    992.6218, 997.4564, 996.6575, 998.7985, 989.6844, 995.7244, 985.7905, 
    988.489, 967.4069, 959.4036, 956.0052, 953.0461, 945.9153, 950.8298, 
    948.8872, 953.5197, 956.4843, 955.0159, 964.141, 960.5753, 979.1465, 
    971.1312, 992.2877, 987.1472, 993.5272, 990.2618, 995.8694, 990.8199, 
    999.5974, 1001.528, 1000.208, 1005.297, 990.5415, 996.1599, 954.9749, 
    955.2141, 956.3297, 951.4432, 951.1456, 946.7076, 950.6545, 952.3442, 
    956.6564, 959.2236, 961.6752, 967.0355, 972.9617, 981.3611, 987.4789, 
    991.6199, 989.0767, 991.3214, 988.8128, 987.641, 1000.804, 993.3727, 
    1004.562, 1003.937, 998.8496, 1004.007, 955.3821, 954.0067, 949.259, 
    952.9709, 946.2264, 949.9917, 952.1687, 960.6501, 962.5308, 964.2813, 
    967.664, 972.0061, 979.7109, 986.5073, 992.7885, 992.3257, 992.4886, 
    993.9015, 990.4089, 994.4771, 995.1632, 993.3715, 1003.853, 1000.837, 
    1003.923, 1001.958, 954.4534, 956.7715, 955.5176, 957.8779, 956.2142, 
    963.6519, 965.8724, 976.1727, 971.9205, 978.7036, 972.6053, 973.6809, 
    978.9274, 972.9329, 986.1307, 977.1479, 993.9565, 984.8542, 994.5322, 
    992.7612, 995.6964, 998.3395, 1001.683, 1007.909, 1006.461, 1011.71, 
    960.2455, 963.2866, 963.0177, 966.1769, 968.4763, 973.4944, 981.6445, 
    978.5648, 984.232, 985.3773, 976.7724, 982.0394, 965.3206, 967.9865, 
    966.3973, 960.485, 979.2735, 969.6259, 987.5807, 982.2493, 997.9619, 
    990.0898, 1005.665, 1012.468, 1018.949, 1026.627, 964.953, 962.8785, 
    966.5458, 971.5637, 976.2614, 982.5731, 983.2229, 984.4153, 987.5162, 
    990.1378, 984.7935, 990.797, 968.6077, 980.1191, 962.0967, 967.5277, 
    971.2664, 969.6226, 978.2138, 980.2593, 988.6546, 984.2978, 1010.781, 
    998.9001, 1032.433, 1022.927, 962.1557, 964.9456, 974.4469, 969.9058, 
    982.9969, 986.2699, 988.9453, 992.3859, 992.7584, 994.8089, 991.4529, 
    994.6758, 982.5866, 987.9547, 973.3519, 976.8693, 975.2481, 973.4758, 
    978.9649, 984.8773, 985.0035, 986.9141, 992.3367, 983.0505, 1012.336, 
    994.0604, 967.9055, 973.1718, 973.9274, 971.8784, 985.9409, 980.8022, 
    994.7587, 990.9501, 997.2047, 994.0875, 993.6304, 989.6568, 987.1981, 
    981.0369, 976.0761, 972.1749, 973.0794, 977.3737, 985.2409, 992.7924, 
    991.1291, 996.7267, 982.0367, 988.1472, 985.7773, 991.979, 978.4833, 
    989.9561, 975.5907, 976.8345, 980.7007, 988.5648, 990.3194, 992.2008, 
    991.0389, 985.442, 984.5304, 980.6062, 979.5282, 976.5634, 974.1218, 
    976.3524, 978.7052, 985.444, 991.592, 998.3773, 1000.051, 1008.119, 
    1001.543, 1012.44, 1003.163, 1019.325, 990.6274, 1002.891, 980.877, 
    983.2048, 987.4421, 997.2896, 991.9496, 998.1997, 984.4946, 977.5229, 
    975.7331, 972.4114, 975.8093, 975.532, 978.8024, 977.7492, 985.6693, 
    981.4001, 993.6192, 998.1498, 1011.158, 1019.293, 1027.704, 1031.382, 
    1032.494, 1032.959,
  1829.891, 1849.353, 1845.525, 1861.55, 1852.613, 1863.175, 1833.791, 
    1850.138, 1839.657, 1831.62, 1893.772, 1862.273, 1928.095, 1906.814, 
    1960.691, 1924.741, 1968.121, 1959.632, 1985.507, 1977.992, 2012.212, 
    1989.003, 2030.648, 2006.596, 2010.304, 1988.252, 1868.494, 1889.771, 
    1867.255, 1870.243, 1868.9, 1852.797, 1844.827, 1828.425, 1831.373, 
    1843.433, 1871.591, 1861.899, 1886.589, 1886.022, 1914.579, 1901.556, 
    1950.848, 1936.759, 1978.304, 1967.612, 1977.798, 1974.693, 1977.839, 
    1962.226, 1968.871, 1955.293, 1903.977, 1918.863, 1875.39, 1850.529, 
    1834.5, 1823.354, 1824.919, 1827.912, 1843.504, 1858.497, 1870.15, 
    1878.058, 1885.94, 1910.376, 1923.666, 1953.734, 1948.261, 1957.557, 
    1966.558, 1981.947, 1979.389, 1986.256, 1957.309, 1976.409, 1945.164, 
    1953.567, 1888.107, 1864.5, 1854.715, 1846.26, 1826.124, 1839.966, 
    1834.475, 1847.609, 1856.09, 1851.882, 1878.275, 1867.892, 1924.461, 
    1899.519, 1965.502, 1949.38, 1969.423, 1959.121, 1976.872, 1960.875, 
    1988.829, 1995.074, 1990.801, 2007.361, 1960, 1977.799, 1851.764, 
    1852.449, 1855.646, 1841.704, 1840.86, 1828.345, 1839.469, 1844.263, 
    1856.584, 1863.98, 1871.086, 1886.974, 1905.169, 1931.447, 1950.414, 
    1963.395, 1955.405, 1962.454, 1954.579, 1950.919, 1992.728, 1968.934, 
    2004.954, 2002.91, 1986.421, 2003.14, 1852.93, 1848.998, 1835.524, 
    1846.046, 1826.996, 1837.594, 1843.764, 1868.109, 1873.575, 1878.686, 
    1888.891, 1902.216, 1926.238, 1947.389, 1967.085, 1965.622, 1966.136, 
    1970.611, 1959.583, 1972.438, 1974.621, 1968.93, 2002.637, 1992.835, 
    2002.867, 1996.466, 1850.273, 1856.914, 1853.318, 1860.097, 1855.315, 
    1876.846, 1883.436, 1915.146, 1901.952, 1923.069, 1904.067, 1907.396, 
    1923.773, 1905.08, 1946.22, 1918.193, 1970.785, 1942.263, 1972.614, 
    1966.998, 1976.32, 1984.781, 1995.575, 2015.958, 2011.183, 2028.584, 
    1866.936, 1875.779, 1874.995, 1884.361, 1891.372, 1906.819, 1932.344, 
    1922.633, 1940.339, 1943.882, 1917.018, 1933.586, 1881.761, 1889.876, 
    1885.031, 1867.631, 1924.861, 1894.893, 1950.731, 1934.231, 1983.568, 
    1958.581, 2008.569, 2031.119, 2053.034, 2079.24, 1880.652, 1874.589, 
    1885.483, 1900.852, 1915.423, 1935.226, 1937.226, 1940.906, 1950.53, 
    1958.732, 1942.075, 1960.803, 1891.774, 1927.524, 1872.311, 1888.475, 
    1899.936, 1894.883, 1921.532, 1927.967, 1954.084, 1940.542, 2025.485, 
    1986.584, 2099.509, 2066.705, 1872.483, 1880.631, 1909.773, 1895.752, 
    1936.53, 1946.652, 1954.993, 1965.812, 1966.989, 1973.493, 1962.868, 
    1973.07, 1935.267, 1951.898, 1906.377, 1917.321, 1912.264, 1906.761, 
    1923.891, 1942.334, 1942.725, 1948.655, 1965.657, 1936.695, 2030.677, 
    1971.115, 1889.628, 1905.819, 1908.161, 1901.822, 1945.63, 1929.68, 
    1973.334, 1961.285, 1981.141, 1971.201, 1969.751, 1957.222, 1949.539, 
    1930.422, 1914.845, 1902.738, 1905.534, 1918.899, 1943.46, 1967.097, 
    1961.848, 1979.611, 1933.577, 1952.499, 1945.123, 1964.527, 1922.378, 
    1958.161, 1913.331, 1917.213, 1929.359, 1953.803, 1959.302, 1965.227, 
    1961.564, 1944.083, 1941.261, 1929.061, 1925.662, 1916.366, 1908.764, 
    1915.707, 1923.074, 1944.089, 1963.307, 1984.902, 1990.293, 2016.649, 
    1995.121, 2031.025, 2000.386, 2054.321, 1960.27, 1999.5, 1929.917, 
    1937.17, 1950.299, 1981.412, 1964.434, 1984.332, 1941.151, 1919.366, 
    1913.775, 1903.468, 1914.012, 1913.149, 1923.38, 1920.075, 1944.788, 
    1931.57, 1969.715, 1984.171, 2026.74, 2054.213, 2082.9, 2095.761, 
    2099.724, 2101.388,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.536768, 4.555262, 4.551662, 4.566609, 4.558312, 4.568107, 4.540512, 
    4.555998, 4.546107, 4.53843, 4.595716, 4.567276, 4.625376, 4.607146, 
    4.65303, 4.622537, 4.659195, 4.652147, 4.673377, 4.667288, 4.694517, 
    4.676189, 4.70867, 4.690135, 4.693032, 4.675585, 4.572988, 4.592169, 
    4.571854, 4.574585, 4.573359, 4.558485, 4.551003, 4.535356, 4.538193, 
    4.549686, 4.575813, 4.566931, 4.589335, 4.588828, 4.613858, 4.602561, 
    4.644767, 4.632744, 4.667542, 4.658775, 4.66713, 4.664596, 4.667163, 
    4.65431, 4.659814, 4.648513, 4.604676, 4.617531, 4.579264, 4.556363, 
    4.541191, 4.530447, 4.531965, 4.53486, 4.549754, 4.563786, 4.5745, 
    4.581676, 4.588755, 4.610233, 4.621624, 4.647202, 4.642577, 4.650412, 
    4.657903, 4.6705, 4.668425, 4.673981, 4.650204, 4.665998, 4.639945, 
    4.647061, 4.590688, 4.569326, 4.560273, 4.552354, 4.533133, 4.546401, 
    4.541167, 4.553624, 4.561552, 4.557629, 4.581873, 4.572437, 4.6223, 
    4.600777, 4.657029, 4.643526, 4.660269, 4.65172, 4.666376, 4.653184, 
    4.676049, 4.681039, 4.677629, 4.690734, 4.652454, 4.667131, 4.557519, 
    4.558159, 4.561139, 4.54805, 4.54725, 4.535278, 4.545929, 4.55047, 
    4.562011, 4.568848, 4.575353, 4.589678, 4.605715, 4.628201, 4.644401, 
    4.655281, 4.648607, 4.654499, 4.647913, 4.644828, 4.679169, 4.659866, 
    4.688848, 4.687241, 4.674113, 4.687422, 4.558608, 4.554928, 4.54217, 
    4.552152, 4.533976, 4.544145, 4.549999, 4.572636, 4.577618, 4.582243, 
    4.591386, 4.603139, 4.623806, 4.641838, 4.658339, 4.657128, 4.657555, 
    4.661246, 4.652106, 4.662748, 4.664536, 4.659863, 4.687026, 4.679255, 
    4.687206, 4.682146, 4.556124, 4.562318, 4.55897, 4.565267, 4.560831, 
    4.580582, 4.586514, 4.614345, 4.602908, 4.621117, 4.604754, 4.607651, 
    4.621715, 4.605637, 4.640843, 4.616958, 4.66139, 4.637469, 4.662892, 
    4.658267, 4.665925, 4.672791, 4.681437, 4.697421, 4.693717, 4.707103, 
    4.571562, 4.579617, 4.578906, 4.587343, 4.59359, 4.60715, 4.628954, 
    4.620746, 4.635821, 4.638853, 4.615952, 4.630004, 4.585011, 4.592262, 
    4.587943, 4.572198, 4.622639, 4.596706, 4.644669, 4.630562, 4.671812, 
    4.651268, 4.691678, 4.709027, 4.725387, 4.74456, 4.584015, 4.578537, 
    4.588347, 4.601945, 4.614583, 4.631422, 4.633147, 4.636307, 4.644499, 
    4.651395, 4.637308, 4.653124, 4.593947, 4.624894, 4.576469, 4.591016, 
    4.601142, 4.596697, 4.619809, 4.625268, 4.647497, 4.635996, 4.704742, 
    4.674244, 4.759188, 4.735351, 4.576625, 4.583995, 4.609712, 4.597464, 
    4.632547, 4.641211, 4.648261, 4.657286, 4.65826, 4.663613, 4.654843, 
    4.663266, 4.631458, 4.645654, 4.606766, 4.616211, 4.611864, 4.6071, 
    4.621815, 4.63753, 4.637864, 4.642911, 4.657158, 4.632689, 4.708693, 
    4.661662, 4.592041, 4.606281, 4.608315, 4.602794, 4.640342, 4.626713, 
    4.663483, 4.653525, 4.669847, 4.661732, 4.660539, 4.650131, 4.643661, 
    4.627338, 4.614086, 4.603594, 4.606032, 4.617562, 4.638492, 4.65835, 
    4.653995, 4.668605, 4.629997, 4.646161, 4.63991, 4.656221, 4.620529, 
    4.650918, 4.612783, 4.616118, 4.626443, 4.64726, 4.651871, 4.656802, 
    4.653759, 4.639024, 4.636611, 4.626192, 4.623318, 4.615392, 4.608837, 
    4.614826, 4.621121, 4.639029, 4.655208, 4.672889, 4.677222, 4.697956, 
    4.681077, 4.708956, 4.685251, 4.726333, 4.652679, 4.68455, 4.626913, 
    4.633099, 4.644304, 4.670067, 4.656144, 4.672429, 4.636517, 4.617961, 
    4.613165, 4.604232, 4.61337, 4.612626, 4.621381, 4.618566, 4.639624, 
    4.628304, 4.66051, 4.672299, 4.705699, 4.726254, 4.747232, 4.756515, 
    4.759342, 4.760524,
  5.626039, 5.649297, 5.644769, 5.66357, 5.653134, 5.665454, 5.630748, 
    5.650223, 5.637784, 5.628129, 5.700191, 5.66441, 5.737524, 5.714577, 
    5.772345, 5.73395, 5.780109, 5.771232, 5.797972, 5.790303, 5.824607, 
    5.801515, 5.842442, 5.819085, 5.822735, 5.800755, 5.671595, 5.695728, 
    5.670168, 5.673604, 5.672061, 5.653351, 5.64394, 5.624263, 5.627831, 
    5.642285, 5.675149, 5.663976, 5.692163, 5.691525, 5.723025, 5.708807, 
    5.761939, 5.746801, 5.790622, 5.77958, 5.790104, 5.786911, 5.790145, 
    5.773956, 5.780889, 5.766656, 5.711468, 5.727648, 5.679491, 5.650682, 
    5.631601, 5.618092, 5.62, 5.62364, 5.642369, 5.660018, 5.673497, 
    5.682526, 5.691433, 5.718462, 5.732801, 5.765005, 5.759181, 5.769048, 
    5.778482, 5.794349, 5.791735, 5.798733, 5.768785, 5.788677, 5.755867, 
    5.764827, 5.693865, 5.666988, 5.6556, 5.64564, 5.621468, 5.638153, 
    5.631571, 5.647237, 5.657208, 5.652275, 5.682773, 5.670902, 5.733652, 
    5.706561, 5.777381, 5.760376, 5.781462, 5.770695, 5.789153, 5.772539, 
    5.801339, 5.807625, 5.803329, 5.81984, 5.771619, 5.790105, 5.652137, 
    5.652941, 5.65669, 5.640227, 5.639221, 5.624166, 5.637559, 5.643271, 
    5.657786, 5.666387, 5.674571, 5.692595, 5.712776, 5.741081, 5.761477, 
    5.775179, 5.766774, 5.774194, 5.7659, 5.762015, 5.805269, 5.780953, 
    5.817463, 5.815438, 5.7989, 5.815666, 5.653506, 5.648878, 5.632832, 
    5.645386, 5.622528, 5.635315, 5.642679, 5.671152, 5.67742, 5.683239, 
    5.694743, 5.709534, 5.735547, 5.75825, 5.77903, 5.777506, 5.778043, 
    5.782693, 5.771181, 5.784584, 5.786837, 5.78095, 5.815167, 5.805377, 
    5.815395, 5.809019, 5.650382, 5.658173, 5.653962, 5.661882, 5.656302, 
    5.681149, 5.688613, 5.723638, 5.709242, 5.732163, 5.711567, 5.715213, 
    5.732915, 5.712678, 5.756999, 5.726927, 5.782874, 5.752749, 5.784765, 
    5.778941, 5.788586, 5.797235, 5.808127, 5.828266, 5.823598, 5.840467, 
    5.669801, 5.679934, 5.67904, 5.689656, 5.697517, 5.714581, 5.742029, 
    5.731696, 5.750675, 5.754491, 5.72566, 5.743351, 5.686722, 5.695845, 
    5.690411, 5.670601, 5.734078, 5.701437, 5.761815, 5.744053, 5.796001, 
    5.770126, 5.82103, 5.842893, 5.863514, 5.887687, 5.685468, 5.678577, 
    5.690919, 5.708031, 5.723937, 5.745136, 5.747307, 5.751287, 5.761601, 
    5.770285, 5.752547, 5.772463, 5.697966, 5.736917, 5.675974, 5.694278, 
    5.70702, 5.701427, 5.730515, 5.737388, 5.765376, 5.750895, 5.837492, 
    5.799065, 5.906134, 5.876075, 5.676171, 5.685444, 5.717806, 5.702391, 
    5.746552, 5.757461, 5.766339, 5.777705, 5.778931, 5.785674, 5.774628, 
    5.785236, 5.745181, 5.763056, 5.714098, 5.725987, 5.720515, 5.714518, 
    5.733041, 5.752826, 5.753247, 5.759602, 5.777543, 5.746732, 5.842471, 
    5.783216, 5.695569, 5.713488, 5.716048, 5.709099, 5.756367, 5.739208, 
    5.785509, 5.772968, 5.793526, 5.783304, 5.781801, 5.768694, 5.760545, 
    5.739994, 5.723311, 5.710106, 5.713175, 5.727687, 5.754037, 5.779044, 
    5.77356, 5.791961, 5.743342, 5.763694, 5.755823, 5.776363, 5.731422, 
    5.769684, 5.721673, 5.72587, 5.738868, 5.765079, 5.770885, 5.777094, 
    5.773262, 5.754707, 5.75167, 5.738551, 5.734934, 5.724956, 5.716706, 
    5.724244, 5.732168, 5.754714, 5.775087, 5.797358, 5.802817, 5.82894, 
    5.807672, 5.842803, 5.812931, 5.864706, 5.771903, 5.812049, 5.739459, 
    5.747247, 5.761355, 5.793803, 5.776267, 5.796778, 5.751551, 5.72819, 
    5.722154, 5.710909, 5.722411, 5.721475, 5.732495, 5.728951, 5.755463, 
    5.741211, 5.781765, 5.796615, 5.838698, 5.864606, 5.891056, 5.902761, 
    5.906327, 5.907819,
  8.094118, 8.128306, 8.12165, 8.149295, 8.133948, 8.152065, 8.101038, 
    8.129667, 8.111381, 8.097189, 8.203166, 8.150529, 8.258118, 8.224336, 
    8.309403, 8.252855, 8.320842, 8.307764, 8.347167, 8.335863, 8.386434, 
    8.352388, 8.412737, 8.37829, 8.383674, 8.351268, 8.161097, 8.196599, 
    8.158998, 8.164051, 8.161782, 8.134267, 8.120432, 8.091507, 8.096751, 
    8.117997, 8.166325, 8.149891, 8.191352, 8.190413, 8.236772, 8.215843, 
    8.294074, 8.271778, 8.336335, 8.320062, 8.33557, 8.330865, 8.335631, 
    8.311776, 8.321991, 8.301023, 8.21976, 8.243577, 8.17271, 8.130343, 
    8.102293, 8.082438, 8.085243, 8.090592, 8.118122, 8.144072, 8.163894, 
    8.177176, 8.190279, 8.230056, 8.251163, 8.29859, 8.290011, 8.304545, 
    8.318444, 8.341826, 8.337974, 8.348289, 8.304159, 8.333468, 8.285129, 
    8.298328, 8.193857, 8.154321, 8.137574, 8.12293, 8.0874, 8.111923, 
    8.102249, 8.125278, 8.139939, 8.132685, 8.177539, 8.160077, 8.252416, 
    8.212539, 8.316822, 8.291771, 8.322835, 8.306972, 8.334169, 8.309689, 
    8.352129, 8.361395, 8.355062, 8.379404, 8.308333, 8.335571, 8.132482, 
    8.133665, 8.139176, 8.114973, 8.113493, 8.091364, 8.111052, 8.119448, 
    8.140789, 8.153437, 8.165473, 8.191988, 8.221685, 8.263354, 8.293393, 
    8.313579, 8.301196, 8.312127, 8.299909, 8.294186, 8.357923, 8.322086, 
    8.375899, 8.372914, 8.348535, 8.373251, 8.134496, 8.12769, 8.104102, 
    8.122557, 8.088957, 8.107752, 8.118576, 8.160445, 8.169664, 8.178225, 
    8.195149, 8.216914, 8.255207, 8.28864, 8.319253, 8.317007, 8.317798, 
    8.324649, 8.307688, 8.327436, 8.330756, 8.322081, 8.372515, 8.358081, 
    8.37285, 8.36345, 8.129901, 8.141356, 8.135165, 8.146812, 8.138606, 
    8.175149, 8.186131, 8.237674, 8.216486, 8.250224, 8.219907, 8.225273, 
    8.251332, 8.221541, 8.286797, 8.242516, 8.324916, 8.280539, 8.327703, 
    8.31912, 8.333333, 8.34608, 8.362136, 8.391829, 8.384945, 8.409823, 
    8.158458, 8.173363, 8.172048, 8.187665, 8.199231, 8.224343, 8.264751, 
    8.249537, 8.277483, 8.283104, 8.240651, 8.266698, 8.183348, 8.196771, 
    8.188775, 8.159635, 8.253044, 8.205, 8.293891, 8.267732, 8.344262, 
    8.306134, 8.381158, 8.413401, 8.443824, 8.479502, 8.181503, 8.171366, 
    8.189523, 8.214703, 8.238114, 8.269326, 8.272523, 8.278383, 8.293576, 
    8.306368, 8.28024, 8.309577, 8.199891, 8.257224, 8.167538, 8.194465, 
    8.213216, 8.204983, 8.247799, 8.257916, 8.299136, 8.277806, 8.405437, 
    8.348778, 8.506738, 8.46236, 8.167827, 8.181468, 8.22909, 8.206403, 
    8.271412, 8.287477, 8.300555, 8.3173, 8.319107, 8.329042, 8.312767, 
    8.328398, 8.269392, 8.295719, 8.223632, 8.241133, 8.233077, 8.22425, 
    8.251517, 8.280651, 8.281271, 8.290631, 8.317061, 8.271676, 8.412779, 
    8.325419, 8.196363, 8.222733, 8.226501, 8.216275, 8.285866, 8.260596, 
    8.328799, 8.310322, 8.340613, 8.32555, 8.323336, 8.304025, 8.292021, 
    8.261755, 8.237193, 8.217757, 8.222273, 8.243635, 8.282435, 8.319272, 
    8.311193, 8.338308, 8.266685, 8.296659, 8.285065, 8.315323, 8.249133, 
    8.305483, 8.234781, 8.240959, 8.260096, 8.298698, 8.307252, 8.316401, 
    8.310754, 8.283422, 8.278949, 8.259629, 8.254304, 8.239614, 8.227469, 
    8.238565, 8.250232, 8.283431, 8.313443, 8.346262, 8.354307, 8.392823, 
    8.361465, 8.413268, 8.369218, 8.445583, 8.308752, 8.367917, 8.260966, 
    8.272434, 8.293214, 8.341022, 8.315181, 8.345407, 8.278773, 8.244374, 
    8.235489, 8.218939, 8.235868, 8.234489, 8.250712, 8.245497, 8.284535, 
    8.263547, 8.323281, 8.345167, 8.407215, 8.445436, 8.484475, 8.501758, 
    8.507023, 8.509225,
  12.66552, 12.72099, 12.71019, 12.75506, 12.73015, 12.75956, 12.67674, 
    12.7232, 12.69352, 12.6705, 12.84257, 12.75706, 12.93193, 12.87698, 
    13.01541, 12.92337, 13.03404, 13.01274, 13.07694, 13.05852, 13.14096, 
    13.08545, 13.18388, 13.12768, 13.13646, 13.08362, 12.77422, 12.83189, 
    12.77081, 12.77902, 12.77534, 12.73066, 12.70821, 12.66129, 12.66979, 
    12.70426, 12.78271, 12.75603, 12.82337, 12.82185, 12.8972, 12.86318, 
    12.99045, 12.95416, 13.05929, 13.03277, 13.05804, 13.05037, 13.05814, 
    13.01928, 13.03592, 13.00176, 12.86954, 12.90827, 12.79309, 12.72429, 
    12.67878, 12.64658, 12.65113, 12.6598, 12.70446, 12.74658, 12.77876, 
    12.80034, 12.82163, 12.88628, 12.92061, 12.9978, 12.98384, 13.0075, 
    13.03014, 13.06824, 13.06196, 13.07877, 13.00687, 13.05462, 12.97589, 
    12.99738, 12.82744, 12.76322, 12.73603, 12.71226, 12.65462, 12.6944, 
    12.67871, 12.71607, 12.73987, 12.72809, 12.80093, 12.77257, 12.92265, 
    12.8578, 13.0275, 12.9867, 13.03729, 13.01145, 13.05576, 13.01588, 
    13.08503, 13.10013, 13.08981, 13.1295, 13.01367, 13.05804, 12.72777, 
    12.72968, 12.73863, 12.69935, 12.69695, 12.66105, 12.69299, 12.70661, 
    12.74125, 12.76178, 12.78133, 12.8244, 12.87267, 12.94045, 12.98934, 
    13.02221, 13.00205, 13.01985, 12.99995, 12.99063, 13.09447, 13.03607, 
    13.12378, 13.11891, 13.07917, 13.11946, 12.73103, 12.71999, 12.68172, 
    12.71166, 12.65715, 12.68764, 12.7052, 12.77316, 12.78814, 12.80204, 
    12.82954, 12.86492, 12.92719, 12.9816, 13.03146, 13.0278, 13.02909, 
    13.04025, 13.01262, 13.04479, 13.0502, 13.03606, 13.11826, 13.09473, 
    13.11881, 13.10348, 12.72358, 12.74217, 12.73212, 12.75103, 12.73771, 
    12.79704, 12.81489, 12.89867, 12.86422, 12.91909, 12.86978, 12.87851, 
    12.92089, 12.87244, 12.9786, 12.90655, 13.04068, 12.96841, 13.04522, 
    13.03124, 13.05439, 13.07517, 13.10134, 13.14977, 13.13854, 13.17913, 
    12.76994, 12.79414, 12.79201, 12.81738, 12.83617, 12.87699, 12.94272, 
    12.91797, 12.96344, 12.97259, 12.90351, 12.94589, 12.81037, 12.83218, 
    12.81918, 12.77185, 12.92367, 12.84555, 12.99015, 12.94757, 13.0722, 
    13.01009, 13.13236, 13.18496, 13.23463, 13.29292, 12.80737, 12.7909, 
    12.8204, 12.86132, 12.89939, 12.95017, 12.95537, 12.96491, 12.98964, 
    13.01047, 12.96793, 13.0157, 12.83725, 12.93047, 12.78468, 12.82843, 
    12.8589, 12.84552, 12.91514, 12.9316, 12.99869, 12.96397, 13.17197, 
    13.07957, 13.33744, 13.26491, 12.78515, 12.80731, 12.88471, 12.84783, 
    12.95356, 12.97971, 13.001, 13.02827, 13.03122, 13.0474, 13.02089, 
    13.04635, 12.95027, 12.99313, 12.87584, 12.9043, 12.8912, 12.87684, 
    12.92119, 12.9686, 12.96961, 12.98484, 13.02789, 12.95399, 13.18395, 
    13.0415, 12.83151, 12.87438, 12.8805, 12.86388, 12.97709, 12.93596, 
    13.04701, 13.01691, 13.06626, 13.04171, 13.03811, 13.00665, 12.98711, 
    12.93785, 12.89789, 12.86629, 12.87363, 12.90837, 12.9715, 13.03149, 
    13.01833, 13.0625, 12.94587, 12.99466, 12.97578, 13.02505, 12.91731, 
    13.00903, 12.89397, 12.90402, 12.93515, 12.99798, 13.01191, 13.02681, 
    13.01761, 12.97311, 12.96583, 12.93439, 12.92572, 12.90183, 12.88208, 
    12.90012, 12.9191, 12.97312, 13.02199, 13.07546, 13.08858, 13.15139, 
    13.10025, 13.18475, 13.11289, 13.2375, 13.01435, 13.11077, 12.93656, 
    12.95522, 12.98905, 13.06693, 13.02482, 13.07407, 12.96554, 12.90957, 
    12.89512, 12.86821, 12.89573, 12.89349, 12.91988, 12.9114, 12.97492, 
    12.94076, 13.03802, 13.07368, 13.17487, 13.23726, 13.30105, 13.3293, 
    13.33791, 13.34151,
  20.5999, 20.69597, 20.67725, 20.75504, 20.71184, 20.76284, 20.61933, 
    20.6998, 20.64839, 20.60852, 20.90694, 20.75851, 21.06236, 20.96676, 
    21.20783, 21.04745, 21.24033, 21.20317, 21.31522, 21.28305, 21.42712, 
    21.33008, 21.50222, 21.40389, 21.41924, 21.32689, 20.78828, 20.8884, 
    20.78236, 20.7966, 20.79021, 20.71274, 20.67383, 20.59257, 20.6073, 
    20.66698, 20.80301, 20.75671, 20.87359, 20.87094, 21.00193, 20.94276, 
    21.1643, 21.10106, 21.28439, 21.23812, 21.28222, 21.26883, 21.28239, 
    21.21457, 21.2436, 21.18403, 20.95382, 21.02119, 20.82101, 20.7017, 
    20.62286, 20.56712, 20.57499, 20.59, 20.66733, 20.74033, 20.79616, 
    20.8336, 20.87056, 20.98293, 21.04266, 21.17712, 21.15278, 21.19403, 
    21.23352, 21.30001, 21.28905, 21.31841, 21.19294, 21.27624, 21.13892, 
    21.17638, 20.88066, 20.76919, 20.72204, 20.68085, 20.58105, 20.64991, 
    20.62273, 20.68745, 20.7287, 20.70829, 20.83462, 20.78541, 21.04621, 
    20.93342, 21.22891, 21.15777, 21.246, 21.20092, 21.27823, 21.20864, 
    21.32934, 21.35573, 21.3377, 21.40707, 21.20479, 21.28222, 20.70772, 
    20.71104, 20.72655, 20.65848, 20.65433, 20.59217, 20.64746, 20.67106, 
    20.73109, 20.7667, 20.80061, 20.87539, 20.95927, 21.07719, 21.16237, 
    21.21969, 21.18452, 21.21557, 21.18087, 21.16462, 21.34584, 21.24387, 
    21.39707, 21.38856, 21.31911, 21.38952, 20.71338, 20.69424, 20.62794, 
    20.6798, 20.58541, 20.63819, 20.66861, 20.78644, 20.81242, 20.83656, 
    20.88431, 20.94578, 21.05411, 21.14888, 21.23582, 21.22943, 21.23168, 
    21.25116, 21.20296, 21.25908, 21.26852, 21.24385, 21.38742, 21.34629, 
    21.38838, 21.36159, 20.70046, 20.73269, 20.71527, 20.74804, 20.72495, 
    20.82788, 20.85886, 21.00448, 20.94457, 21.04, 20.95424, 20.96941, 
    21.04314, 20.95886, 21.14365, 21.01818, 21.25191, 21.1259, 21.25984, 
    21.23544, 21.27585, 21.31212, 21.35784, 21.44251, 21.42287, 21.4939, 
    20.78084, 20.82285, 20.81914, 20.86319, 20.89583, 20.96678, 21.08115, 
    21.03806, 21.11724, 21.13318, 21.01291, 21.08667, 20.85101, 20.88889, 
    20.86632, 20.78416, 21.04799, 20.91212, 21.16379, 21.0896, 21.30695, 
    21.19854, 21.41207, 21.50412, 21.59113, 21.69336, 20.84581, 20.81722, 
    20.86843, 20.93953, 21.00573, 21.09411, 21.10318, 21.11979, 21.16289, 
    21.19921, 21.12506, 21.20832, 20.8977, 21.05983, 20.80643, 20.88238, 
    20.93533, 20.91208, 21.03314, 21.06179, 21.17867, 21.11815, 21.48136, 
    21.3198, 21.77155, 21.64422, 20.80724, 20.84571, 20.9802, 20.91608, 
    21.10003, 21.14559, 21.1827, 21.23026, 21.2354, 21.26365, 21.21739, 
    21.26181, 21.0943, 21.16897, 20.96477, 21.01427, 20.99148, 20.96652, 
    21.04366, 21.12622, 21.12798, 21.15453, 21.22959, 21.10077, 21.50234, 
    21.25335, 20.88774, 20.96223, 20.97288, 20.94398, 21.14101, 21.06938, 
    21.26296, 21.21044, 21.29656, 21.25372, 21.24742, 21.19255, 21.15848, 
    21.07266, 21.00312, 20.94816, 20.96093, 21.02135, 21.13128, 21.23587, 
    21.21291, 21.29, 21.08663, 21.17164, 21.13874, 21.22465, 21.03692, 
    21.1967, 20.9963, 21.01378, 21.06796, 21.17743, 21.20172, 21.22771, 
    21.21167, 21.13408, 21.12139, 21.06664, 21.05156, 21.00997, 20.97562, 
    21.00701, 21.04003, 21.13411, 21.21931, 21.31264, 21.33555, 21.44535, 
    21.35593, 21.50374, 21.37803, 21.59616, 21.20598, 21.37432, 21.07043, 
    21.10292, 21.16186, 21.29773, 21.22425, 21.31021, 21.1209, 21.02345, 
    20.9983, 20.9515, 20.99937, 20.99547, 21.04139, 21.02662, 21.13724, 
    21.07774, 21.24727, 21.30952, 21.48644, 21.59574, 21.70763, 21.75724, 
    21.77237, 21.7787,
  34.64178, 34.82256, 34.7873, 34.9339, 34.85246, 34.94862, 34.67832, 
    34.82977, 34.73297, 34.65799, 35.22099, 34.94046, 35.51581, 35.33433, 
    35.79281, 35.48749, 35.85484, 35.78393, 35.99794, 35.93644, 36.21229, 
    36.02638, 36.3565, 36.16775, 36.19719, 36.02028, 34.99663, 35.18589, 
    34.98547, 35.01235, 35.00028, 34.85415, 34.78085, 34.62801, 34.65569, 
    34.76797, 35.02445, 34.93707, 35.15787, 35.15286, 35.40105, 35.28883, 
    35.70983, 35.58942, 35.939, 35.85061, 35.93484, 35.90927, 35.93518, 
    35.80567, 35.86108, 35.74743, 35.30981, 35.43761, 35.05846, 34.83335, 
    34.68494, 34.5802, 34.59498, 34.62318, 34.76863, 34.90616, 35.01151, 
    35.08224, 35.15214, 35.365, 35.47839, 35.73426, 35.68786, 35.7665, 
    35.84183, 35.96887, 35.94791, 36.00405, 35.76441, 35.92341, 35.66148, 
    35.73284, 35.17124, 34.96061, 34.87169, 34.79408, 34.60635, 34.73584, 
    34.68471, 34.80651, 34.88423, 34.84576, 35.08418, 34.99121, 35.48513, 
    35.27114, 35.83303, 35.69738, 35.86566, 35.77964, 35.92722, 35.79436, 
    36.02497, 36.07548, 36.04095, 36.17384, 35.78702, 35.93485, 34.84468, 
    34.85096, 34.88018, 34.75196, 34.74414, 34.62726, 34.73122, 34.77564, 
    34.88874, 34.9559, 35.01992, 35.16127, 35.32013, 35.54402, 35.70615, 
    35.81544, 35.74836, 35.80758, 35.74139, 35.71043, 36.05655, 35.8616, 
    36.15468, 36.13837, 36.00539, 36.14021, 34.85536, 34.81929, 34.6945, 
    34.7921, 34.61456, 34.71379, 34.77103, 34.99316, 35.04223, 35.08784, 
    35.17815, 35.29456, 35.50015, 35.68045, 35.84622, 35.83403, 35.83833, 
    35.87551, 35.78352, 35.89064, 35.90867, 35.86156, 36.13618, 36.05741, 
    36.13802, 36.0867, 34.83101, 34.89175, 34.85891, 34.92071, 34.87716, 
    35.07145, 35.13, 35.4059, 35.29227, 35.47334, 35.31059, 35.33936, 
    35.4793, 35.31936, 35.67049, 35.4319, 35.87695, 35.63669, 35.89209, 
    35.8455, 35.92268, 35.99202, 36.07952, 36.24184, 36.20415, 36.3405, 
    34.9826, 35.06193, 35.05492, 35.13819, 35.19995, 35.33437, 35.55154, 
    35.46964, 35.6202, 35.65054, 35.42189, 35.56203, 35.11515, 35.18681, 
    35.14411, 34.98885, 35.48851, 35.2308, 35.70884, 35.5676, 35.98212, 
    35.7751, 36.18343, 36.36015, 36.52758, 36.7248, 35.10532, 35.05129, 
    35.14811, 35.28272, 35.40826, 35.5762, 35.59344, 35.62506, 35.70713, 
    35.77637, 35.63508, 35.79375, 35.20348, 35.511, 35.03091, 35.17449, 
    35.27476, 35.23071, 35.4603, 35.51473, 35.73722, 35.62194, 36.31643, 
    36.00671, 36.876, 36.62993, 35.03245, 35.10513, 35.35983, 35.2383, 
    35.58744, 35.67417, 35.74489, 35.83562, 35.84542, 35.89936, 35.81104, 
    35.89586, 35.57656, 35.71873, 35.33056, 35.42447, 35.38122, 35.33387, 
    35.4803, 35.6373, 35.64064, 35.69121, 35.83433, 35.58887, 36.35673, 
    35.87968, 35.18464, 35.32574, 35.34594, 35.29114, 35.66546, 35.52916, 
    35.89804, 35.79779, 35.96227, 35.8804, 35.86838, 35.76368, 35.69873, 
    35.5354, 35.40332, 35.29908, 35.32327, 35.43792, 35.64693, 35.84632, 
    35.80251, 35.94973, 35.56196, 35.72381, 35.66113, 35.8249, 35.46748, 
    35.77157, 35.39036, 35.42354, 35.52647, 35.73484, 35.78116, 35.83075, 
    35.80013, 35.65226, 35.62811, 35.52395, 35.49529, 35.41631, 35.35114, 
    35.41068, 35.47338, 35.65231, 35.81471, 35.99301, 36.03684, 36.24728, 
    36.07586, 36.35942, 36.11818, 36.53728, 35.78928, 36.11108, 35.53115, 
    35.59296, 35.70518, 35.96449, 35.82413, 35.98836, 35.62716, 35.44189, 
    35.39416, 35.3054, 35.39619, 35.3888, 35.47597, 35.44792, 35.65827, 
    35.54505, 35.86808, 35.98705, 36.32619, 36.53647, 36.75238, 36.84832, 
    36.87759, 36.88984,
  60.67866, 61.07138, 60.99464, 61.31427, 61.13654, 61.34644, 60.75787, 
    61.08709, 60.87651, 60.71379, 61.94415, 61.3286, 62.59654, 62.19429, 
    63.21474, 62.53363, 63.35389, 63.19484, 63.67592, 63.53733, 64.16097, 
    63.74009, 64.48915, 64.05992, 64.12669, 63.72631, 61.45146, 61.86686, 
    61.42703, 61.48588, 61.45945, 61.14022, 60.9806, 60.64882, 60.70879, 
    60.95258, 61.51238, 61.32119, 61.80522, 61.7942, 62.34192, 62.09377, 
    63.02899, 62.76031, 63.54311, 63.34439, 63.53375, 63.4762, 63.5345, 
    63.24357, 63.36789, 63.11309, 62.1401, 62.42293, 61.58691, 61.09489, 
    60.77224, 60.54533, 60.5773, 60.63837, 60.95401, 61.2537, 61.48405, 
    61.6391, 61.79262, 62.26212, 62.51342, 63.08363, 62.97991, 63.15579, 
    63.32469, 63.61038, 63.56317, 63.68969, 63.15111, 63.50803, 62.92099, 
    63.08046, 61.83464, 61.37265, 61.17847, 61.00938, 60.60192, 60.88274, 
    60.77174, 61.03644, 61.20583, 61.12193, 61.64335, 61.4396, 62.52837, 
    62.05472, 63.30494, 63.00117, 63.37819, 63.18523, 63.5166, 63.21821, 
    63.7369, 63.85101, 63.77299, 64.07372, 63.20175, 63.53376, 61.11959, 
    61.13326, 61.197, 60.91779, 60.90078, 60.64719, 60.87272, 60.96927, 
    61.21567, 61.36237, 61.50245, 61.81269, 62.16289, 62.65925, 63.02077, 
    63.26548, 63.11519, 63.24784, 63.0996, 63.03035, 63.80822, 63.36906, 
    64.03029, 63.99333, 63.69271, 63.99749, 61.14286, 61.06427, 60.79298, 
    61.00508, 60.61969, 60.83485, 60.95924, 61.44387, 61.55134, 61.65136, 
    61.84983, 62.10643, 62.56173, 62.96335, 63.33453, 63.30719, 63.31681, 
    63.40031, 63.19391, 63.43432, 63.47487, 63.36899, 63.98838, 63.81017, 
    63.99254, 63.87637, 61.08979, 61.22225, 61.1506, 61.28547, 61.19041, 
    61.6154, 61.74396, 62.35265, 62.10136, 62.5022, 62.14183, 62.20539, 
    62.51543, 62.16119, 62.9411, 62.41028, 63.40356, 62.86567, 63.43758, 
    63.33292, 63.50638, 63.66257, 63.86015, 64.22809, 64.14249, 64.45267, 
    61.42075, 61.59453, 61.57916, 61.76195, 61.89783, 62.19437, 62.67599, 
    62.494, 62.8289, 62.89658, 62.38808, 62.69933, 61.71135, 61.86889, 
    61.77497, 61.43444, 62.53588, 61.96577, 63.02679, 62.71174, 63.64025, 
    63.17506, 64.09548, 64.49747, 64.88044, 65.3342, 61.68975, 61.57121, 
    61.78375, 62.08028, 62.35789, 62.73087, 62.76927, 62.83974, 63.02298, 
    63.1779, 62.86208, 63.21685, 61.9056, 62.58585, 61.52654, 61.84178, 
    62.06271, 61.96557, 62.47326, 62.59414, 63.09025, 62.83279, 64.3978, 
    63.6957, 65.68405, 65.11556, 61.5299, 61.68932, 62.25066, 61.98231, 
    62.75591, 62.94933, 63.10743, 63.31075, 63.33276, 63.45393, 63.25561, 
    63.44606, 62.73167, 63.04889, 62.18595, 62.39381, 62.298, 62.19328, 
    62.51765, 62.86703, 62.87449, 62.9874, 63.30784, 62.75908, 64.48967, 
    63.4097, 61.8641, 62.17531, 62.21996, 62.09887, 62.92989, 62.62622, 
    63.45097, 63.22589, 63.59551, 63.4113, 63.38429, 63.14947, 63.00418, 
    62.64008, 62.34694, 62.1164, 62.16985, 62.42362, 62.88852, 63.33477, 
    63.23648, 63.56726, 62.69917, 63.06026, 62.92022, 63.2867, 62.48919, 
    63.16716, 62.31825, 62.39175, 62.62022, 63.08494, 63.18863, 63.29981, 
    63.23115, 62.90041, 62.84653, 62.61464, 62.55093, 62.37573, 62.23145, 
    62.36326, 62.5023, 62.90052, 63.26383, 63.6648, 63.7637, 64.24046, 
    63.85188, 64.4958, 63.9476, 64.90269, 63.20683, 63.93153, 62.63064, 
    62.7682, 63.0186, 63.60052, 63.28497, 63.6543, 62.84442, 62.43243, 
    62.32666, 62.13037, 62.33117, 62.31479, 62.50804, 62.4458, 62.91383, 
    62.66155, 63.38363, 63.65136, 64.42004, 64.90083, 65.39787, 65.61987, 
    65.68774, 65.71616,
  116.3177, 117.5456, 117.3041, 118.3152, 117.7513, 118.4177, 116.5638, 
    117.5952, 116.9339, 116.4268, 120.3482, 118.3608, 122.5137, 121.1711, 
    124.6258, 122.3021, 125.1096, 124.5568, 126.2418, 125.7524, 127.9808, 
    126.4695, 129.1813, 127.6151, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9487, 118.3372, 119.895, 119.8592, 121.661, 120.8393, 
    123.9848, 123.0674, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7258, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9053, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3958, 122.2342, 124.1728, 123.8164, 124.4217, 
    125.0078, 126.01, 125.8434, 126.2906, 124.4056, 125.6494, 123.6147, 
    124.1619, 119.9907, 118.5013, 117.8839, 117.3505, 116.0801, 116.9533, 
    116.607, 117.4356, 117.9707, 117.7052, 119.3704, 118.7153, 122.2845, 
    120.7108, 124.9391, 123.8893, 125.1945, 124.5236, 125.6795, 124.6378, 
    126.4582, 126.8648, 126.5865, 127.6649, 124.5808, 125.7399, 117.6978, 
    117.741, 117.9427, 117.063, 117.0098, 116.2202, 116.922, 117.2245, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9566, 
    124.8018, 124.2816, 124.7406, 124.2278, 123.9895, 126.712, 125.1626, 
    127.5082, 127.3751, 126.3013, 127.3901, 117.7713, 117.5232, 116.6731, 
    117.337, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.881, 122.3966, 123.7596, 125.0421, 124.9469, 124.9804, 
    125.2718, 124.5536, 125.3908, 125.5329, 125.1623, 127.3573, 126.719, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9218, 
    119.2802, 119.696, 121.6967, 120.8643, 122.1966, 120.9977, 121.2078, 
    122.241, 121.0616, 123.6834, 121.889, 125.2831, 123.4258, 125.4022, 
    125.0365, 125.6436, 126.1945, 126.8974, 128.2247, 127.9138, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1968, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8149, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3097, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4884, 127.7436, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7949, 121.7142, 122.9675, 123.0978, 123.3374, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.014, 
    120.7371, 120.4183, 122.0996, 122.5056, 124.1956, 123.3137, 128.8452, 
    126.3119, 133.7281, 131.5293, 119.005, 119.5191, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2548, 124.9593, 125.0359, 125.4595, 124.7676, 
    125.4319, 122.9702, 124.0532, 121.1435, 121.834, 121.5149, 121.1677, 
    122.2484, 123.4304, 123.4559, 123.842, 124.9492, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1083, 121.256, 120.8561, 123.6451, 122.6137, 
    125.4491, 124.6645, 125.9575, 125.3102, 125.2158, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.043, 
    124.7011, 125.8578, 122.8602, 124.0923, 123.612, 124.8756, 122.153, 
    124.4611, 121.5822, 121.8271, 122.5935, 124.1773, 124.5353, 124.9212, 
    124.6827, 123.5443, 123.3605, 122.5747, 122.3602, 121.7737, 121.2941, 
    121.7321, 122.197, 123.5447, 124.7961, 126.2024, 126.5535, 128.2698, 
    126.8678, 129.2059, 127.2107, 130.7229, 124.5984, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9752, 124.8696, 126.1653, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5902, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6129, 133.4765, 
    133.7426, 133.8544,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02028661, -0.01995555, -0.02001946, -0.01975575, -0.01990158, 
    -0.01972957, -0.02021903, -0.01994251, -0.02011857, -0.02025658, 
    -0.01925455, -0.01974408, -0.01876002, -0.01906207, -0.01831312, 
    -0.01880666, -0.01821532, -0.0183272, -0.01799279, -0.01808791, 
    -0.01766731, -0.01794907, -0.01745352, -0.01773418, -0.01768994, 
    -0.01795844, -0.01964453, -0.01931477, -0.01966425, -0.01961681, 
    -0.01963809, -0.01989855, -0.02003119, -0.02031218, -0.02026086, 
    -0.02005464, -0.01959551, -0.01975011, -0.01936305, -0.0193717, 
    -0.01895016, -0.01913898, -0.01844525, -0.01863963, -0.01808393, 
    -0.01822197, -0.01809038, -0.01813018, -0.01808986, -0.01829278, 
    -0.01820554, -0.01838521, -0.01910346, -0.01888927, -0.01953586, 
    -0.01993605, -0.02020681, -0.02040132, -0.0203737, -0.02032115, 
    -0.02005344, -0.01980523, -0.01961828, -0.01949429, -0.01937295, 
    -0.01901049, -0.01882169, -0.0184062, -0.01848047, -0.01835486, 
    -0.01823577, -0.01803765, -0.0180701, -0.01798338, -0.01835819, 
    -0.01810815, -0.01852292, -0.01840846, -0.01933998, -0.01970828, 
    -0.019867, -0.02000715, -0.02035249, -0.02011332, -0.02020724, 
    -0.0199846, -0.01984449, -0.01991366, -0.01949091, -0.0196541, 
    -0.01881056, -0.01916902, -0.01824961, -0.0184652, -0.01819835, 
    -0.018334, -0.01810222, -0.01831068, -0.01795123, -0.01787397, 
    -0.01792673, -0.01772502, -0.0183223, -0.01809037, -0.0199156, 
    -0.01990429, -0.01985175, -0.02008383, -0.02009813, -0.02031358, 
    -0.02012176, -0.02004066, -0.01983641, -0.01971663, -0.01960349, 
    -0.01935719, -0.01908603, -0.01871374, -0.01845114, -0.01827735, 
    -0.01838371, -0.01828977, -0.01839482, -0.01844428, -0.01790287, 
    -0.01820472, -0.01775388, -0.01777851, -0.01798132, -0.01777573, 
    -0.01989637, -0.01996146, -0.0201892, -0.02001074, -0.02033719, 
    -0.02015374, -0.02004906, -0.01965065, -0.01956429, -0.01948454, 
    -0.01932809, -0.01912927, -0.0187858, -0.01849238, -0.01822887, 
    -0.01824804, -0.01824128, -0.01818292, -0.01832785, -0.01815925, 
    -0.0181311, -0.01820477, -0.01778181, -0.01790155, -0.01777903, 
    -0.01785689, -0.01994028, -0.01983101, -0.01988997, -0.01977925, 
    -0.01985718, -0.01951315, -0.01941125, -0.01894207, -0.01913316, 
    -0.01883004, -0.01910214, -0.01905361, -0.01882019, -0.01908733, 
    -0.01850841, -0.01889875, -0.01818066, -0.01856294, -0.01815698, 
    -0.01823, -0.01810929, -0.01800191, -0.01786781, -0.01762318, 
    -0.01767951, -0.01747704, -0.01966932, -0.01952978, -0.01954205, 
    -0.01939707, -0.0192906, -0.01906201, -0.01870143, -0.01883616, 
    -0.01858964, -0.01854056, -0.01891541, -0.01868428, -0.01943701, 
    -0.01931319, -0.01938682, -0.01965826, -0.01880499, -0.01923778, 
    -0.01844683, -0.01867518, -0.01801717, -0.0183412, -0.01771059, 
    -0.01744816, -0.01720512, -0.01692564, -0.0194541, -0.0195484, 
    -0.01937992, -0.01914935, -0.01893812, -0.01866116, -0.01863308, 
    -0.01858176, -0.01844956, -0.01833919, -0.01856555, -0.01831163, 
    -0.01928455, -0.01876793, -0.01958416, -0.01933439, -0.01916287, 
    -0.01923793, -0.01885163, -0.0187618, -0.01840148, -0.01858681, 
    -0.01751252, -0.01797928, -0.01671622, -0.01705918, -0.01958146, 
    -0.01945443, -0.01901919, -0.01922496, -0.01864284, -0.01850248, 
    -0.01838924, -0.01824554, -0.01823011, -0.01814562, -0.01828429, 
    -0.01815109, -0.01866058, -0.01843101, -0.01906843, -0.01891111, 
    -0.01898332, -0.01906284, -0.01881855, -0.01856195, -0.01855655, 
    -0.01847509, -0.01824757, -0.01864052, -0.01745318, -0.01817637, 
    -0.01931693, -0.01907655, -0.01904252, -0.01913507, -0.0185165, 
    -0.01873809, -0.01814768, -0.01830525, -0.01804786, -0.01817526, 
    -0.01819409, -0.01835935, -0.01846304, -0.01872787, -0.01894637, 
    -0.01912162, -0.01908072, -0.01888875, -0.01854639, -0.0182287, 
    -0.01829778, -0.01806728, -0.0186844, -0.01842288, -0.01852348, 
    -0.01826242, -0.01883974, -0.01834679, -0.01896801, -0.01891266, 
    -0.01874252, -0.01840526, -0.01833159, -0.01825322, -0.01830154, 
    -0.01853779, -0.01857683, -0.01874665, -0.01879381, -0.0189247, 
    -0.01903379, -0.01893408, -0.01882997, -0.01853771, -0.0182785, 
    -0.01800038, -0.01793303, -0.01761506, -0.01787339, -0.01744924, 
    -0.01780907, -0.01719121, -0.01831871, -0.01781984, -0.01873483, 
    -0.01863387, -0.0184527, -0.01804441, -0.01826364, -0.01800755, 
    -0.01857836, -0.01888215, -0.01896166, -0.01911091, -0.01895826, 
    -0.01897063, -0.01882569, -0.01887214, -0.01852809, -0.01871205, 
    -0.01819455, -0.01800957, -0.01749812, -0.01719238, -0.01688715, 
    -0.01675426, -0.01671404, -0.01669725,
  -0.05424561, -0.05319658, -0.05339885, -0.05256495, -0.05302586, 
    -0.05248226, -0.05403123, -0.05315533, -0.05371277, -0.05415035, 
    -0.05098546, -0.05252808, -0.04943406, -0.05038077, -0.04803829, 
    -0.04958008, -0.04773362, -0.04808215, -0.04704147, -0.04733715, 
    -0.04603188, -0.04690566, -0.04537049, -0.04623903, -0.04610197, 
    -0.04693477, -0.05221383, -0.05117485, -0.05227605, -0.05212636, 
    -0.0521935, -0.05301626, -0.05343598, -0.05432675, -0.0541639, 
    -0.05351026, -0.0520592, -0.05254713, -0.05132678, -0.05135401, 
    -0.05002971, -0.05062228, -0.04845035, -0.04905746, -0.04732477, 
    -0.04775432, -0.04734484, -0.04746862, -0.04734323, -0.04797489, 
    -0.04770316, -0.04826302, -0.05051072, -0.04983884, -0.05187109, 
    -0.05313487, -0.05399247, -0.0546098, -0.05452207, -0.05435523, 
    -0.05350646, -0.05272127, -0.05213102, -0.05174008, -0.05135792, 
    -0.05021893, -0.04962715, -0.0483285, -0.04856027, -0.04816839, 
    -0.04779728, -0.04718089, -0.04728178, -0.04701226, -0.04817876, 
    -0.04740009, -0.04869279, -0.04833554, -0.05125417, -0.05241504, 
    -0.05291651, -0.05335989, -0.05445472, -0.05369613, -0.05399383, 
    -0.05328851, -0.05284534, -0.05306406, -0.05172944, -0.05224403, 
    -0.0495923, -0.05071663, -0.04784041, -0.04851261, -0.04768078, 
    -0.04810335, -0.04738167, -0.04803066, -0.04691239, -0.04667253, 
    -0.0468363, -0.04621063, -0.0480669, -0.04734481, -0.05307018, 
    -0.05303444, -0.0528683, -0.05360271, -0.05364801, -0.05433121, 
    -0.05372288, -0.05346599, -0.0528198, -0.0524414, -0.05208435, 
    -0.05130833, -0.050456, -0.04928926, -0.04846873, -0.0479268, 
    -0.04825836, -0.04796551, -0.04829299, -0.04844731, -0.04676223, 
    -0.04770061, -0.04630008, -0.04637643, -0.04700585, -0.04636782, 
    -0.05300936, -0.05321528, -0.05393665, -0.05337124, -0.05440616, 
    -0.05382423, -0.05349258, -0.05223314, -0.05196073, -0.05170936, 
    -0.05121676, -0.05059177, -0.04951476, -0.04859745, -0.0477758, 
    -0.04783551, -0.04781447, -0.04763275, -0.04808418, -0.04755907, 
    -0.0474715, -0.04770077, -0.04638667, -0.04675814, -0.04637806, 
    -0.04661953, -0.05314826, -0.05280274, -0.05298914, -0.05263917, 
    -0.05288545, -0.0517995, -0.05147852, -0.05000434, -0.05060397, 
    -0.0496533, -0.05050656, -0.05035422, -0.04962245, -0.05046008, 
    -0.04864749, -0.04986856, -0.0476257, -0.0488178, -0.04755202, 
    -0.04777932, -0.04740365, -0.04706981, -0.04665342, -0.04589524, 
    -0.04606965, -0.04544317, -0.05229207, -0.05185194, -0.0518906, 
    -0.05143388, -0.05109882, -0.05038058, -0.04925073, -0.04967244, 
    -0.04890121, -0.04874789, -0.04992079, -0.04919709, -0.05155962, 
    -0.05116987, -0.0514016, -0.05225717, -0.04957483, -0.05093272, 
    -0.04845528, -0.04916863, -0.04711725, -0.0481258, -0.04616595, 
    -0.04535395, -0.04460386, -0.04374361, -0.05161346, -0.05191064, 
    -0.05137987, -0.05065484, -0.04999197, -0.04912479, -0.04903701, 
    -0.04887661, -0.0484638, -0.04811953, -0.04882594, -0.04803364, 
    -0.05107979, -0.04945882, -0.05202339, -0.05123658, -0.0506973, 
    -0.0509332, -0.04972091, -0.04943962, -0.04831377, -0.04889238, 
    -0.04555288, -0.04699952, -0.04310065, -0.04415433, -0.05201487, 
    -0.05161452, -0.05024622, -0.05089242, -0.04906751, -0.04862898, 
    -0.0482756, -0.04782772, -0.04777968, -0.04751668, -0.04794845, 
    -0.04753368, -0.04912296, -0.04840591, -0.05040074, -0.0499073, 
    -0.05013369, -0.05038321, -0.04961729, -0.04881472, -0.04879783, 
    -0.04854348, -0.04783406, -0.04906026, -0.04536945, -0.04761238, 
    -0.05118165, -0.05042623, -0.05031943, -0.05060997, -0.04867275, 
    -0.04936545, -0.04752309, -0.04801374, -0.04721263, -0.04760892, 
    -0.04766752, -0.04818238, -0.04850586, -0.04933343, -0.05001784, 
    -0.05056774, -0.05043931, -0.04983722, -0.0487661, -0.04777528, 
    -0.04799047, -0.04727301, -0.04919747, -0.04838054, -0.04869454, 
    -0.04788031, -0.04968368, -0.04814325, -0.05008569, -0.04991214, 
    -0.0493793, -0.04832558, -0.04809585, -0.04785163, -0.04800219, 
    -0.04873925, -0.04886119, -0.0493922, -0.04953984, -0.04994988, 
    -0.05029202, -0.0499793, -0.04965307, -0.04873898, -0.04793041, 
    -0.04706506, -0.04685586, -0.04587012, -0.04667073, -0.04535725, 
    -0.04647119, -0.04456096, -0.0480557, -0.0465046, -0.04935523, 
    -0.04903945, -0.04847359, -0.04720191, -0.04788411, -0.04708736, 
    -0.04886598, -0.04981653, -0.05006577, -0.0505341, -0.05005512, 
    -0.0500939, -0.04963968, -0.04978518, -0.04870894, -0.04928396, 
    -0.04766896, -0.04709362, -0.04550836, -0.04456457, -0.04362532, 
    -0.04321733, -0.04309396, -0.0430425,
  -0.07888652, -0.07723158, -0.0775505, -0.07623623, -0.07696247, -0.076106, 
    -0.07854813, -0.07716656, -0.07804563, -0.07873614, -0.07375098, 
    -0.07617816, -0.07131527, -0.07280098, -0.06912857, -0.07154429, 
    -0.06865185, -0.06919722, -0.06756967, -0.06803183, -0.06599323, 
    -0.06735747, -0.06496184, -0.06631649, -0.06610259, -0.06740295, 
    -0.07568329, -0.07404868, -0.07578127, -0.07554559, -0.07565129, 
    -0.07694734, -0.07760905, -0.07901463, -0.07875753, -0.07772619, 
    -0.07543988, -0.07620817, -0.07428756, -0.07433038, -0.0722498, 
    -0.0731803, -0.06977365, -0.07072483, -0.06801248, -0.06868424, 
    -0.06804386, -0.06823739, -0.06804134, -0.06902935, -0.06860421, 
    -0.06948034, -0.07300506, -0.07195025, -0.07514382, -0.0771343, 
    -0.07848696, -0.0794616, -0.07932305, -0.0790596, -0.0777202, 
    -0.07648248, -0.07555293, -0.07493766, -0.07433654, -0.07254685, 
    -0.07161812, -0.06958286, -0.0699458, -0.06933221, -0.06875145, 
    -0.06778757, -0.06794526, -0.06752402, -0.06934843, -0.06813025, 
    -0.07015339, -0.06959389, -0.07417341, -0.07600013, -0.07679013, 
    -0.07748907, -0.07921669, -0.07801938, -0.0784891, -0.07737651, 
    -0.07667799, -0.07702267, -0.07492092, -0.07573085, -0.07156347, 
    -0.07332853, -0.06881893, -0.06987116, -0.06856919, -0.06923041, 
    -0.06810144, -0.06911663, -0.06736799, -0.0669933, -0.0672491, 
    -0.06627217, -0.06917335, -0.06804381, -0.07703232, -0.07697599, 
    -0.07671416, -0.07787202, -0.07794347, -0.07902166, -0.07806159, 
    -0.07765638, -0.07663774, -0.07604163, -0.07547947, -0.07425856, 
    -0.07291912, -0.07108821, -0.06980244, -0.0689541, -0.06947305, 
    -0.06901468, -0.06952727, -0.06976891, -0.0671334, -0.06860023, 
    -0.06641176, -0.06653097, -0.06751402, -0.06651752, -0.07693646, 
    -0.07726105, -0.07839886, -0.07750696, -0.07914001, -0.07822149, 
    -0.07769831, -0.07571369, -0.07528488, -0.07488934, -0.07411458, 
    -0.07313237, -0.07144184, -0.07000404, -0.06871784, -0.06881125, 
    -0.06877834, -0.06849407, -0.0692004, -0.06837884, -0.0682419, 
    -0.06860047, -0.06654694, -0.06712701, -0.0665335, -0.06691053, 
    -0.0771554, -0.07661085, -0.07690459, -0.07635316, -0.07674117, 
    -0.07503116, -0.07452621, -0.07220999, -0.07315154, -0.07165914, 
    -0.07299853, -0.07275929, -0.07161076, -0.07292552, -0.07008242, 
    -0.0719969, -0.06848305, -0.07034925, -0.06836782, -0.06872335, 
    -0.0681358, -0.06761396, -0.06696346, -0.06578006, -0.06605216, 
    -0.06507512, -0.07580648, -0.07511368, -0.07517452, -0.074456, 
    -0.07392918, -0.07280067, -0.07102779, -0.07168919, -0.07047994, 
    -0.07023972, -0.07207885, -0.07094371, -0.07465377, -0.07404087, 
    -0.07440524, -0.07575153, -0.07153606, -0.07366809, -0.06978138, 
    -0.07089909, -0.0676881, -0.06926554, -0.06620243, -0.06493605, 
    -0.06376769, -0.06242949, -0.07473847, -0.07520604, -0.07437106, 
    -0.07323145, -0.07219058, -0.07083037, -0.07069276, -0.0704414, 
    -0.06979471, -0.06925572, -0.07036201, -0.06912129, -0.07389925, 
    -0.0713541, -0.07538351, -0.07414576, -0.07329817, -0.07366884, 
    -0.07176521, -0.07132399, -0.06955981, -0.07046612, -0.06524616, 
    -0.06750413, -0.06143053, -0.06306817, -0.0753701, -0.07474012, 
    -0.07258969, -0.07360476, -0.07074057, -0.07005343, -0.06950004, 
    -0.06879908, -0.06872392, -0.06831256, -0.06898798, -0.06833914, 
    -0.0708275, -0.06970408, -0.07283233, -0.07205769, -0.07241302, 
    -0.0728048, -0.07160266, -0.07034442, -0.07031796, -0.0699195, 
    -0.06880899, -0.07072921, -0.06496022, -0.06846222, -0.07405937, 
    -0.07287236, -0.07270464, -0.07316097, -0.070122, -0.07120766, 
    -0.06832257, -0.06909016, -0.06783717, -0.06845681, -0.06854846, 
    -0.06935409, -0.06986059, -0.07115748, -0.07223117, -0.07309463, 
    -0.07289291, -0.07194772, -0.07026824, -0.06871704, -0.06905374, 
    -0.06793156, -0.07094429, -0.06966434, -0.07015613, -0.06888136, 
    -0.07170681, -0.06929285, -0.07233769, -0.07206529, -0.0712294, 
    -0.06957829, -0.06921865, -0.06883649, -0.06907208, -0.07022618, 
    -0.07041723, -0.07124963, -0.07148118, -0.07212451, -0.07266161, 
    -0.07217068, -0.07165879, -0.07022575, -0.06895975, -0.06760654, 
    -0.06727967, -0.06574088, -0.06699049, -0.06494121, -0.0666789, 
    -0.06370091, -0.06915583, -0.06673106, -0.07119166, -0.0706966, 
    -0.06981005, -0.06782043, -0.0688873, -0.06764139, -0.07042474, 
    -0.07191525, -0.07230642, -0.0730418, -0.0722897, -0.07235057, 
    -0.07163779, -0.07186606, -0.07017869, -0.07107989, -0.06855072, 
    -0.06765118, -0.06517676, -0.06370652, -0.06224562, -0.06161173, 
    -0.06142015, -0.06134024,
  -0.08614745, -0.08423818, -0.08460601, -0.08309054, -0.08392785, 
    -0.08294041, -0.08575694, -0.0841632, -0.08517716, -0.0859739, 
    -0.08022729, -0.0830236, -0.07742436, -0.07913367, -0.07491082, 
    -0.07768777, -0.07436323, -0.07498969, -0.07312064, -0.07365122, 
    -0.07131182, -0.07287706, -0.07012921, -0.07168259, -0.07143723, 
    -0.07292926, -0.08245321, -0.08057011, -0.08256613, -0.08229453, 
    -0.08241633, -0.0839104, -0.08467355, -0.08629531, -0.08599859, 
    -0.08480866, -0.08217271, -0.08305819, -0.08084521, -0.08089452, 
    -0.07849939, -0.07957028, -0.07565203, -0.07674539, -0.073629, 
    -0.07440042, -0.07366502, -0.07388725, -0.07366213, -0.07479684, 
    -0.07430851, -0.07531499, -0.07936856, -0.07815475, -0.08183157, 
    -0.084126, -0.08568637, -0.08681123, -0.0866513, -0.08634721, 
    -0.08480175, -0.08337442, -0.08230299, -0.08159406, -0.08090162, 
    -0.07884121, -0.07777269, -0.07543279, -0.07584988, -0.07514479, 
    -0.07447762, -0.07337077, -0.07355182, -0.07306824, -0.07516342, 
    -0.07376422, -0.07608847, -0.07544546, -0.08071374, -0.08281839, 
    -0.08372913, -0.08453515, -0.08652852, -0.08514688, -0.08568884, 
    -0.08440533, -0.08359981, -0.08399726, -0.08157476, -0.08250801, 
    -0.07770982, -0.07974092, -0.07455512, -0.0757641, -0.07426829, 
    -0.07502782, -0.07373113, -0.0748971, -0.07288913, -0.07245912, 
    -0.07275269, -0.07163174, -0.07496227, -0.07366496, -0.0840084, 
    -0.08394343, -0.08364152, -0.08497688, -0.08505931, -0.08630342, 
    -0.08519557, -0.08472814, -0.08355342, -0.08286622, -0.08221833, 
    -0.0808118, -0.07926965, -0.07716323, -0.07568512, -0.07471039, 
    -0.0753066, -0.07477998, -0.07536891, -0.07564659, -0.07261991, 
    -0.07430393, -0.07179189, -0.07192864, -0.07305676, -0.07191321, 
    -0.08389786, -0.08427217, -0.08558471, -0.08455578, -0.08644002, 
    -0.08538005, -0.0847765, -0.08248825, -0.08199411, -0.08153838, 
    -0.08064598, -0.07951511, -0.07756992, -0.07591681, -0.07443902, 
    -0.07454631, -0.07450851, -0.07418202, -0.07499335, -0.07404967, 
    -0.07389243, -0.07430421, -0.07194696, -0.07261257, -0.07193154, 
    -0.07236414, -0.08415033, -0.08352242, -0.08386111, -0.08322532, 
    -0.08367268, -0.08170178, -0.08112007, -0.07845359, -0.07953718, 
    -0.07781987, -0.07936104, -0.07908568, -0.07776422, -0.07927702, 
    -0.0760069, -0.07820842, -0.07416935, -0.07631361, -0.07403702, 
    -0.07444534, -0.07377059, -0.07317148, -0.07242487, -0.07106733, 
    -0.0713794, -0.07025906, -0.0825952, -0.08179685, -0.08186694, 
    -0.08103921, -0.08043247, -0.07913332, -0.07709375, -0.07785442, 
    -0.07646386, -0.07618771, -0.0783027, -0.07699706, -0.08126701, 
    -0.08056109, -0.08098073, -0.08253186, -0.0776783, -0.08013185, 
    -0.07566091, -0.07694576, -0.07325658, -0.07506818, -0.07155176, 
    -0.07009964, -0.06876083, -0.0672285, -0.08136457, -0.08190326, 
    -0.08094137, -0.07962915, -0.07843125, -0.07686674, -0.07670853, 
    -0.07641953, -0.07567624, -0.0750569, -0.07632828, -0.07490247, 
    -0.08039802, -0.07746901, -0.08210775, -0.08068188, -0.07970596, 
    -0.08013272, -0.07794188, -0.07743438, -0.0754063, -0.07644796, 
    -0.07045514, -0.0730454, -0.0660854, -0.06795969, -0.0820923, 
    -0.08136648, -0.0788905, -0.08005892, -0.0767635, -0.07597358, 
    -0.07533762, -0.07453232, -0.07444599, -0.07397356, -0.07474931, 
    -0.07400409, -0.07686344, -0.07557207, -0.07916975, -0.07827836, 
    -0.0786872, -0.07913806, -0.0777549, -0.07630806, -0.07627764, 
    -0.07581966, -0.07454372, -0.07675043, -0.07012735, -0.07414544, 
    -0.08058241, -0.07921582, -0.07902279, -0.07954802, -0.07605239, 
    -0.07730061, -0.07398506, -0.07486669, -0.07342772, -0.07413922, 
    -0.07424447, -0.07516993, -0.07575195, -0.07724288, -0.07847796, 
    -0.07947166, -0.07923948, -0.07815184, -0.0762205, -0.0744381, 
    -0.07482486, -0.07353609, -0.07699774, -0.07552642, -0.07609162, 
    -0.07462684, -0.07787471, -0.07509957, -0.07860051, -0.07828709, 
    -0.07732559, -0.07542753, -0.07501432, -0.0745753, -0.07484592, 
    -0.07617214, -0.07639176, -0.07734887, -0.07761516, -0.07835524, 
    -0.07897326, -0.07840835, -0.07781947, -0.07617165, -0.07471689, 
    -0.07316296, -0.07278777, -0.0710224, -0.0724559, -0.07010557, 
    -0.07209837, -0.06868434, -0.07494214, -0.07215822, -0.07728219, 
    -0.07671294, -0.07569387, -0.07340851, -0.07463366, -0.07320297, 
    -0.07640039, -0.07811449, -0.07856454, -0.07941084, -0.07854529, 
    -0.07861535, -0.07779531, -0.07805789, -0.07611755, -0.07715367, 
    -0.07424707, -0.0732142, -0.07037557, -0.06869076, -0.06701805, 
    -0.0662927, -0.06607352, -0.06598211,
  -0.06724854, -0.06570274, -0.06600055, -0.06477354, -0.06545148, -0.064652, 
    -0.06693238, -0.06564203, -0.06646297, -0.06710804, -0.06245522, 
    -0.06471935, -0.06018564, -0.0615697, -0.05815036, -0.06039893, 
    -0.05770696, -0.05821422, -0.0567008, -0.05713043, -0.05523618, 
    -0.05650358, -0.05427864, -0.0555364, -0.05533773, -0.05654585, 
    -0.06425752, -0.0627328, -0.06434895, -0.06412905, -0.06422766, 
    -0.06543735, -0.06605524, -0.06736824, -0.06712802, -0.06616463, 
    -0.0640304, -0.06474736, -0.06295554, -0.06299547, -0.06105611, 
    -0.06192322, -0.05875054, -0.05963586, -0.05711243, -0.05773707, 
    -0.0571416, -0.05732155, -0.05713926, -0.05805806, -0.05766265, 
    -0.05847763, -0.06175989, -0.06077706, -0.06375419, -0.06561191, 
    -0.06687524, -0.06778593, -0.06765645, -0.06741027, -0.06615902, 
    -0.0650034, -0.06413589, -0.06356188, -0.06300122, -0.0613329, 
    -0.06046769, -0.05857301, -0.05891074, -0.05833981, -0.05779958, 
    -0.05690334, -0.05704994, -0.05665838, -0.0583549, -0.05722193, 
    -0.05910393, -0.05858327, -0.0628491, -0.06455319, -0.06529059, 
    -0.06594318, -0.06755706, -0.06643846, -0.06687724, -0.06583808, 
    -0.06518589, -0.06550768, -0.06354626, -0.06430189, -0.06041678, 
    -0.0620614, -0.05786234, -0.05884128, -0.05763008, -0.05824509, 
    -0.05719513, -0.05813925, -0.05651335, -0.05616517, -0.05640287, 
    -0.05549523, -0.05819201, -0.05714156, -0.0655167, -0.06546409, 
    -0.06521966, -0.06630082, -0.06636755, -0.06737481, -0.06647788, 
    -0.06609943, -0.06514832, -0.06459193, -0.06406734, -0.06292849, 
    -0.0616798, -0.0599742, -0.05877733, -0.05798807, -0.05847083, 
    -0.05804441, -0.05852128, -0.05874613, -0.05629535, -0.05765894, 
    -0.0556249, -0.05573562, -0.05664908, -0.05572313, -0.0654272, 
    -0.06573026, -0.06679294, -0.06595989, -0.06748541, -0.06662723, 
    -0.06613858, -0.0642859, -0.06388579, -0.0635168, -0.06279422, 
    -0.06187855, -0.0603035, -0.05896494, -0.05776833, -0.0578552, 
    -0.0578246, -0.05756022, -0.05821718, -0.05745307, -0.05732574, 
    -0.05765917, -0.05575046, -0.05628941, -0.05573798, -0.05608825, 
    -0.06563161, -0.06512322, -0.06539745, -0.06488267, -0.06524488, 
    -0.0636491, -0.06317811, -0.06101903, -0.06189642, -0.06050589, 
    -0.06175381, -0.06153084, -0.06046084, -0.06168577, -0.05903789, 
    -0.06082051, -0.05754997, -0.05928624, -0.05744282, -0.05777345, 
    -0.05722709, -0.05674197, -0.05613744, -0.05503822, -0.0552909, 
    -0.05438378, -0.06437248, -0.06372607, -0.06378283, -0.06311262, 
    -0.06262136, -0.06156942, -0.05991794, -0.06053387, -0.05940789, 
    -0.05918429, -0.06089685, -0.05983965, -0.06329708, -0.0627255, 
    -0.06306528, -0.0643212, -0.06039126, -0.06237794, -0.05875773, 
    -0.0597981, -0.05681088, -0.05827778, -0.05543046, -0.0542547, 
    -0.0531707, -0.05193007, -0.06337607, -0.06381224, -0.0630334, 
    -0.0619709, -0.06100094, -0.05973412, -0.05960601, -0.059372, 
    -0.05877014, -0.05826864, -0.05929811, -0.05814359, -0.06259346, 
    -0.06022179, -0.06397781, -0.0628233, -0.06203309, -0.06237864, 
    -0.06060469, -0.06019375, -0.05855156, -0.05939502, -0.05454254, 
    -0.05663989, -0.05100461, -0.05252206, -0.0639653, -0.06337761, 
    -0.06137281, -0.06231889, -0.05965052, -0.0590109, -0.05849595, 
    -0.05784388, -0.05777398, -0.05739143, -0.05801958, -0.05741615, 
    -0.05973145, -0.05868579, -0.06159892, -0.06087714, -0.06120819, 
    -0.06157326, -0.06045329, -0.05928174, -0.05925711, -0.05888627, 
    -0.05785311, -0.05963994, -0.05427714, -0.05753061, -0.06274275, 
    -0.06163623, -0.06147993, -0.06190521, -0.05907472, -0.06008543, 
    -0.05740075, -0.05811463, -0.05694946, -0.05752557, -0.0576108, 
    -0.05836016, -0.05883145, -0.06003869, -0.06103876, -0.06184337, 
    -0.06165538, -0.0607747, -0.05921084, -0.05776758, -0.05808076, 
    -0.05703721, -0.05984019, -0.05864882, -0.05910648, -0.05792041, 
    -0.06055029, -0.0583032, -0.06113799, -0.06088421, -0.06010567, 
    -0.05856876, -0.05823416, -0.05787868, -0.05809781, -0.05917168, 
    -0.05934951, -0.06012451, -0.06034014, -0.06093939, -0.06143982, 
    -0.0609824, -0.06050557, -0.05917129, -0.05799333, -0.05673507, 
    -0.05643127, -0.05500184, -0.05616255, -0.0542595, -0.05587307, 
    -0.05310878, -0.05817572, -0.05592152, -0.06007052, -0.05960958, 
    -0.05878441, -0.0569339, -0.05792593, -0.05676747, -0.0593565, 
    -0.06074445, -0.06110886, -0.06179413, -0.06109329, -0.06115, -0.060486, 
    -0.06069862, -0.05912748, -0.05996645, -0.0576129, -0.05677657, 
    -0.05447811, -0.05311397, -0.05175968, -0.05117244, -0.050995, -0.05092099,
  -0.06388779, -0.0621957, -0.06252144, -0.0611801, -0.06192096, -0.06104733, 
    -0.06354145, -0.0621293, -0.06302749, -0.06373385, -0.0586514, 
    -0.06112089, -0.05618334, -0.05768753, -0.05397669, -0.05641495, 
    -0.05349682, -0.05404583, -0.05240908, -0.05287334, -0.0508287, 
    -0.05219606, -0.04979744, -0.05115234, -0.05093816, -0.05224171, 
    -0.0606166, -0.05895376, -0.06071641, -0.06047636, -0.060584, 
    -0.06190551, -0.06258127, -0.06401895, -0.06375575, -0.06270096, 
    -0.0603687, -0.06115149, -0.05919647, -0.05923999, -0.05712903, 
    -0.05807219, -0.05462673, -0.05558663, -0.05285389, -0.0535294, 
    -0.05288542, -0.05307996, -0.05288289, -0.05387678, -0.05344888, 
    -0.05433108, -0.05789445, -0.05682573, -0.06006731, -0.06209637, 
    -0.06347887, -0.06447677, -0.06433482, -0.064065, -0.06269484, 
    -0.06143121, -0.06048382, -0.05985753, -0.05924625, -0.05742997, 
    -0.05648964, -0.0544344, -0.05480034, -0.05418182, -0.05359703, 
    -0.05262791, -0.05278634, -0.05236325, -0.05419815, -0.05297225, 
    -0.05500975, -0.05444551, -0.05908048, -0.06093943, -0.06174508, 
    -0.06245868, -0.06422587, -0.06300065, -0.06348106, -0.06234371, 
    -0.06163064, -0.0619824, -0.05984049, -0.06066504, -0.05643434, 
    -0.05822258, -0.05366495, -0.05472506, -0.05341365, -0.05407925, 
    -0.05294329, -0.05396466, -0.05220662, -0.05183069, -0.05208731, 
    -0.05110795, -0.05402179, -0.05288537, -0.06199226, -0.06193475, 
    -0.06166754, -0.06285001, -0.06292304, -0.06402615, -0.0630438, 
    -0.06262963, -0.06158958, -0.06098172, -0.06040901, -0.05916699, 
    -0.05780731, -0.05595379, -0.05465576, -0.05380101, -0.05432372, 
    -0.053862, -0.05437836, -0.05462195, -0.05197123, -0.05344487, 
    -0.05124778, -0.0513672, -0.05235321, -0.05135374, -0.06189441, 
    -0.06222579, -0.06338874, -0.06247696, -0.06414735, -0.06320731, 
    -0.06267247, -0.06064757, -0.06021089, -0.05980837, -0.05902068, 
    -0.05802357, -0.05631131, -0.05485908, -0.05356321, -0.05365722, 
    -0.0536241, -0.05333808, -0.05404903, -0.05322219, -0.05308449, 
    -0.05344511, -0.05138322, -0.05196481, -0.05136975, -0.05174768, 
    -0.06211791, -0.06156215, -0.06186188, -0.06129931, -0.06169511, 
    -0.05995267, -0.05943906, -0.05708872, -0.05804302, -0.05653113, 
    -0.05788783, -0.05764526, -0.05648219, -0.0578138, -0.05493816, 
    -0.05687295, -0.053327, -0.05520742, -0.0532111, -0.05356875, 
    -0.05297783, -0.05245356, -0.05180076, -0.05061536, -0.05088767, 
    -0.04991059, -0.0607421, -0.06003664, -0.06009855, -0.05936768, 
    -0.05883234, -0.05768722, -0.05589272, -0.05656153, -0.05533935, 
    -0.05509686, -0.05695592, -0.05580776, -0.05956877, -0.0589458, 
    -0.05931608, -0.06068612, -0.05640662, -0.05856723, -0.05463452, 
    -0.05576267, -0.05252801, -0.05411465, -0.05103812, -0.04977168, 
    -0.04860621, -0.04727495, -0.0596549, -0.06013064, -0.05928133, 
    -0.05812408, -0.05706906, -0.05569324, -0.05555425, -0.05530042, 
    -0.05464797, -0.05410476, -0.05522029, -0.05396936, -0.05880197, 
    -0.05622259, -0.0603113, -0.05905237, -0.05819177, -0.05856798, 
    -0.05663845, -0.05619214, -0.05441116, -0.05532538, -0.0500815, 
    -0.05234328, -0.04628376, -0.04790984, -0.06029765, -0.05965658, 
    -0.05747337, -0.05850292, -0.05560254, -0.0549089, -0.05435092, 
    -0.05364497, -0.05356933, -0.05315553, -0.05383512, -0.05318226, 
    -0.05569034, -0.05455658, -0.05771931, -0.05693449, -0.05729436, 
    -0.0576914, -0.05647399, -0.05520254, -0.05517583, -0.05477382, 
    -0.05365496, -0.05559106, -0.04979583, -0.05330605, -0.0589646, 
    -0.0577599, -0.05758987, -0.05805258, -0.05497808, -0.05607454, 
    -0.0531656, -0.053938, -0.05267774, -0.0533006, -0.05339279, -0.05420386, 
    -0.0547144, -0.0560238, -0.05711016, -0.05798528, -0.05778073, 
    -0.05682317, -0.05512566, -0.05356241, -0.05390134, -0.05277258, 
    -0.05580835, -0.05451653, -0.05501251, -0.05372779, -0.05657936, 
    -0.05414217, -0.05721804, -0.05694218, -0.05609651, -0.05442979, 
    -0.05406742, -0.05368262, -0.0539198, -0.0550832, -0.05527603, 
    -0.05611696, -0.0563511, -0.05700215, -0.05754625, -0.0570489, 
    -0.05653077, -0.05508277, -0.0538067, -0.0524461, -0.05211798, 
    -0.05057617, -0.05182787, -0.04977684, -0.05151549, -0.0485397, 
    -0.05400415, -0.05156776, -0.05605835, -0.05555812, -0.05466343, 
    -0.05266093, -0.05373377, -0.0524811, -0.05528361, -0.05679031, 
    -0.05718638, -0.0579317, -0.05716944, -0.0572311, -0.05650952, 
    -0.05674051, -0.05503528, -0.05594538, -0.05339506, -0.05249093, 
    -0.05001213, -0.04854528, -0.04709234, -0.04646338, -0.04627346, 
    -0.04619427,
  -0.04035017, -0.03907184, -0.03931778, -0.03830553, -0.03886447, 
    -0.0382054, -0.04008836, -0.03902173, -0.03969999, -0.0402338, 
    -0.03640078, -0.03826088, -0.03454657, -0.03567605, -0.0328932, 
    -0.03472036, -0.03253425, -0.03294493, -0.03172141, -0.03206819, 
    -0.03054259, -0.03156237, -0.02977479, -0.03078379, -0.03062415, 
    -0.03159644, -0.03788066, -0.03662828, -0.0379559, -0.03777496, 
    -0.03785609, -0.03885281, -0.03936297, -0.04044933, -0.04025035, 
    -0.03945336, -0.03769382, -0.03828395, -0.03681095, -0.03684371, 
    -0.03525646, -0.03596519, -0.0333798, -0.03409905, -0.03205366, 
    -0.03255861, -0.03207722, -0.0322226, -0.03207533, -0.03281844, 
    -0.0324984, -0.03315843, -0.03583157, -0.0350287, -0.03746673, 
    -0.03899687, -0.04004107, -0.04079557, -0.04068821, -0.04048416, 
    -0.03944873, -0.03849493, -0.03778059, -0.03730871, -0.03684842, 
    -0.03548251, -0.03477641, -0.03323578, -0.03350982, -0.03304671, 
    -0.03260919, -0.03188484, -0.03200319, -0.03168719, -0.03305893, 
    -0.03214211, -0.03366669, -0.0332441, -0.03672365, -0.03812404, 
    -0.03873174, -0.03927039, -0.04060581, -0.03967972, -0.04004272, 
    -0.03918359, -0.03864539, -0.03891084, -0.03729587, -0.03791717, 
    -0.03473491, -0.03607827, -0.03265998, -0.03345343, -0.03247205, 
    -0.03296995, -0.03212046, -0.0328842, -0.03157025, -0.03128969, 
    -0.03148119, -0.0307507, -0.03292694, -0.03207718, -0.03891828, 
    -0.03887488, -0.03867324, -0.03956592, -0.0396211, -0.04045478, 
    -0.03971232, -0.03939948, -0.03861441, -0.03815593, -0.0377242, 
    -0.03678877, -0.03576607, -0.03437437, -0.03340153, -0.03276176, 
    -0.03315292, -0.03280739, -0.03319383, -0.03337621, -0.03139455, 
    -0.0324954, -0.03085493, -0.03094397, -0.03167969, -0.03093393, 
    -0.03884443, -0.03909456, -0.03997295, -0.03928419, -0.04054642, 
    -0.03983586, -0.03943183, -0.03790401, -0.03757491, -0.03727167, 
    -0.03667865, -0.03592864, -0.03464259, -0.03355382, -0.03258389, 
    -0.0326542, -0.03262943, -0.03241555, -0.03294734, -0.03232891, 
    -0.03222599, -0.03249558, -0.03095591, -0.03138977, -0.03094587, 
    -0.03122775, -0.03901312, -0.03859372, -0.03881989, -0.03839545, 
    -0.03869404, -0.03738037, -0.03699357, -0.03522618, -0.03594326, 
    -0.03480755, -0.03582659, -0.03564429, -0.03477082, -0.03577095, 
    -0.03361305, -0.03506416, -0.03240726, -0.0338148, -0.03232063, 
    -0.03258804, -0.03214628, -0.03175462, -0.03126735, -0.03038366, 
    -0.03058653, -0.02985898, -0.03797527, -0.03744362, -0.03749027, 
    -0.03693983, -0.03653692, -0.03567581, -0.03432857, -0.03483037, 
    -0.03391368, -0.03373196, -0.03512646, -0.03426485, -0.03709124, 
    -0.0366223, -0.03690099, -0.03793306, -0.03471411, -0.03633747, 
    -0.03338563, -0.03423104, -0.03181022, -0.03299643, -0.03069865, 
    -0.02975563, -0.0288894, -0.02790193, -0.03715609, -0.03751444, 
    -0.03687483, -0.0360042, -0.03521141, -0.03417898, -0.03407476, 
    -0.0338845, -0.0333957, -0.03298903, -0.03382445, -0.03288772, 
    -0.03651407, -0.03457602, -0.03765057, -0.0367025, -0.0360551, 
    -0.03633804, -0.03488811, -0.03455317, -0.03321838, -0.03390321, 
    -0.02998617, -0.03167228, -0.02716813, -0.02837259, -0.03764028, 
    -0.03715736, -0.03551513, -0.0362891, -0.03411097, -0.03359114, 
    -0.03317328, -0.03264504, -0.03258847, -0.03227909, -0.03278728, 
    -0.03229907, -0.03417681, -0.03332726, -0.03569993, -0.03511037, 
    -0.03538064, -0.03567896, -0.03476467, -0.03381114, -0.03379113, 
    -0.03348995, -0.03265251, -0.03410236, -0.0297736, -0.03239161, 
    -0.03663645, -0.03573044, -0.03560267, -0.03595044, -0.03364296, 
    -0.03446495, -0.03228661, -0.03286425, -0.03192206, -0.03238753, 
    -0.03245645, -0.0330632, -0.03344545, -0.03442689, -0.03524229, 
    -0.03589985, -0.03574609, -0.03502678, -0.03375353, -0.03258329, 
    -0.03283682, -0.03199291, -0.03426529, -0.03329727, -0.03366876, 
    -0.03270698, -0.03484375, -0.03301704, -0.03532331, -0.03511614, 
    -0.03448142, -0.03323233, -0.03296109, -0.0326732, -0.03285063, 
    -0.03372172, -0.03386622, -0.03449677, -0.03467244, -0.03516117, 
    -0.03556988, -0.03519628, -0.03480728, -0.0337214, -0.03276602, 
    -0.03174906, -0.03150408, -0.03035447, -0.03128758, -0.02975948, 
    -0.03105455, -0.02884002, -0.03291374, -0.03109353, -0.0344528, 
    -0.03407767, -0.03340728, -0.03190951, -0.03271146, -0.0317752, 
    -0.0338719, -0.0350021, -0.03529953, -0.03585957, -0.03528681, 
    -0.03533312, -0.03479134, -0.03496472, -0.03368582, -0.03436807, 
    -0.03245816, -0.03178253, -0.02993454, -0.02884416, -0.02776664, 
    -0.02730101, -0.02716052, -0.02710195,
  -0.01970495, -0.01870051, -0.01889313, -0.01810233, -0.01853834, 
    -0.01802441, -0.01949858, -0.0186613, -0.01919307, -0.01961318, 
    -0.01662921, -0.01806758, -0.01521542, -0.01607413, -0.01397334, 
    -0.01534703, -0.01370616, -0.01401192, -0.01310461, -0.01336065, 
    -0.01224113, -0.01298748, -0.01168475, -0.01241691, -0.01230052, 
    -0.01301256, -0.01777202, -0.01680408, -0.01783044, -0.01768999, 
    -0.01775294, -0.01852923, -0.01892854, -0.0197832, -0.01962623, 
    -0.01899943, -0.01762706, -0.01808554, -0.01694472, -0.01696996, 
    -0.0157542, -0.01629521, -0.01433697, -0.01487742, -0.01334991, 
    -0.01372426, -0.01336733, -0.01347495, -0.01336593, -0.01391762, 
    -0.01367953, -0.01417134, -0.01619298, -0.015581, -0.01745114, 
    -0.01864185, -0.01946134, -0.02005678, -0.01997189, -0.01981069, 
    -0.0189958, -0.0182499, -0.01769435, -0.01732889, -0.01697359, 
    -0.01592643, -0.01538952, -0.01422918, -0.01443441, -0.01408788, 
    -0.01376187, -0.01322516, -0.01331259, -0.01307939, -0.01409701, 
    -0.01341534, -0.01455213, -0.0142354, -0.01687748, -0.01796112, 
    -0.01843466, -0.01885599, -0.01990677, -0.01917714, -0.01946264, 
    -0.01878799, -0.01836725, -0.01857458, -0.01731896, -0.01780037, 
    -0.01535806, -0.0163818, -0.01379965, -0.01439214, -0.01365996, 
    -0.01403058, -0.01339933, -0.01396663, -0.01299328, -0.01278711, 
    -0.01292777, -0.01239277, -0.0139985, -0.0133673, -0.0185804, 
    -0.01854647, -0.01838898, -0.01908777, -0.01913109, -0.0197875, 
    -0.01920275, -0.01895718, -0.01834308, -0.01798592, -0.01765062, 
    -0.01692763, -0.01614291, -0.01508521, -0.01435325, -0.0138754, 
    -0.01416722, -0.01390938, -0.0141978, -0.01433429, -0.0128641, 
    -0.0136773, -0.01246885, -0.01253391, -0.01307387, -0.01252657, 
    -0.01852268, -0.01871829, -0.01940772, -0.0188668, -0.01985986, 
    -0.01929986, -0.01898255, -0.01779014, -0.01753491, -0.01730026, 
    -0.01684284, -0.01626723, -0.01528811, -0.01446741, -0.01374306, 
    -0.01379535, -0.01377692, -0.01361802, -0.01401371, -0.01355374, 
    -0.01347746, -0.01367744, -0.01254264, -0.01286059, -0.0125353, 
    -0.01274168, -0.01865457, -0.01832693, -0.0185035, -0.01817236, 
    -0.01840522, -0.01738431, -0.01708551, -0.01573116, -0.01627842, 
    -0.01541313, -0.01618917, -0.01604987, -0.01538528, -0.01614663, 
    -0.01451186, -0.01560794, -0.01361187, -0.01466342, -0.0135476, 
    -0.01374614, -0.01341843, -0.01312909, -0.01277073, -0.01212556, 
    -0.01227312, -0.01174552, -0.01784549, -0.01743325, -0.01746936, 
    -0.01704405, -0.01673382, -0.01607395, -0.01505061, -0.01543043, 
    -0.0147378, -0.01460116, -0.0156553, -0.0150025, -0.01716087, 
    -0.01679948, -0.0170141, -0.0178127, -0.01534229, -0.01658059, 
    -0.01434134, -0.01497698, -0.0131701, -0.01405035, -0.01235481, 
    -0.01167093, -0.01104941, -0.0103492, -0.01721095, -0.01748808, 
    -0.01699394, -0.01632508, -0.01571992, -0.0149377, -0.01485912, 
    -0.01471585, -0.01434888, -0.01404482, -0.01467068, -0.01396925, 
    -0.01671625, -0.01523771, -0.01759354, -0.01686119, -0.01636406, 
    -0.01658102, -0.01547424, -0.01522042, -0.01421617, -0.01472993, 
    -0.01183743, -0.0130684, -0.009834953, -0.01068181, -0.01758556, 
    -0.01721193, -0.0159513, -0.01654346, -0.01488641, -0.01449541, 
    -0.01418244, -0.01378853, -0.01374646, -0.0135168, -0.01389441, 
    -0.01353161, -0.01493606, -0.01429764, -0.01609237, -0.01564306, 
    -0.01584878, -0.01607635, -0.01538061, -0.01466068, -0.01464562, 
    -0.01441952, -0.01379409, -0.01487992, -0.01168389, -0.01360025, 
    -0.01681037, -0.01611568, -0.0160181, -0.01628392, -0.01453431, 
    -0.01515368, -0.01352238, -0.01395176, -0.01325265, -0.01359722, 
    -0.01364838, -0.0141002, -0.01438616, -0.0151249, -0.01574342, 
    -0.01624521, -0.01612764, -0.01557954, -0.01461737, -0.01374261, 
    -0.01393131, -0.01330499, -0.01500283, -0.01427519, -0.01455368, 
    -0.01383462, -0.01544059, -0.01406572, -0.01580511, -0.01564746, 
    -0.01516614, -0.0142266, -0.01402398, -0.01380948, -0.01394161, 
    -0.01459346, -0.0147021, -0.01517775, -0.01531073, -0.0156817, 
    -0.01599308, -0.01570841, -0.01541293, -0.01459322, -0.01387857, 
    -0.01312499, -0.0129446, -0.01210436, -0.01278557, -0.0116737, 
    -0.0126148, -0.01101418, -0.01398866, -0.01264334, -0.0151445, 
    -0.01486131, -0.01435756, -0.01324338, -0.01383795, -0.01314426, 
    -0.01470637, -0.01556079, -0.01578699, -0.0162144, -0.01577731, 
    -0.01581258, -0.01540083, -0.0155324, -0.01456649, -0.01508045, 
    -0.01364964, -0.01314967, -0.01180011, -0.01101713, -0.01025399, 
    -0.009927681, -0.009829647, -0.009788836,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  365.4042, 367.2402, 366.8827, 368.3649, 367.543, 368.5133, 365.7758, 
    367.3133, 366.3313, 365.5691, 371.2495, 368.431, 374.1903, 372.3824, 
    376.9343, 373.9088, 377.5461, 376.8464, 378.954, 378.3494, 381.0539, 
    379.2332, 382.46, 380.6184, 380.9062, 379.1733, 368.9968, 370.8979, 
    368.8844, 369.1551, 369.0335, 367.5601, 366.8174, 365.2639, 365.5456, 
    366.6866, 369.2768, 368.3968, 370.6167, 370.5664, 373.0479, 371.9277, 
    376.1141, 374.9211, 378.3746, 377.5043, 378.3338, 378.0821, 378.3371, 
    377.0611, 377.6075, 376.4858, 372.1374, 373.4122, 369.6187, 367.3497, 
    365.8432, 364.7769, 364.9275, 365.2148, 366.6933, 368.0851, 369.1465, 
    369.8577, 370.5592, 372.6887, 373.8182, 376.3557, 375.8967, 376.6743, 
    377.4178, 378.6684, 378.4623, 379.014, 376.6536, 378.2214, 375.6355, 
    376.3417, 370.7512, 368.634, 367.7374, 366.9514, 365.0434, 366.3604, 
    365.8409, 367.0775, 367.8638, 367.4752, 369.8771, 368.9422, 373.8852, 
    371.7509, 377.331, 375.9909, 377.6526, 376.804, 378.2589, 376.9494, 
    379.2194, 379.7149, 379.3763, 380.6779, 376.8769, 378.3339, 367.4643, 
    367.5278, 367.823, 366.5242, 366.4447, 365.2563, 366.3135, 366.7645, 
    367.9093, 368.5866, 369.2311, 370.6508, 372.2405, 374.4705, 376.0777, 
    377.1575, 376.4951, 377.0798, 376.4262, 376.12, 379.5293, 377.6126, 
    380.4905, 380.3308, 379.0272, 380.3488, 367.5723, 367.207, 365.9404, 
    366.9314, 365.127, 366.1364, 366.7177, 368.962, 369.4555, 369.9139, 
    370.82, 371.985, 374.0345, 375.8234, 377.461, 377.3409, 377.3831, 
    377.7497, 376.8423, 377.8987, 378.0763, 377.6123, 380.3094, 379.5377, 
    380.3274, 379.8247, 367.3257, 367.9398, 367.6082, 368.2319, 367.7925, 
    369.7493, 370.3373, 373.0963, 371.9621, 373.7679, 372.1452, 372.4325, 
    373.8274, 372.2327, 375.7249, 373.3555, 377.7639, 375.3901, 377.913, 
    377.4539, 378.2141, 378.8959, 379.7545, 381.3423, 380.9742, 382.3042, 
    368.8555, 369.6536, 369.5831, 370.4193, 371.0385, 372.3827, 374.5452, 
    373.731, 375.2264, 375.5272, 373.2555, 374.6494, 370.1882, 370.9069, 
    370.4788, 368.9185, 373.9188, 371.3474, 376.1043, 374.7047, 378.7986, 
    376.7594, 380.7717, 382.4956, 384.1092, 386.001, 370.0894, 369.5466, 
    370.5187, 371.8668, 373.1198, 374.79, 374.961, 375.2746, 376.0874, 
    376.7718, 375.374, 376.9434, 371.0741, 374.1425, 369.3417, 370.7834, 
    371.7871, 371.3464, 373.638, 374.1794, 376.385, 375.2437, 382.0699, 
    379.0403, 387.4445, 385.0922, 369.3571, 370.0875, 372.6368, 371.4224, 
    374.9016, 375.7612, 376.4608, 377.3566, 377.4532, 377.9846, 377.114, 
    377.9501, 374.7935, 376.2021, 372.3446, 373.2813, 372.8501, 372.3777, 
    373.837, 375.3961, 375.4291, 375.9299, 377.3443, 374.9157, 382.4627, 
    377.7913, 370.8849, 372.2967, 372.4982, 371.9508, 375.675, 374.3229, 
    377.9716, 376.9832, 378.6035, 377.7978, 377.6794, 376.6464, 376.0042, 
    374.3849, 373.0705, 372.0301, 372.2719, 373.4152, 375.4915, 377.4621, 
    377.0299, 378.4802, 374.6486, 376.2524, 375.6321, 377.2508, 373.7095, 
    376.7249, 372.9413, 373.272, 374.2961, 376.3616, 376.819, 377.3085, 
    377.0063, 375.5442, 375.3048, 374.2711, 373.9861, 373.2, 372.55, 
    373.1439, 373.7683, 375.5447, 377.1503, 378.9056, 379.3358, 381.3956, 
    379.7188, 382.4889, 380.1338, 384.2029, 376.8995, 380.0639, 374.3426, 
    374.9563, 376.0682, 378.6255, 377.2432, 378.86, 375.2954, 373.4549, 
    372.9792, 372.0934, 372.9995, 372.9257, 373.7939, 373.5148, 375.6038, 
    374.4807, 377.6765, 378.8471, 382.1648, 384.1948, 386.2644, 387.1805, 
    387.4596, 387.5764 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.195739e-08, 6.223058e-08, 6.217748e-08, 6.239782e-08, 6.22756e-08, 
    6.241988e-08, 6.201279e-08, 6.224143e-08, 6.209547e-08, 6.198199e-08, 
    6.282544e-08, 6.240766e-08, 6.325951e-08, 6.299303e-08, 6.36625e-08, 
    6.321804e-08, 6.375213e-08, 6.364969e-08, 6.395803e-08, 6.38697e-08, 
    6.426407e-08, 6.39988e-08, 6.446854e-08, 6.420073e-08, 6.424262e-08, 
    6.399005e-08, 6.249174e-08, 6.277342e-08, 6.247505e-08, 6.251522e-08, 
    6.24972e-08, 6.227812e-08, 6.216771e-08, 6.193653e-08, 6.19785e-08, 
    6.21483e-08, 6.253328e-08, 6.240261e-08, 6.273198e-08, 6.272454e-08, 
    6.309124e-08, 6.29259e-08, 6.354229e-08, 6.33671e-08, 6.387339e-08, 
    6.374605e-08, 6.38674e-08, 6.38306e-08, 6.386788e-08, 6.368114e-08, 
    6.376114e-08, 6.359683e-08, 6.295686e-08, 6.314493e-08, 6.258403e-08, 
    6.224678e-08, 6.202281e-08, 6.186388e-08, 6.188635e-08, 6.192918e-08, 
    6.21493e-08, 6.235626e-08, 6.2514e-08, 6.261951e-08, 6.272347e-08, 
    6.303814e-08, 6.320472e-08, 6.357771e-08, 6.351041e-08, 6.362443e-08, 
    6.373339e-08, 6.39163e-08, 6.388619e-08, 6.396677e-08, 6.362144e-08, 
    6.385094e-08, 6.347207e-08, 6.357569e-08, 6.275169e-08, 6.243786e-08, 
    6.230444e-08, 6.218769e-08, 6.190362e-08, 6.209979e-08, 6.202245e-08, 
    6.220644e-08, 6.232334e-08, 6.226553e-08, 6.262239e-08, 6.248365e-08, 
    6.321459e-08, 6.289974e-08, 6.372068e-08, 6.352423e-08, 6.376777e-08, 
    6.36435e-08, 6.385643e-08, 6.366479e-08, 6.399677e-08, 6.406906e-08, 
    6.401966e-08, 6.420943e-08, 6.365416e-08, 6.38674e-08, 6.226391e-08, 
    6.227334e-08, 6.231727e-08, 6.212414e-08, 6.211233e-08, 6.193537e-08, 
    6.209284e-08, 6.215989e-08, 6.233013e-08, 6.243081e-08, 6.252654e-08, 
    6.273701e-08, 6.297206e-08, 6.330077e-08, 6.353696e-08, 6.369527e-08, 
    6.35982e-08, 6.368391e-08, 6.35881e-08, 6.354319e-08, 6.404196e-08, 
    6.376189e-08, 6.418213e-08, 6.415888e-08, 6.396869e-08, 6.41615e-08, 
    6.227996e-08, 6.222569e-08, 6.203729e-08, 6.218473e-08, 6.19161e-08, 
    6.206646e-08, 6.215291e-08, 6.248654e-08, 6.255986e-08, 6.262782e-08, 
    6.276207e-08, 6.293436e-08, 6.323661e-08, 6.349962e-08, 6.373973e-08, 
    6.372213e-08, 6.372833e-08, 6.378196e-08, 6.36491e-08, 6.380377e-08, 
    6.382973e-08, 6.376186e-08, 6.415576e-08, 6.404323e-08, 6.415839e-08, 
    6.408511e-08, 6.224334e-08, 6.233464e-08, 6.22853e-08, 6.237808e-08, 
    6.231271e-08, 6.260337e-08, 6.269052e-08, 6.309833e-08, 6.293097e-08, 
    6.319734e-08, 6.295803e-08, 6.300043e-08, 6.320601e-08, 6.297097e-08, 
    6.348511e-08, 6.313651e-08, 6.378404e-08, 6.343591e-08, 6.380586e-08, 
    6.373869e-08, 6.384992e-08, 6.394953e-08, 6.407485e-08, 6.43061e-08, 
    6.425255e-08, 6.444595e-08, 6.247078e-08, 6.25892e-08, 6.257878e-08, 
    6.270273e-08, 6.27944e-08, 6.29931e-08, 6.331179e-08, 6.319195e-08, 
    6.341197e-08, 6.345614e-08, 6.312188e-08, 6.33271e-08, 6.266848e-08, 
    6.277487e-08, 6.271153e-08, 6.248011e-08, 6.321955e-08, 6.284005e-08, 
    6.354086e-08, 6.333526e-08, 6.393532e-08, 6.363688e-08, 6.422307e-08, 
    6.447366e-08, 6.470955e-08, 6.498519e-08, 6.265385e-08, 6.257338e-08, 
    6.271748e-08, 6.291684e-08, 6.310184e-08, 6.33478e-08, 6.337297e-08, 
    6.341904e-08, 6.35384e-08, 6.363876e-08, 6.34336e-08, 6.366392e-08, 
    6.279953e-08, 6.32525e-08, 6.254295e-08, 6.275658e-08, 6.290509e-08, 
    6.283995e-08, 6.317826e-08, 6.325799e-08, 6.358201e-08, 6.341452e-08, 
    6.44118e-08, 6.397055e-08, 6.51951e-08, 6.485286e-08, 6.254526e-08, 
    6.265358e-08, 6.303058e-08, 6.28512e-08, 6.336422e-08, 6.34905e-08, 
    6.359317e-08, 6.37244e-08, 6.373858e-08, 6.381633e-08, 6.368892e-08, 
    6.38113e-08, 6.334832e-08, 6.355521e-08, 6.298749e-08, 6.312566e-08, 
    6.30621e-08, 6.299238e-08, 6.320757e-08, 6.343683e-08, 6.344175e-08, 
    6.351525e-08, 6.372239e-08, 6.33663e-08, 6.446873e-08, 6.378785e-08, 
    6.27717e-08, 6.298033e-08, 6.301015e-08, 6.292932e-08, 6.347784e-08, 
    6.327909e-08, 6.381444e-08, 6.366975e-08, 6.390682e-08, 6.378902e-08, 
    6.377169e-08, 6.362038e-08, 6.352618e-08, 6.32882e-08, 6.309457e-08, 
    6.294105e-08, 6.297675e-08, 6.314539e-08, 6.345086e-08, 6.373985e-08, 
    6.367654e-08, 6.388881e-08, 6.332702e-08, 6.356257e-08, 6.347153e-08, 
    6.370894e-08, 6.318876e-08, 6.363167e-08, 6.307555e-08, 6.312431e-08, 
    6.327515e-08, 6.357854e-08, 6.364569e-08, 6.371736e-08, 6.367314e-08, 
    6.345861e-08, 6.342348e-08, 6.327148e-08, 6.322951e-08, 6.31137e-08, 
    6.301781e-08, 6.310542e-08, 6.319741e-08, 6.345871e-08, 6.369419e-08, 
    6.395094e-08, 6.401378e-08, 6.431375e-08, 6.406955e-08, 6.447252e-08, 
    6.412989e-08, 6.472303e-08, 6.365737e-08, 6.411983e-08, 6.328201e-08, 
    6.337227e-08, 6.353551e-08, 6.390996e-08, 6.370782e-08, 6.394423e-08, 
    6.34221e-08, 6.315121e-08, 6.308114e-08, 6.295038e-08, 6.308413e-08, 
    6.307325e-08, 6.320123e-08, 6.316011e-08, 6.346739e-08, 6.330233e-08, 
    6.377125e-08, 6.394237e-08, 6.442568e-08, 6.472197e-08, 6.502361e-08, 
    6.515678e-08, 6.519732e-08, 6.521426e-08 ;

 SOM_C_LEACHED =
  4.936022e-21, 4.1143e-20, 4.041273e-20, 1.724337e-20, 5.857769e-20, 
    -9.818658e-20, 1.260552e-20, -8.411525e-21, -7.421965e-20, 3.192002e-20, 
    3.089081e-20, 6.664967e-22, 3.764863e-20, -2.756924e-20, 5.182015e-20, 
    6.319044e-21, -4.87961e-20, 2.227307e-20, 6.496721e-21, 6.283585e-20, 
    -5.986705e-20, 2.893463e-22, 7.045066e-20, 7.163681e-20, 2.268712e-20, 
    2.34715e-20, -1.948031e-20, -1.86402e-21, 1.244342e-20, -2.160986e-20, 
    -5.158285e-20, 1.51006e-20, -2.175008e-20, 5.761332e-21, -2.239059e-21, 
    -4.726187e-20, -3.080681e-20, 2.042081e-20, -1.00094e-20, 7.512718e-21, 
    -2.726049e-20, 5.393755e-20, 1.569108e-20, 5.903489e-21, -8.053157e-21, 
    -5.620685e-20, -2.79531e-20, 4.141649e-20, -1.185704e-20, -1.532275e-20, 
    3.369727e-21, 1.829032e-20, 5.394022e-20, 1.032682e-20, 4.35798e-20, 
    -2.613179e-20, -1.360893e-20, -2.007421e-21, -1.166803e-20, 3.194618e-20, 
    -1.458973e-20, -3.522284e-20, -6.150691e-20, -2.598597e-20, 3.242856e-20, 
    5.271661e-20, -4.806081e-20, 4.616914e-20, -6.050366e-20, 1.596313e-20, 
    -1.479888e-21, 3.342885e-20, 8.066896e-21, -1.022811e-20, 5.310882e-21, 
    -6.101345e-20, 4.432733e-20, 6.915926e-20, -3.074092e-20, 5.775661e-20, 
    2.194357e-20, 1.721979e-20, -2.114508e-21, -1.836131e-20, 6.871203e-20, 
    4.082698e-20, -3.370014e-20, -2.039437e-20, 4.787554e-20, 4.00391e-21, 
    -8.90438e-21, 7.301519e-20, 4.308223e-20, -4.928739e-20, 5.026662e-20, 
    4.52041e-20, -5.045248e-20, -2.590601e-20, 2.439756e-21, 3.049714e-20, 
    -1.703082e-20, -3.453504e-20, -3.866252e-20, -1.623826e-20, 1.780795e-20, 
    5.572143e-20, 1.599129e-20, -1.096841e-20, 8.054167e-21, 1.032612e-20, 
    4.393568e-20, 2.018816e-20, 8.220296e-21, 2.872957e-21, -2.036067e-20, 
    -7.195225e-20, 8.932931e-21, 4.738013e-20, -2.147204e-20, 6.912473e-21, 
    -4.932925e-20, 5.823491e-21, -7.962205e-21, -3.540523e-20, -2.016731e-20, 
    3.601378e-21, 1.739535e-20, 3.003485e-20, -1.942525e-20, -1.359487e-20, 
    -7.606421e-20, 6.008606e-20, -7.865649e-20, -1.918209e-20, -2.153492e-21, 
    2.591715e-20, 5.713385e-21, -1.51939e-20, -6.9144e-20, -1.755212e-20, 
    4.707441e-20, -7.406931e-20, 4.389548e-21, -2.220484e-20, 2.995039e-20, 
    -2.617486e-20, 1.984529e-20, -3.018379e-20, 1.609011e-20, 1.178868e-20, 
    3.703619e-20, 1.396621e-20, -1.229911e-20, -2.600728e-20, 2.557692e-20, 
    3.768063e-20, 7.2552e-21, 5.901804e-20, -2.174714e-20, -1.966715e-20, 
    7.186326e-21, -1.93271e-20, -3.658474e-20, -7.339851e-20, -8.835773e-21, 
    -5.84002e-22, 4.365369e-20, 3.546331e-20, 1.110534e-20, -6.352029e-20, 
    -2.990431e-20, 9.297429e-21, 5.231636e-20, -5.788125e-20, -6.339914e-20, 
    1.688907e-20, -1.252197e-20, -1.656602e-20, -4.981973e-20, 2.868155e-20, 
    2.593004e-20, -1.072038e-20, 1.308235e-20, -1.994897e-20, 2.985635e-20, 
    -1.93161e-20, 2.398089e-20, -1.340709e-20, -7.56551e-21, 6.245498e-21, 
    5.477421e-20, 2.641034e-20, 5.825902e-20, 8.48525e-20, -2.128646e-21, 
    -1.427208e-21, -5.471941e-21, 2.278079e-20, 5.573683e-20, -1.535009e-20, 
    2.727595e-20, -2.0704e-20, 3.866939e-20, -1.762106e-20, -6.437288e-21, 
    7.130648e-21, 3.886405e-20, 3.178412e-20, -6.021011e-20, -1.365408e-20, 
    5.882012e-20, -7.948039e-20, 9.354384e-21, 5.148082e-20, -2.038714e-21, 
    8.018991e-20, 2.365529e-20, 3.029312e-20, 8.58454e-20, 2.888958e-20, 
    4.255222e-20, -5.549672e-20, -9.281552e-21, -4.719338e-21, 4.105127e-20, 
    1.148445e-20, -1.090389e-20, -8.551764e-22, 3.595354e-20, 3.109447e-20, 
    -6.904247e-20, 4.249718e-20, 3.303014e-20, 4.057555e-20, 1.175251e-20, 
    -2.612678e-20, 3.29934e-20, 1.824175e-20, -1.93711e-20, -3.646712e-20, 
    3.858886e-20, 1.965875e-20, 1.512953e-20, 5.968859e-21, 2.382168e-20, 
    -3.238044e-20, -5.28958e-21, -2.506083e-20, -2.068301e-20, 2.454346e-22, 
    -5.530857e-20, -8.636876e-21, 3.016687e-20, 5.223514e-20, 3.378449e-20, 
    -7.988966e-20, 1.146258e-20, -2.207504e-20, -5.003001e-20, 3.962294e-20, 
    -5.445707e-20, 8.315752e-21, -5.560796e-20, 1.226091e-20, -1.464468e-21, 
    -1.466811e-20, -1.939512e-20, -6.025069e-20, 1.108805e-20, -1.820541e-21, 
    1.495962e-20, 1.896723e-20, -3.587005e-20, 6.785333e-20, -4.517911e-20, 
    -3.59591e-20, 4.58524e-21, -1.232457e-21, -1.404046e-20, 2.150462e-20, 
    8.870867e-20, 1.400404e-21, -2.658322e-21, -4.073259e-20, 3.70481e-20, 
    -3.830821e-20, -9.87815e-20, -5.510503e-20, 2.88352e-20, -1.368548e-20, 
    4.335473e-21, -3.944456e-20, 2.279656e-20, 4.391462e-20, -2.935374e-20, 
    -2.876125e-21, -3.438794e-20, -5.356528e-20, 1.420026e-20, -3.244247e-20, 
    1.652792e-20, -2.215282e-20, -9.801052e-21, -1.868588e-20, -3.886962e-20, 
    2.259528e-20, -1.226247e-20, -4.589298e-20, 3.536982e-20, -1.325736e-20, 
    -1.626931e-20, -1.162202e-21, -5.046714e-21, 1.703564e-20, -6.847972e-20, 
    4.101231e-20, -3.484779e-20, -1.752131e-20, 2.364135e-20, -8.127667e-20, 
    2.094305e-20, -3.293405e-20, 1.100529e-20, 7.334848e-20, 3.911678e-20, 
    -1.156062e-21, 3.679084e-20, -9.708978e-20, -1.118218e-20, -3.348546e-20, 
    4.027695e-20, 8.112065e-20, 1.200472e-20, 2.465105e-20, -5.844556e-20, 
    5.75043e-20, -3.564532e-20, -1.891769e-20 ;

 SR =
  6.195836e-08, 6.223155e-08, 6.217844e-08, 6.23988e-08, 6.227657e-08, 
    6.242085e-08, 6.201375e-08, 6.224239e-08, 6.209643e-08, 6.198296e-08, 
    6.282642e-08, 6.240863e-08, 6.326049e-08, 6.2994e-08, 6.366348e-08, 
    6.321901e-08, 6.375311e-08, 6.365067e-08, 6.395901e-08, 6.387068e-08, 
    6.426506e-08, 6.399979e-08, 6.446953e-08, 6.420172e-08, 6.424361e-08, 
    6.399104e-08, 6.249272e-08, 6.27744e-08, 6.247603e-08, 6.251619e-08, 
    6.249817e-08, 6.227909e-08, 6.216867e-08, 6.193749e-08, 6.197946e-08, 
    6.214927e-08, 6.253426e-08, 6.240357e-08, 6.273295e-08, 6.272551e-08, 
    6.309222e-08, 6.292688e-08, 6.354328e-08, 6.336808e-08, 6.387437e-08, 
    6.374704e-08, 6.386838e-08, 6.383159e-08, 6.386886e-08, 6.368212e-08, 
    6.376213e-08, 6.359781e-08, 6.295784e-08, 6.314591e-08, 6.2585e-08, 
    6.224774e-08, 6.202378e-08, 6.186485e-08, 6.188731e-08, 6.193014e-08, 
    6.215026e-08, 6.235724e-08, 6.251497e-08, 6.262048e-08, 6.272445e-08, 
    6.303911e-08, 6.32057e-08, 6.357869e-08, 6.351139e-08, 6.362541e-08, 
    6.373437e-08, 6.391728e-08, 6.388717e-08, 6.396776e-08, 6.362242e-08, 
    6.385192e-08, 6.347305e-08, 6.357667e-08, 6.275266e-08, 6.243883e-08, 
    6.23054e-08, 6.218865e-08, 6.190459e-08, 6.210075e-08, 6.202342e-08, 
    6.220741e-08, 6.232432e-08, 6.22665e-08, 6.262336e-08, 6.248462e-08, 
    6.321557e-08, 6.290072e-08, 6.372166e-08, 6.352521e-08, 6.376875e-08, 
    6.364448e-08, 6.385741e-08, 6.366577e-08, 6.399775e-08, 6.407004e-08, 
    6.402064e-08, 6.421042e-08, 6.365515e-08, 6.386838e-08, 6.226487e-08, 
    6.22743e-08, 6.231824e-08, 6.212511e-08, 6.21133e-08, 6.193633e-08, 
    6.20938e-08, 6.216086e-08, 6.23311e-08, 6.243179e-08, 6.252751e-08, 
    6.273797e-08, 6.297304e-08, 6.330175e-08, 6.353794e-08, 6.369626e-08, 
    6.359918e-08, 6.368489e-08, 6.358908e-08, 6.354417e-08, 6.404295e-08, 
    6.376287e-08, 6.418312e-08, 6.415987e-08, 6.396967e-08, 6.416249e-08, 
    6.228093e-08, 6.222666e-08, 6.203825e-08, 6.21857e-08, 6.191706e-08, 
    6.206743e-08, 6.215388e-08, 6.248751e-08, 6.256082e-08, 6.262879e-08, 
    6.276304e-08, 6.293534e-08, 6.323759e-08, 6.35006e-08, 6.374071e-08, 
    6.372311e-08, 6.372931e-08, 6.378295e-08, 6.365008e-08, 6.380476e-08, 
    6.383071e-08, 6.376284e-08, 6.415675e-08, 6.404422e-08, 6.415937e-08, 
    6.40861e-08, 6.22443e-08, 6.233561e-08, 6.228627e-08, 6.237905e-08, 
    6.231368e-08, 6.260434e-08, 6.269149e-08, 6.309931e-08, 6.293195e-08, 
    6.319831e-08, 6.2959e-08, 6.300141e-08, 6.320698e-08, 6.297194e-08, 
    6.348608e-08, 6.313749e-08, 6.378503e-08, 6.343689e-08, 6.380684e-08, 
    6.373967e-08, 6.38509e-08, 6.395051e-08, 6.407584e-08, 6.430709e-08, 
    6.425354e-08, 6.444694e-08, 6.247174e-08, 6.259017e-08, 6.257976e-08, 
    6.270371e-08, 6.279537e-08, 6.299408e-08, 6.331277e-08, 6.319293e-08, 
    6.341295e-08, 6.345712e-08, 6.312285e-08, 6.332808e-08, 6.266944e-08, 
    6.277585e-08, 6.27125e-08, 6.248108e-08, 6.322053e-08, 6.284102e-08, 
    6.354184e-08, 6.333624e-08, 6.393631e-08, 6.363786e-08, 6.422406e-08, 
    6.447465e-08, 6.471054e-08, 6.498618e-08, 6.265482e-08, 6.257435e-08, 
    6.271845e-08, 6.291781e-08, 6.310282e-08, 6.334877e-08, 6.337395e-08, 
    6.342002e-08, 6.353938e-08, 6.363974e-08, 6.343458e-08, 6.36649e-08, 
    6.28005e-08, 6.325348e-08, 6.254392e-08, 6.275756e-08, 6.290607e-08, 
    6.284093e-08, 6.317924e-08, 6.325897e-08, 6.358299e-08, 6.341549e-08, 
    6.44128e-08, 6.397154e-08, 6.519609e-08, 6.485385e-08, 6.254623e-08, 
    6.265455e-08, 6.303155e-08, 6.285217e-08, 6.33652e-08, 6.349148e-08, 
    6.359415e-08, 6.372539e-08, 6.373956e-08, 6.381732e-08, 6.36899e-08, 
    6.381229e-08, 6.33493e-08, 6.355619e-08, 6.298847e-08, 6.312663e-08, 
    6.306308e-08, 6.299335e-08, 6.320855e-08, 6.343781e-08, 6.344272e-08, 
    6.351623e-08, 6.372337e-08, 6.336728e-08, 6.446972e-08, 6.378883e-08, 
    6.277267e-08, 6.298131e-08, 6.301112e-08, 6.29303e-08, 6.347882e-08, 
    6.328006e-08, 6.381542e-08, 6.367073e-08, 6.390781e-08, 6.379e-08, 
    6.377267e-08, 6.362136e-08, 6.352716e-08, 6.328918e-08, 6.309555e-08, 
    6.294202e-08, 6.297773e-08, 6.314637e-08, 6.345184e-08, 6.374083e-08, 
    6.367753e-08, 6.388979e-08, 6.3328e-08, 6.356355e-08, 6.347251e-08, 
    6.370992e-08, 6.318974e-08, 6.363265e-08, 6.307653e-08, 6.312529e-08, 
    6.327612e-08, 6.357952e-08, 6.364667e-08, 6.371835e-08, 6.367412e-08, 
    6.345959e-08, 6.342446e-08, 6.327246e-08, 6.323049e-08, 6.311468e-08, 
    6.301879e-08, 6.310639e-08, 6.319839e-08, 6.345969e-08, 6.369518e-08, 
    6.395192e-08, 6.401477e-08, 6.431474e-08, 6.407053e-08, 6.447351e-08, 
    6.413087e-08, 6.472403e-08, 6.365835e-08, 6.412082e-08, 6.328299e-08, 
    6.337325e-08, 6.353649e-08, 6.391095e-08, 6.37088e-08, 6.394522e-08, 
    6.342308e-08, 6.315219e-08, 6.308211e-08, 6.295136e-08, 6.30851e-08, 
    6.307422e-08, 6.320221e-08, 6.316108e-08, 6.346837e-08, 6.33033e-08, 
    6.377223e-08, 6.394335e-08, 6.442666e-08, 6.472296e-08, 6.502461e-08, 
    6.515778e-08, 6.519831e-08, 6.521526e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999957, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 
    0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999957, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3396233, -0.339628, -0.3396271, -0.339631, -0.3396289, -0.3396314, 
    -0.3396243, -0.3396282, -0.3396257, -0.3396237, -0.3396385, -0.3396312, 
    -0.3396466, -0.3396418, -0.3396539, -0.3396458, -0.3396555, -0.3396538, 
    -0.3396594, -0.3396578, -0.3396648, -0.3396602, -0.3396686, -0.3396638, 
    -0.3396645, -0.33966, -0.3396328, -0.3396376, -0.3396325, -0.3396332, 
    -0.3396329, -0.3396289, -0.3396268, -0.339623, -0.3396237, -0.3396266, 
    -0.3396335, -0.3396312, -0.3396372, -0.339637, -0.3396436, -0.3396406, 
    -0.3396518, -0.3396487, -0.3396579, -0.3396555, -0.3396578, -0.3396571, 
    -0.3396578, -0.3396543, -0.3396558, -0.3396528, -0.3396412, -0.3396446, 
    -0.3396344, -0.3396282, -0.3396244, -0.3396217, -0.3396221, -0.3396228, 
    -0.3396266, -0.3396303, -0.3396332, -0.3396351, -0.339637, -0.3396425, 
    -0.3396456, -0.3396524, -0.3396513, -0.3396533, -0.3396553, -0.3396586, 
    -0.3396581, -0.3396595, -0.3396533, -0.3396574, -0.3396506, -0.3396524, 
    -0.3396372, -0.3396318, -0.3396292, -0.3396273, -0.3396224, -0.3396257, 
    -0.3396244, -0.3396277, -0.3396297, -0.3396287, -0.3396352, -0.3396326, 
    -0.3396458, -0.3396401, -0.3396551, -0.3396515, -0.3396559, -0.3396537, 
    -0.3396575, -0.3396541, -0.3396601, -0.3396614, -0.3396605, -0.339664, 
    -0.3396539, -0.3396577, -0.3396287, -0.3396288, -0.3396297, -0.3396262, 
    -0.339626, -0.3396229, -0.3396257, -0.3396268, -0.3396299, -0.3396317, 
    -0.3396334, -0.3396372, -0.3396414, -0.3396474, -0.3396517, -0.3396546, 
    -0.3396529, -0.3396544, -0.3396527, -0.3396519, -0.3396609, -0.3396558, 
    -0.3396635, -0.3396631, -0.3396595, -0.3396631, -0.339629, -0.339628, 
    -0.3396247, -0.3396273, -0.3396226, -0.3396252, -0.3396266, -0.3396326, 
    -0.339634, -0.3396352, -0.3396377, -0.3396408, -0.3396462, -0.339651, 
    -0.3396554, -0.3396551, -0.3396552, -0.3396562, -0.3396538, -0.3396566, 
    -0.339657, -0.3396558, -0.339663, -0.3396609, -0.3396631, -0.3396617, 
    -0.3396283, -0.3396299, -0.3396291, -0.3396307, -0.3396295, -0.3396347, 
    -0.3396363, -0.3396437, -0.3396407, -0.3396455, -0.3396412, -0.339642, 
    -0.3396455, -0.3396415, -0.3396507, -0.3396443, -0.3396562, -0.3396497, 
    -0.3396566, -0.3396554, -0.3396575, -0.3396592, -0.3396615, -0.3396657, 
    -0.3396647, -0.3396683, -0.3396324, -0.3396345, -0.3396344, -0.3396366, 
    -0.3396382, -0.3396419, -0.3396476, -0.3396455, -0.3396495, -0.3396503, 
    -0.3396442, -0.3396479, -0.3396359, -0.3396378, -0.3396367, -0.3396325, 
    -0.3396459, -0.339639, -0.3396518, -0.3396481, -0.339659, -0.3396535, 
    -0.3396642, -0.3396686, -0.3396731, -0.339678, -0.3396357, -0.3396343, 
    -0.3396369, -0.3396404, -0.3396438, -0.3396483, -0.3396488, -0.3396496, 
    -0.3396518, -0.3396536, -0.3396498, -0.3396541, -0.3396381, -0.3396465, 
    -0.3396337, -0.3396375, -0.3396402, -0.3396391, -0.3396452, -0.3396467, 
    -0.3396525, -0.3396495, -0.3396675, -0.3396595, -0.3396819, -0.3396756, 
    -0.3396338, -0.3396357, -0.3396425, -0.3396393, -0.3396486, -0.3396509, 
    -0.3396528, -0.3396551, -0.3396554, -0.3396568, -0.3396545, -0.3396567, 
    -0.3396483, -0.3396521, -0.3396418, -0.3396443, -0.3396431, -0.3396419, 
    -0.3396458, -0.3396498, -0.33965, -0.3396513, -0.3396547, -0.3396486, 
    -0.3396683, -0.339656, -0.3396379, -0.3396415, -0.3396422, -0.3396407, 
    -0.3396506, -0.339647, -0.3396568, -0.3396542, -0.3396585, -0.3396563, 
    -0.339656, -0.3396533, -0.3396515, -0.3396472, -0.3396437, -0.3396409, 
    -0.3396416, -0.3396446, -0.3396501, -0.3396554, -0.3396542, -0.3396581, 
    -0.3396479, -0.3396522, -0.3396505, -0.3396549, -0.3396454, -0.3396531, 
    -0.3396434, -0.3396443, -0.339647, -0.3396524, -0.3396537, -0.339655, 
    -0.3396542, -0.3396502, -0.3396496, -0.3396469, -0.3396461, -0.3396441, 
    -0.3396423, -0.3396439, -0.3396455, -0.3396503, -0.3396546, -0.3396592, 
    -0.3396604, -0.3396657, -0.3396612, -0.3396684, -0.3396621, -0.3396731, 
    -0.3396537, -0.3396621, -0.3396471, -0.3396488, -0.3396516, -0.3396584, 
    -0.3396548, -0.339659, -0.3396496, -0.3396446, -0.3396435, -0.3396411, 
    -0.3396435, -0.3396433, -0.3396457, -0.3396449, -0.3396505, -0.3396475, 
    -0.339656, -0.339659, -0.3396679, -0.3396732, -0.3396789, -0.3396813, 
    -0.339682, -0.3396823 ;

 TAUY =
  -0.3396233, -0.339628, -0.3396271, -0.339631, -0.3396289, -0.3396314, 
    -0.3396243, -0.3396282, -0.3396257, -0.3396237, -0.3396385, -0.3396312, 
    -0.3396466, -0.3396418, -0.3396539, -0.3396458, -0.3396555, -0.3396538, 
    -0.3396594, -0.3396578, -0.3396648, -0.3396602, -0.3396686, -0.3396638, 
    -0.3396645, -0.33966, -0.3396328, -0.3396376, -0.3396325, -0.3396332, 
    -0.3396329, -0.3396289, -0.3396268, -0.339623, -0.3396237, -0.3396266, 
    -0.3396335, -0.3396312, -0.3396372, -0.339637, -0.3396436, -0.3396406, 
    -0.3396518, -0.3396487, -0.3396579, -0.3396555, -0.3396578, -0.3396571, 
    -0.3396578, -0.3396543, -0.3396558, -0.3396528, -0.3396412, -0.3396446, 
    -0.3396344, -0.3396282, -0.3396244, -0.3396217, -0.3396221, -0.3396228, 
    -0.3396266, -0.3396303, -0.3396332, -0.3396351, -0.339637, -0.3396425, 
    -0.3396456, -0.3396524, -0.3396513, -0.3396533, -0.3396553, -0.3396586, 
    -0.3396581, -0.3396595, -0.3396533, -0.3396574, -0.3396506, -0.3396524, 
    -0.3396372, -0.3396318, -0.3396292, -0.3396273, -0.3396224, -0.3396257, 
    -0.3396244, -0.3396277, -0.3396297, -0.3396287, -0.3396352, -0.3396326, 
    -0.3396458, -0.3396401, -0.3396551, -0.3396515, -0.3396559, -0.3396537, 
    -0.3396575, -0.3396541, -0.3396601, -0.3396614, -0.3396605, -0.339664, 
    -0.3396539, -0.3396577, -0.3396287, -0.3396288, -0.3396297, -0.3396262, 
    -0.339626, -0.3396229, -0.3396257, -0.3396268, -0.3396299, -0.3396317, 
    -0.3396334, -0.3396372, -0.3396414, -0.3396474, -0.3396517, -0.3396546, 
    -0.3396529, -0.3396544, -0.3396527, -0.3396519, -0.3396609, -0.3396558, 
    -0.3396635, -0.3396631, -0.3396595, -0.3396631, -0.339629, -0.339628, 
    -0.3396247, -0.3396273, -0.3396226, -0.3396252, -0.3396266, -0.3396326, 
    -0.339634, -0.3396352, -0.3396377, -0.3396408, -0.3396462, -0.339651, 
    -0.3396554, -0.3396551, -0.3396552, -0.3396562, -0.3396538, -0.3396566, 
    -0.339657, -0.3396558, -0.339663, -0.3396609, -0.3396631, -0.3396617, 
    -0.3396283, -0.3396299, -0.3396291, -0.3396307, -0.3396295, -0.3396347, 
    -0.3396363, -0.3396437, -0.3396407, -0.3396455, -0.3396412, -0.339642, 
    -0.3396455, -0.3396415, -0.3396507, -0.3396443, -0.3396562, -0.3396497, 
    -0.3396566, -0.3396554, -0.3396575, -0.3396592, -0.3396615, -0.3396657, 
    -0.3396647, -0.3396683, -0.3396324, -0.3396345, -0.3396344, -0.3396366, 
    -0.3396382, -0.3396419, -0.3396476, -0.3396455, -0.3396495, -0.3396503, 
    -0.3396442, -0.3396479, -0.3396359, -0.3396378, -0.3396367, -0.3396325, 
    -0.3396459, -0.339639, -0.3396518, -0.3396481, -0.339659, -0.3396535, 
    -0.3396642, -0.3396686, -0.3396731, -0.339678, -0.3396357, -0.3396343, 
    -0.3396369, -0.3396404, -0.3396438, -0.3396483, -0.3396488, -0.3396496, 
    -0.3396518, -0.3396536, -0.3396498, -0.3396541, -0.3396381, -0.3396465, 
    -0.3396337, -0.3396375, -0.3396402, -0.3396391, -0.3396452, -0.3396467, 
    -0.3396525, -0.3396495, -0.3396675, -0.3396595, -0.3396819, -0.3396756, 
    -0.3396338, -0.3396357, -0.3396425, -0.3396393, -0.3396486, -0.3396509, 
    -0.3396528, -0.3396551, -0.3396554, -0.3396568, -0.3396545, -0.3396567, 
    -0.3396483, -0.3396521, -0.3396418, -0.3396443, -0.3396431, -0.3396419, 
    -0.3396458, -0.3396498, -0.33965, -0.3396513, -0.3396547, -0.3396486, 
    -0.3396683, -0.339656, -0.3396379, -0.3396415, -0.3396422, -0.3396407, 
    -0.3396506, -0.339647, -0.3396568, -0.3396542, -0.3396585, -0.3396563, 
    -0.339656, -0.3396533, -0.3396515, -0.3396472, -0.3396437, -0.3396409, 
    -0.3396416, -0.3396446, -0.3396501, -0.3396554, -0.3396542, -0.3396581, 
    -0.3396479, -0.3396522, -0.3396505, -0.3396549, -0.3396454, -0.3396531, 
    -0.3396434, -0.3396443, -0.339647, -0.3396524, -0.3396537, -0.339655, 
    -0.3396542, -0.3396502, -0.3396496, -0.3396469, -0.3396461, -0.3396441, 
    -0.3396423, -0.3396439, -0.3396455, -0.3396503, -0.3396546, -0.3396592, 
    -0.3396604, -0.3396657, -0.3396612, -0.3396684, -0.3396621, -0.3396731, 
    -0.3396537, -0.3396621, -0.3396471, -0.3396488, -0.3396516, -0.3396584, 
    -0.3396548, -0.339659, -0.3396496, -0.3396446, -0.3396435, -0.3396411, 
    -0.3396435, -0.3396433, -0.3396457, -0.3396449, -0.3396505, -0.3396475, 
    -0.339656, -0.339659, -0.3396679, -0.3396732, -0.3396789, -0.3396813, 
    -0.339682, -0.3396823 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.114, 261.1351, 261.131, 261.1479, 261.1385, 261.1497, 261.1183, 
    261.1359, 261.1247, 261.1159, 261.1808, 261.1487, 261.2143, 261.1938, 
    261.2453, 261.2111, 261.2521, 261.2443, 261.268, 261.2612, 261.2915, 
    261.2711, 261.3072, 261.2866, 261.2898, 261.2704, 261.1552, 261.1768, 
    261.1539, 261.157, 261.1556, 261.1387, 261.1302, 261.1124, 261.1157, 
    261.1287, 261.1584, 261.1483, 261.1737, 261.1731, 261.2014, 261.1886, 
    261.236, 261.2226, 261.2615, 261.2517, 261.261, 261.2582, 261.261, 
    261.2467, 261.2528, 261.2402, 261.191, 261.2055, 261.1623, 261.1363, 
    261.1191, 261.1068, 261.1086, 261.1118, 261.1288, 261.1448, 261.1569, 
    261.165, 261.173, 261.1972, 261.2101, 261.2387, 261.2336, 261.2423, 
    261.2507, 261.2648, 261.2625, 261.2686, 261.2421, 261.2597, 261.2307, 
    261.2386, 261.1752, 261.1511, 261.1407, 261.1318, 261.1099, 261.125, 
    261.119, 261.1332, 261.1422, 261.1378, 261.1653, 261.1546, 261.2108, 
    261.1866, 261.2498, 261.2346, 261.2534, 261.2438, 261.2602, 261.2455, 
    261.271, 261.2765, 261.2727, 261.2873, 261.2446, 261.261, 261.1377, 
    261.1384, 261.1418, 261.1269, 261.126, 261.1123, 261.1245, 261.1296, 
    261.1428, 261.1505, 261.1579, 261.1741, 261.1922, 261.2175, 261.2356, 
    261.2478, 261.2403, 261.2469, 261.2396, 261.2361, 261.2744, 261.2529, 
    261.2852, 261.2834, 261.2688, 261.2836, 261.1389, 261.1347, 261.1202, 
    261.1316, 261.1108, 261.1224, 261.1291, 261.1548, 261.1605, 261.1657, 
    261.176, 261.1893, 261.2125, 261.2328, 261.2512, 261.2498, 261.2503, 
    261.2545, 261.2442, 261.2561, 261.2581, 261.2529, 261.2832, 261.2745, 
    261.2834, 261.2777, 261.1361, 261.1431, 261.1393, 261.1465, 261.1414, 
    261.1638, 261.1705, 261.2019, 261.189, 261.2095, 261.1911, 261.1944, 
    261.2101, 261.1921, 261.2316, 261.2048, 261.2546, 261.2278, 261.2563, 
    261.2511, 261.2597, 261.2673, 261.2769, 261.2947, 261.2906, 261.3054, 
    261.1536, 261.1627, 261.1619, 261.1714, 261.1785, 261.1938, 261.2183, 
    261.2091, 261.226, 261.2294, 261.2037, 261.2195, 261.1688, 261.177, 
    261.1721, 261.1543, 261.2112, 261.182, 261.2359, 261.2201, 261.2662, 
    261.2433, 261.2883, 261.3076, 261.3257, 261.3468, 261.1677, 261.1615, 
    261.1726, 261.1879, 261.2021, 261.2211, 261.223, 261.2266, 261.2357, 
    261.2434, 261.2277, 261.2454, 261.1789, 261.2137, 261.1591, 261.1756, 
    261.187, 261.182, 261.208, 261.2142, 261.2391, 261.2262, 261.3028, 
    261.2689, 261.3629, 261.3366, 261.1593, 261.1677, 261.1967, 261.1829, 
    261.2224, 261.2321, 261.24, 261.25, 261.2511, 261.2571, 261.2473, 
    261.2567, 261.2211, 261.237, 261.1934, 261.204, 261.1991, 261.1938, 
    261.2103, 261.2279, 261.2283, 261.2339, 261.2498, 261.2225, 261.3071, 
    261.2549, 261.1768, 261.1928, 261.1951, 261.1889, 261.2311, 261.2158, 
    261.257, 261.2458, 261.264, 261.255, 261.2537, 261.242, 261.2348, 
    261.2165, 261.2016, 261.1898, 261.1925, 261.2055, 261.229, 261.2512, 
    261.2463, 261.2627, 261.2195, 261.2376, 261.2306, 261.2488, 261.2089, 
    261.2429, 261.2001, 261.2039, 261.2155, 261.2388, 261.244, 261.2495, 
    261.2461, 261.2296, 261.2269, 261.2152, 261.212, 261.2031, 261.1957, 
    261.2024, 261.2095, 261.2296, 261.2477, 261.2674, 261.2723, 261.2953, 
    261.2765, 261.3074, 261.2811, 261.3267, 261.2448, 261.2804, 261.216, 
    261.223, 261.2355, 261.2643, 261.2487, 261.2669, 261.2268, 261.206, 
    261.2006, 261.1905, 261.2008, 261.2, 261.2098, 261.2066, 261.2303, 
    261.2176, 261.2536, 261.2668, 261.3039, 261.3266, 261.3497, 261.3599, 
    261.363, 261.3643 ;

 TG_R =
  261.114, 261.1351, 261.131, 261.1479, 261.1385, 261.1497, 261.1183, 
    261.1359, 261.1247, 261.1159, 261.1808, 261.1487, 261.2143, 261.1938, 
    261.2453, 261.2111, 261.2521, 261.2443, 261.268, 261.2612, 261.2915, 
    261.2711, 261.3072, 261.2866, 261.2898, 261.2704, 261.1552, 261.1768, 
    261.1539, 261.157, 261.1556, 261.1387, 261.1302, 261.1124, 261.1157, 
    261.1287, 261.1584, 261.1483, 261.1737, 261.1731, 261.2014, 261.1886, 
    261.236, 261.2226, 261.2615, 261.2517, 261.261, 261.2582, 261.261, 
    261.2467, 261.2528, 261.2402, 261.191, 261.2055, 261.1623, 261.1363, 
    261.1191, 261.1068, 261.1086, 261.1118, 261.1288, 261.1448, 261.1569, 
    261.165, 261.173, 261.1972, 261.2101, 261.2387, 261.2336, 261.2423, 
    261.2507, 261.2648, 261.2625, 261.2686, 261.2421, 261.2597, 261.2307, 
    261.2386, 261.1752, 261.1511, 261.1407, 261.1318, 261.1099, 261.125, 
    261.119, 261.1332, 261.1422, 261.1378, 261.1653, 261.1546, 261.2108, 
    261.1866, 261.2498, 261.2346, 261.2534, 261.2438, 261.2602, 261.2455, 
    261.271, 261.2765, 261.2727, 261.2873, 261.2446, 261.261, 261.1377, 
    261.1384, 261.1418, 261.1269, 261.126, 261.1123, 261.1245, 261.1296, 
    261.1428, 261.1505, 261.1579, 261.1741, 261.1922, 261.2175, 261.2356, 
    261.2478, 261.2403, 261.2469, 261.2396, 261.2361, 261.2744, 261.2529, 
    261.2852, 261.2834, 261.2688, 261.2836, 261.1389, 261.1347, 261.1202, 
    261.1316, 261.1108, 261.1224, 261.1291, 261.1548, 261.1605, 261.1657, 
    261.176, 261.1893, 261.2125, 261.2328, 261.2512, 261.2498, 261.2503, 
    261.2545, 261.2442, 261.2561, 261.2581, 261.2529, 261.2832, 261.2745, 
    261.2834, 261.2777, 261.1361, 261.1431, 261.1393, 261.1465, 261.1414, 
    261.1638, 261.1705, 261.2019, 261.189, 261.2095, 261.1911, 261.1944, 
    261.2101, 261.1921, 261.2316, 261.2048, 261.2546, 261.2278, 261.2563, 
    261.2511, 261.2597, 261.2673, 261.2769, 261.2947, 261.2906, 261.3054, 
    261.1536, 261.1627, 261.1619, 261.1714, 261.1785, 261.1938, 261.2183, 
    261.2091, 261.226, 261.2294, 261.2037, 261.2195, 261.1688, 261.177, 
    261.1721, 261.1543, 261.2112, 261.182, 261.2359, 261.2201, 261.2662, 
    261.2433, 261.2883, 261.3076, 261.3257, 261.3468, 261.1677, 261.1615, 
    261.1726, 261.1879, 261.2021, 261.2211, 261.223, 261.2266, 261.2357, 
    261.2434, 261.2277, 261.2454, 261.1789, 261.2137, 261.1591, 261.1756, 
    261.187, 261.182, 261.208, 261.2142, 261.2391, 261.2262, 261.3028, 
    261.2689, 261.3629, 261.3366, 261.1593, 261.1677, 261.1967, 261.1829, 
    261.2224, 261.2321, 261.24, 261.25, 261.2511, 261.2571, 261.2473, 
    261.2567, 261.2211, 261.237, 261.1934, 261.204, 261.1991, 261.1938, 
    261.2103, 261.2279, 261.2283, 261.2339, 261.2498, 261.2225, 261.3071, 
    261.2549, 261.1768, 261.1928, 261.1951, 261.1889, 261.2311, 261.2158, 
    261.257, 261.2458, 261.264, 261.255, 261.2537, 261.242, 261.2348, 
    261.2165, 261.2016, 261.1898, 261.1925, 261.2055, 261.229, 261.2512, 
    261.2463, 261.2627, 261.2195, 261.2376, 261.2306, 261.2488, 261.2089, 
    261.2429, 261.2001, 261.2039, 261.2155, 261.2388, 261.244, 261.2495, 
    261.2461, 261.2296, 261.2269, 261.2152, 261.212, 261.2031, 261.1957, 
    261.2024, 261.2095, 261.2296, 261.2477, 261.2674, 261.2723, 261.2953, 
    261.2765, 261.3074, 261.2811, 261.3267, 261.2448, 261.2804, 261.216, 
    261.223, 261.2355, 261.2643, 261.2487, 261.2669, 261.2268, 261.206, 
    261.2006, 261.1905, 261.2008, 261.2, 261.2098, 261.2066, 261.2303, 
    261.2176, 261.2536, 261.2668, 261.3039, 261.3266, 261.3497, 261.3599, 
    261.363, 261.3643 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.4839, 254.4854, 254.4851, 254.4863, 254.4857, 254.4865, 254.4842, 
    254.4855, 254.4847, 254.4841, 254.4886, 254.4864, 254.491, 254.4896, 
    254.4932, 254.4908, 254.4937, 254.4932, 254.4949, 254.4944, 254.4966, 
    254.4951, 254.4977, 254.4962, 254.4964, 254.4951, 254.4868, 254.4883, 
    254.4868, 254.487, 254.4869, 254.4857, 254.4851, 254.4838, 254.4841, 
    254.485, 254.4871, 254.4864, 254.4882, 254.4881, 254.4901, 254.4892, 
    254.4926, 254.4916, 254.4944, 254.4937, 254.4944, 254.4942, 254.4944, 
    254.4934, 254.4938, 254.4929, 254.4894, 254.4904, 254.4874, 254.4855, 
    254.4843, 254.4834, 254.4836, 254.4838, 254.485, 254.4861, 254.487, 
    254.4875, 254.4881, 254.4898, 254.4907, 254.4928, 254.4924, 254.493, 
    254.4937, 254.4947, 254.4945, 254.4949, 254.493, 254.4943, 254.4922, 
    254.4928, 254.4882, 254.4866, 254.4858, 254.4852, 254.4837, 254.4847, 
    254.4843, 254.4853, 254.4859, 254.4856, 254.4876, 254.4868, 254.4908, 
    254.4891, 254.4936, 254.4925, 254.4939, 254.4932, 254.4943, 254.4933, 
    254.4951, 254.4955, 254.4952, 254.4963, 254.4932, 254.4944, 254.4856, 
    254.4857, 254.4859, 254.4848, 254.4848, 254.4838, 254.4847, 254.485, 
    254.486, 254.4865, 254.487, 254.4882, 254.4895, 254.4913, 254.4926, 
    254.4935, 254.4929, 254.4934, 254.4929, 254.4926, 254.4953, 254.4938, 
    254.4961, 254.496, 254.4949, 254.496, 254.4857, 254.4854, 254.4844, 
    254.4852, 254.4837, 254.4845, 254.485, 254.4868, 254.4872, 254.4876, 
    254.4883, 254.4893, 254.4909, 254.4924, 254.4937, 254.4936, 254.4936, 
    254.4939, 254.4932, 254.494, 254.4942, 254.4938, 254.496, 254.4954, 
    254.496, 254.4956, 254.4855, 254.486, 254.4857, 254.4862, 254.4859, 
    254.4874, 254.4879, 254.4901, 254.4892, 254.4907, 254.4894, 254.4896, 
    254.4907, 254.4895, 254.4923, 254.4903, 254.4939, 254.492, 254.494, 
    254.4937, 254.4943, 254.4948, 254.4955, 254.4968, 254.4965, 254.4976, 
    254.4867, 254.4874, 254.4873, 254.488, 254.4885, 254.4896, 254.4913, 
    254.4907, 254.4919, 254.4921, 254.4903, 254.4914, 254.4878, 254.4884, 
    254.4881, 254.4868, 254.4908, 254.4887, 254.4926, 254.4915, 254.4948, 
    254.4931, 254.4964, 254.4977, 254.4991, 254.5005, 254.4877, 254.4873, 
    254.4881, 254.4892, 254.4902, 254.4915, 254.4917, 254.4919, 254.4926, 
    254.4931, 254.492, 254.4933, 254.4885, 254.491, 254.4871, 254.4883, 
    254.4891, 254.4888, 254.4906, 254.491, 254.4928, 254.4919, 254.4974, 
    254.4949, 254.5017, 254.4998, 254.4872, 254.4877, 254.4898, 254.4888, 
    254.4916, 254.4923, 254.4929, 254.4936, 254.4937, 254.4941, 254.4934, 
    254.4941, 254.4915, 254.4927, 254.4896, 254.4903, 254.49, 254.4896, 
    254.4908, 254.492, 254.4921, 254.4924, 254.4935, 254.4916, 254.4977, 
    254.4939, 254.4884, 254.4895, 254.4897, 254.4892, 254.4922, 254.4911, 
    254.4941, 254.4933, 254.4946, 254.494, 254.4939, 254.493, 254.4925, 
    254.4912, 254.4901, 254.4893, 254.4895, 254.4904, 254.4921, 254.4937, 
    254.4933, 254.4945, 254.4914, 254.4927, 254.4922, 254.4935, 254.4907, 
    254.493, 254.4901, 254.4903, 254.4911, 254.4928, 254.4932, 254.4936, 
    254.4933, 254.4921, 254.4919, 254.4911, 254.4909, 254.4902, 254.4897, 
    254.4902, 254.4907, 254.4921, 254.4934, 254.4948, 254.4952, 254.4968, 
    254.4955, 254.4977, 254.4958, 254.4991, 254.4932, 254.4957, 254.4912, 
    254.4917, 254.4926, 254.4946, 254.4935, 254.4948, 254.4919, 254.4904, 
    254.4901, 254.4893, 254.4901, 254.49, 254.4907, 254.4905, 254.4922, 
    254.4913, 254.4939, 254.4948, 254.4975, 254.4991, 254.5008, 254.5015, 
    254.5018, 254.5019 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24017, 18.24017, 18.24018, 
    18.24017, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24016, 18.24016, 18.24016, 18.24017, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24013, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24017, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24011, 18.24011, 18.24011, 18.2401, 
    18.24009, 18.2401, 18.24009, 18.24011, 18.2401, 18.24011, 18.24011, 
    18.24015, 18.24016, 18.24017, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24018, 18.24017, 18.24017, 18.24016, 18.24016, 18.24013, 18.24014, 
    18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 18.24009, 
    18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24017, 18.24017, 
    18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24015, 18.24014, 18.24012, 18.24011, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24018, 18.24018, 
    18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 18.24008, 
    18.24009, 18.24017, 18.24017, 18.24017, 18.24017, 18.24017, 18.24016, 
    18.24015, 18.24013, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24014, 18.24011, 18.24013, 18.2401, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24007, 18.24008, 18.24007, 18.24016, 
    18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24012, 18.24013, 
    18.24012, 18.24012, 18.24013, 18.24012, 18.24015, 18.24015, 18.24015, 
    18.24016, 18.24013, 18.24014, 18.24011, 18.24012, 18.24009, 18.24011, 
    18.24008, 18.24007, 18.24006, 18.24004, 18.24015, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24012, 18.24012, 18.24012, 18.24011, 18.24011, 
    18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 18.24014, 
    18.24014, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 18.24009, 
    18.24003, 18.24005, 18.24016, 18.24015, 18.24014, 18.24014, 18.24012, 
    18.24011, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 18.2401, 
    18.24015, 18.24014, 18.24014, 18.24014, 18.24011, 18.24012, 18.2401, 
    18.2401, 18.24009, 18.2401, 18.2401, 18.24011, 18.24011, 18.24012, 
    18.24013, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24012, 18.24011, 18.24011, 18.2401, 18.24013, 18.24011, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.24011, 18.2401, 18.2401, 
    18.24012, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.2401, 18.24009, 18.24009, 18.24007, 18.24009, 
    18.24007, 18.24008, 18.24006, 18.24011, 18.24008, 18.24012, 18.24012, 
    18.24011, 18.24009, 18.2401, 18.24009, 18.24012, 18.24013, 18.24013, 
    18.24014, 18.24013, 18.24013, 18.24013, 18.24013, 18.24012, 18.24012, 
    18.2401, 18.24009, 18.24007, 18.24006, 18.24004, 18.24003, 18.24003, 
    18.24003 ;

 TOTCOLCH4 =
  4.303581e-06, 4.166393e-06, 4.192906e-06, 4.083431e-06, 4.143999e-06, 
    4.072551e-06, 4.27561e-06, 4.160982e-06, 4.233996e-06, 4.291159e-06, 
    3.874851e-06, 4.078581e-06, 3.668583e-06, 3.794623e-06, 3.481943e-06, 
    3.688051e-06, 3.441088e-06, 3.487827e-06, 3.348133e-06, 3.387868e-06, 
    3.212222e-06, 3.329872e-06, 3.123027e-06, 3.240138e-06, 3.221669e-06, 
    3.333786e-06, 4.037204e-06, 3.899939e-06, 4.045403e-06, 4.025674e-06, 
    4.034525e-06, 4.142737e-06, 4.197763e-06, 4.314165e-06, 4.292927e-06, 
    4.207493e-06, 4.016817e-06, 4.081092e-06, 3.920069e-06, 3.923672e-06, 
    3.747942e-06, 3.826698e-06, 3.537143e-06, 3.618324e-06, 3.386205e-06, 
    3.443869e-06, 3.3889e-06, 3.405524e-06, 3.388683e-06, 3.473449e-06, 
    3.437005e-06, 3.512062e-06, 3.811885e-06, 3.722533e-06, 3.992002e-06, 
    4.158292e-06, 4.270548e-06, 4.351033e-06, 4.339613e-06, 4.317875e-06, 
    4.206996e-06, 4.103991e-06, 4.026293e-06, 3.974707e-06, 3.92419e-06, 
    3.773101e-06, 3.694327e-06, 3.520827e-06, 3.551855e-06, 3.499382e-06, 
    3.449633e-06, 3.366872e-06, 3.380428e-06, 3.344204e-06, 3.500774e-06, 
    3.396319e-06, 3.569584e-06, 3.521774e-06, 3.91044e-06, 4.063708e-06, 
    4.129634e-06, 4.187801e-06, 4.33084e-06, 4.231817e-06, 4.270724e-06, 
    4.17845e-06, 4.120296e-06, 4.149013e-06, 3.973301e-06, 4.041185e-06, 
    3.689683e-06, 3.839216e-06, 3.455418e-06, 3.545477e-06, 3.434002e-06, 
    3.490671e-06, 3.393845e-06, 3.480927e-06, 3.330776e-06, 3.298506e-06, 
    3.32054e-06, 3.236316e-06, 3.485785e-06, 3.388894e-06, 4.149816e-06, 
    4.145125e-06, 4.123312e-06, 4.219595e-06, 4.225523e-06, 4.314745e-06, 
    4.235319e-06, 4.201699e-06, 4.116942e-06, 4.067177e-06, 4.020138e-06, 
    3.917626e-06, 3.804615e-06, 3.649267e-06, 3.539604e-06, 3.467004e-06, 
    3.511439e-06, 3.472194e-06, 3.516076e-06, 3.53674e-06, 3.310575e-06, 
    3.436662e-06, 3.248364e-06, 3.258649e-06, 3.343342e-06, 3.257489e-06, 
    4.141834e-06, 4.168849e-06, 4.263257e-06, 4.189291e-06, 4.324515e-06, 
    4.248568e-06, 4.205177e-06, 4.039745e-06, 4.003834e-06, 3.970647e-06, 
    3.905505e-06, 3.822648e-06, 3.679348e-06, 3.556827e-06, 3.446752e-06, 
    3.454761e-06, 3.45194e-06, 3.427556e-06, 3.488101e-06, 3.417667e-06, 
    3.405909e-06, 3.436684e-06, 3.260027e-06, 3.310028e-06, 3.258867e-06, 
    3.291377e-06, 4.160061e-06, 4.114699e-06, 4.13918e-06, 4.093197e-06, 
    4.125562e-06, 3.982547e-06, 3.940133e-06, 3.744562e-06, 3.824267e-06, 
    3.697814e-06, 3.811334e-06, 3.791095e-06, 3.693696e-06, 3.805162e-06, 
    3.563517e-06, 3.726485e-06, 3.42661e-06, 3.586288e-06, 3.416721e-06, 
    3.447224e-06, 3.3968e-06, 3.351942e-06, 3.295937e-06, 3.193808e-06, 
    3.217318e-06, 3.132836e-06, 4.047514e-06, 3.989473e-06, 3.99458e-06, 
    3.934237e-06, 3.889887e-06, 3.7946e-06, 3.644126e-06, 3.700371e-06, 
    3.597448e-06, 3.576951e-06, 3.733448e-06, 3.636966e-06, 3.95086e-06, 
    3.899291e-06, 3.929966e-06, 4.042914e-06, 3.687356e-06, 3.867872e-06, 
    3.537803e-06, 3.633168e-06, 3.358318e-06, 3.493673e-06, 3.230294e-06, 
    3.120789e-06, 3.019505e-06, 2.903209e-06, 3.957977e-06, 3.997224e-06, 
    3.927094e-06, 3.831014e-06, 3.742922e-06, 3.627314e-06, 3.615592e-06, 
    3.594159e-06, 3.538945e-06, 3.492838e-06, 3.587383e-06, 3.481327e-06, 
    3.887352e-06, 3.671888e-06, 4.012097e-06, 3.908123e-06, 3.836652e-06, 
    3.86794e-06, 3.706829e-06, 3.669332e-06, 3.518856e-06, 3.596269e-06, 
    3.147631e-06, 3.342487e-06, 2.816246e-06, 2.958746e-06, 4.010976e-06, 
    3.958119e-06, 3.776737e-06, 3.862534e-06, 3.619666e-06, 3.561047e-06, 
    3.513748e-06, 3.453714e-06, 3.447272e-06, 3.411976e-06, 3.469907e-06, 
    3.41426e-06, 3.62707e-06, 3.531196e-06, 3.79728e-06, 3.73165e-06, 
    3.761778e-06, 3.79495e-06, 3.693021e-06, 3.585882e-06, 3.583629e-06, 
    3.549605e-06, 3.454546e-06, 3.618698e-06, 3.12287e-06, 3.424805e-06, 
    3.900858e-06, 3.800658e-06, 3.786472e-06, 3.825066e-06, 3.566902e-06, 
    3.659436e-06, 3.412837e-06, 3.47866e-06, 3.371138e-06, 3.424359e-06, 
    3.432222e-06, 3.501259e-06, 3.544574e-06, 3.655164e-06, 3.746363e-06, 
    3.819459e-06, 3.802404e-06, 3.722319e-06, 3.579382e-06, 3.44668e-06, 
    3.475537e-06, 3.379251e-06, 3.637019e-06, 3.527796e-06, 3.569813e-06, 
    3.460769e-06, 3.701866e-06, 3.495998e-06, 3.755395e-06, 3.732297e-06, 
    3.661284e-06, 3.520433e-06, 3.489664e-06, 3.456921e-06, 3.477112e-06, 
    3.575793e-06, 3.592097e-06, 3.663007e-06, 3.682694e-06, 3.737322e-06, 
    3.782831e-06, 3.741235e-06, 3.697786e-06, 3.575759e-06, 3.467485e-06, 
    3.351302e-06, 3.323174e-06, 3.190413e-06, 3.298257e-06, 3.121224e-06, 
    3.271386e-06, 3.013695e-06, 3.484274e-06, 3.275894e-06, 3.658075e-06, 
    3.615919e-06, 3.540249e-06, 3.369691e-06, 3.461278e-06, 3.354296e-06, 
    3.592738e-06, 3.71956e-06, 3.752744e-06, 3.814992e-06, 3.751327e-06, 
    3.756487e-06, 3.696006e-06, 3.715391e-06, 3.571742e-06, 3.648564e-06, 
    3.432415e-06, 3.35514e-06, 3.141631e-06, 3.01419e-06, 2.887218e-06, 
    2.832032e-06, 2.815343e-06, 2.808381e-06 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24017, 18.24017, 18.24018, 
    18.24017, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24016, 18.24016, 18.24016, 18.24017, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24013, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24017, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24011, 18.24011, 18.24011, 18.2401, 
    18.24009, 18.2401, 18.24009, 18.24011, 18.2401, 18.24011, 18.24011, 
    18.24015, 18.24016, 18.24017, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24018, 18.24017, 18.24017, 18.24016, 18.24016, 18.24013, 18.24014, 
    18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 18.24009, 
    18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24017, 18.24017, 
    18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24015, 18.24014, 18.24012, 18.24011, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24018, 18.24018, 
    18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 18.24008, 
    18.24009, 18.24017, 18.24017, 18.24017, 18.24017, 18.24017, 18.24016, 
    18.24015, 18.24013, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24014, 18.24011, 18.24013, 18.2401, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24007, 18.24008, 18.24007, 18.24016, 
    18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24012, 18.24013, 
    18.24012, 18.24012, 18.24013, 18.24012, 18.24015, 18.24015, 18.24015, 
    18.24016, 18.24013, 18.24014, 18.24011, 18.24012, 18.24009, 18.24011, 
    18.24008, 18.24007, 18.24006, 18.24004, 18.24015, 18.24016, 18.24015, 
    18.24014, 18.24013, 18.24012, 18.24012, 18.24012, 18.24011, 18.24011, 
    18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 18.24014, 
    18.24014, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 18.24009, 
    18.24003, 18.24005, 18.24016, 18.24015, 18.24014, 18.24014, 18.24012, 
    18.24011, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 18.24013, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 18.2401, 
    18.24015, 18.24014, 18.24014, 18.24014, 18.24011, 18.24012, 18.2401, 
    18.2401, 18.24009, 18.2401, 18.2401, 18.24011, 18.24011, 18.24012, 
    18.24013, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 
    18.2401, 18.24012, 18.24011, 18.24011, 18.2401, 18.24013, 18.24011, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.24011, 18.2401, 18.2401, 
    18.24012, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.2401, 18.24009, 18.24009, 18.24007, 18.24009, 
    18.24007, 18.24008, 18.24006, 18.24011, 18.24008, 18.24012, 18.24012, 
    18.24011, 18.24009, 18.2401, 18.24009, 18.24012, 18.24013, 18.24013, 
    18.24014, 18.24013, 18.24013, 18.24013, 18.24013, 18.24012, 18.24012, 
    18.2401, 18.24009, 18.24007, 18.24006, 18.24004, 18.24003, 18.24003, 
    18.24003 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976256e-05, 5.976241e-05, 5.976244e-05, 5.976232e-05, 5.976239e-05, 
    5.976231e-05, 5.976253e-05, 5.976241e-05, 5.976249e-05, 5.976254e-05, 
    5.976209e-05, 5.976231e-05, 5.976186e-05, 5.9762e-05, 5.976164e-05, 
    5.976188e-05, 5.976159e-05, 5.976165e-05, 5.976148e-05, 5.976153e-05, 
    5.976132e-05, 5.976146e-05, 5.976121e-05, 5.976135e-05, 5.976133e-05, 
    5.976146e-05, 5.976227e-05, 5.976212e-05, 5.976228e-05, 5.976226e-05, 
    5.976227e-05, 5.976238e-05, 5.976245e-05, 5.976257e-05, 5.976255e-05, 
    5.976246e-05, 5.976225e-05, 5.976232e-05, 5.976214e-05, 5.976214e-05, 
    5.976195e-05, 5.976203e-05, 5.97617e-05, 5.97618e-05, 5.976153e-05, 
    5.976159e-05, 5.976153e-05, 5.976155e-05, 5.976153e-05, 5.976163e-05, 
    5.976159e-05, 5.976167e-05, 5.976202e-05, 5.976192e-05, 5.976222e-05, 
    5.97624e-05, 5.976252e-05, 5.976261e-05, 5.97626e-05, 5.976257e-05, 
    5.976246e-05, 5.976234e-05, 5.976226e-05, 5.97622e-05, 5.976214e-05, 
    5.976198e-05, 5.976189e-05, 5.976169e-05, 5.976172e-05, 5.976166e-05, 
    5.97616e-05, 5.97615e-05, 5.976152e-05, 5.976148e-05, 5.976166e-05, 
    5.976154e-05, 5.976174e-05, 5.976169e-05, 5.976213e-05, 5.97623e-05, 
    5.976237e-05, 5.976243e-05, 5.976259e-05, 5.976248e-05, 5.976252e-05, 
    5.976242e-05, 5.976236e-05, 5.976239e-05, 5.97622e-05, 5.976227e-05, 
    5.976188e-05, 5.976205e-05, 5.976161e-05, 5.976171e-05, 5.976158e-05, 
    5.976165e-05, 5.976154e-05, 5.976164e-05, 5.976146e-05, 5.976142e-05, 
    5.976145e-05, 5.976135e-05, 5.976165e-05, 5.976153e-05, 5.976239e-05, 
    5.976239e-05, 5.976237e-05, 5.976247e-05, 5.976247e-05, 5.976257e-05, 
    5.976249e-05, 5.976245e-05, 5.976236e-05, 5.97623e-05, 5.976225e-05, 
    5.976214e-05, 5.976201e-05, 5.976183e-05, 5.976171e-05, 5.976162e-05, 
    5.976167e-05, 5.976163e-05, 5.976168e-05, 5.97617e-05, 5.976144e-05, 
    5.976159e-05, 5.976136e-05, 5.976137e-05, 5.976147e-05, 5.976137e-05, 
    5.976238e-05, 5.976241e-05, 5.976251e-05, 5.976243e-05, 5.976258e-05, 
    5.97625e-05, 5.976245e-05, 5.976227e-05, 5.976223e-05, 5.97622e-05, 
    5.976213e-05, 5.976203e-05, 5.976187e-05, 5.976173e-05, 5.97616e-05, 
    5.976161e-05, 5.976161e-05, 5.976158e-05, 5.976165e-05, 5.976157e-05, 
    5.976155e-05, 5.976159e-05, 5.976138e-05, 5.976143e-05, 5.976137e-05, 
    5.976141e-05, 5.976241e-05, 5.976235e-05, 5.976238e-05, 5.976233e-05, 
    5.976237e-05, 5.976221e-05, 5.976216e-05, 5.976194e-05, 5.976203e-05, 
    5.976189e-05, 5.976202e-05, 5.976199e-05, 5.976189e-05, 5.976201e-05, 
    5.976174e-05, 5.976192e-05, 5.976158e-05, 5.976176e-05, 5.976156e-05, 
    5.97616e-05, 5.976154e-05, 5.976149e-05, 5.976142e-05, 5.97613e-05, 
    5.976133e-05, 5.976122e-05, 5.976228e-05, 5.976222e-05, 5.976222e-05, 
    5.976215e-05, 5.976211e-05, 5.9762e-05, 5.976183e-05, 5.976189e-05, 
    5.976178e-05, 5.976175e-05, 5.976193e-05, 5.976182e-05, 5.976218e-05, 
    5.976212e-05, 5.976215e-05, 5.976227e-05, 5.976188e-05, 5.976208e-05, 
    5.976171e-05, 5.976182e-05, 5.976149e-05, 5.976165e-05, 5.976134e-05, 
    5.976121e-05, 5.976108e-05, 5.976093e-05, 5.976218e-05, 5.976223e-05, 
    5.976215e-05, 5.976204e-05, 5.976194e-05, 5.976181e-05, 5.976179e-05, 
    5.976177e-05, 5.976171e-05, 5.976165e-05, 5.976176e-05, 5.976164e-05, 
    5.97621e-05, 5.976186e-05, 5.976224e-05, 5.976213e-05, 5.976205e-05, 
    5.976208e-05, 5.97619e-05, 5.976186e-05, 5.976168e-05, 5.976177e-05, 
    5.976124e-05, 5.976147e-05, 5.976082e-05, 5.9761e-05, 5.976224e-05, 
    5.976218e-05, 5.976198e-05, 5.976207e-05, 5.97618e-05, 5.976173e-05, 
    5.976168e-05, 5.976161e-05, 5.97616e-05, 5.976156e-05, 5.976163e-05, 
    5.976156e-05, 5.976181e-05, 5.97617e-05, 5.9762e-05, 5.976193e-05, 
    5.976196e-05, 5.9762e-05, 5.976189e-05, 5.976176e-05, 5.976176e-05, 
    5.976172e-05, 5.976161e-05, 5.97618e-05, 5.976121e-05, 5.976157e-05, 
    5.976212e-05, 5.976201e-05, 5.976199e-05, 5.976203e-05, 5.976174e-05, 
    5.976185e-05, 5.976156e-05, 5.976163e-05, 5.976151e-05, 5.976157e-05, 
    5.976158e-05, 5.976166e-05, 5.976171e-05, 5.976184e-05, 5.976194e-05, 
    5.976203e-05, 5.976201e-05, 5.976192e-05, 5.976175e-05, 5.97616e-05, 
    5.976163e-05, 5.976152e-05, 5.976182e-05, 5.976169e-05, 5.976174e-05, 
    5.976162e-05, 5.97619e-05, 5.976166e-05, 5.976195e-05, 5.976193e-05, 
    5.976185e-05, 5.976169e-05, 5.976165e-05, 5.976161e-05, 5.976163e-05, 
    5.976175e-05, 5.976177e-05, 5.976185e-05, 5.976187e-05, 5.976194e-05, 
    5.976199e-05, 5.976194e-05, 5.976189e-05, 5.976175e-05, 5.976162e-05, 
    5.976149e-05, 5.976145e-05, 5.976129e-05, 5.976142e-05, 5.976121e-05, 
    5.976139e-05, 5.976107e-05, 5.976164e-05, 5.976139e-05, 5.976185e-05, 
    5.976179e-05, 5.976171e-05, 5.976151e-05, 5.976162e-05, 5.976149e-05, 
    5.976177e-05, 5.976191e-05, 5.976195e-05, 5.976202e-05, 5.976195e-05, 
    5.976196e-05, 5.976189e-05, 5.976191e-05, 5.976174e-05, 5.976183e-05, 
    5.976158e-05, 5.976149e-05, 5.976123e-05, 5.976107e-05, 5.976091e-05, 
    5.976084e-05, 5.976082e-05, 5.976081e-05 ;

 TOTLITC_1m =
  5.976256e-05, 5.976241e-05, 5.976244e-05, 5.976232e-05, 5.976239e-05, 
    5.976231e-05, 5.976253e-05, 5.976241e-05, 5.976249e-05, 5.976254e-05, 
    5.976209e-05, 5.976231e-05, 5.976186e-05, 5.9762e-05, 5.976164e-05, 
    5.976188e-05, 5.976159e-05, 5.976165e-05, 5.976148e-05, 5.976153e-05, 
    5.976132e-05, 5.976146e-05, 5.976121e-05, 5.976135e-05, 5.976133e-05, 
    5.976146e-05, 5.976227e-05, 5.976212e-05, 5.976228e-05, 5.976226e-05, 
    5.976227e-05, 5.976238e-05, 5.976245e-05, 5.976257e-05, 5.976255e-05, 
    5.976246e-05, 5.976225e-05, 5.976232e-05, 5.976214e-05, 5.976214e-05, 
    5.976195e-05, 5.976203e-05, 5.97617e-05, 5.97618e-05, 5.976153e-05, 
    5.976159e-05, 5.976153e-05, 5.976155e-05, 5.976153e-05, 5.976163e-05, 
    5.976159e-05, 5.976167e-05, 5.976202e-05, 5.976192e-05, 5.976222e-05, 
    5.97624e-05, 5.976252e-05, 5.976261e-05, 5.97626e-05, 5.976257e-05, 
    5.976246e-05, 5.976234e-05, 5.976226e-05, 5.97622e-05, 5.976214e-05, 
    5.976198e-05, 5.976189e-05, 5.976169e-05, 5.976172e-05, 5.976166e-05, 
    5.97616e-05, 5.97615e-05, 5.976152e-05, 5.976148e-05, 5.976166e-05, 
    5.976154e-05, 5.976174e-05, 5.976169e-05, 5.976213e-05, 5.97623e-05, 
    5.976237e-05, 5.976243e-05, 5.976259e-05, 5.976248e-05, 5.976252e-05, 
    5.976242e-05, 5.976236e-05, 5.976239e-05, 5.97622e-05, 5.976227e-05, 
    5.976188e-05, 5.976205e-05, 5.976161e-05, 5.976171e-05, 5.976158e-05, 
    5.976165e-05, 5.976154e-05, 5.976164e-05, 5.976146e-05, 5.976142e-05, 
    5.976145e-05, 5.976135e-05, 5.976165e-05, 5.976153e-05, 5.976239e-05, 
    5.976239e-05, 5.976237e-05, 5.976247e-05, 5.976247e-05, 5.976257e-05, 
    5.976249e-05, 5.976245e-05, 5.976236e-05, 5.97623e-05, 5.976225e-05, 
    5.976214e-05, 5.976201e-05, 5.976183e-05, 5.976171e-05, 5.976162e-05, 
    5.976167e-05, 5.976163e-05, 5.976168e-05, 5.97617e-05, 5.976144e-05, 
    5.976159e-05, 5.976136e-05, 5.976137e-05, 5.976147e-05, 5.976137e-05, 
    5.976238e-05, 5.976241e-05, 5.976251e-05, 5.976243e-05, 5.976258e-05, 
    5.97625e-05, 5.976245e-05, 5.976227e-05, 5.976223e-05, 5.97622e-05, 
    5.976213e-05, 5.976203e-05, 5.976187e-05, 5.976173e-05, 5.97616e-05, 
    5.976161e-05, 5.976161e-05, 5.976158e-05, 5.976165e-05, 5.976157e-05, 
    5.976155e-05, 5.976159e-05, 5.976138e-05, 5.976143e-05, 5.976137e-05, 
    5.976141e-05, 5.976241e-05, 5.976235e-05, 5.976238e-05, 5.976233e-05, 
    5.976237e-05, 5.976221e-05, 5.976216e-05, 5.976194e-05, 5.976203e-05, 
    5.976189e-05, 5.976202e-05, 5.976199e-05, 5.976189e-05, 5.976201e-05, 
    5.976174e-05, 5.976192e-05, 5.976158e-05, 5.976176e-05, 5.976156e-05, 
    5.97616e-05, 5.976154e-05, 5.976149e-05, 5.976142e-05, 5.97613e-05, 
    5.976133e-05, 5.976122e-05, 5.976228e-05, 5.976222e-05, 5.976222e-05, 
    5.976215e-05, 5.976211e-05, 5.9762e-05, 5.976183e-05, 5.976189e-05, 
    5.976178e-05, 5.976175e-05, 5.976193e-05, 5.976182e-05, 5.976218e-05, 
    5.976212e-05, 5.976215e-05, 5.976227e-05, 5.976188e-05, 5.976208e-05, 
    5.976171e-05, 5.976182e-05, 5.976149e-05, 5.976165e-05, 5.976134e-05, 
    5.976121e-05, 5.976108e-05, 5.976093e-05, 5.976218e-05, 5.976223e-05, 
    5.976215e-05, 5.976204e-05, 5.976194e-05, 5.976181e-05, 5.976179e-05, 
    5.976177e-05, 5.976171e-05, 5.976165e-05, 5.976176e-05, 5.976164e-05, 
    5.97621e-05, 5.976186e-05, 5.976224e-05, 5.976213e-05, 5.976205e-05, 
    5.976208e-05, 5.97619e-05, 5.976186e-05, 5.976168e-05, 5.976177e-05, 
    5.976124e-05, 5.976147e-05, 5.976082e-05, 5.9761e-05, 5.976224e-05, 
    5.976218e-05, 5.976198e-05, 5.976207e-05, 5.97618e-05, 5.976173e-05, 
    5.976168e-05, 5.976161e-05, 5.97616e-05, 5.976156e-05, 5.976163e-05, 
    5.976156e-05, 5.976181e-05, 5.97617e-05, 5.9762e-05, 5.976193e-05, 
    5.976196e-05, 5.9762e-05, 5.976189e-05, 5.976176e-05, 5.976176e-05, 
    5.976172e-05, 5.976161e-05, 5.97618e-05, 5.976121e-05, 5.976157e-05, 
    5.976212e-05, 5.976201e-05, 5.976199e-05, 5.976203e-05, 5.976174e-05, 
    5.976185e-05, 5.976156e-05, 5.976163e-05, 5.976151e-05, 5.976157e-05, 
    5.976158e-05, 5.976166e-05, 5.976171e-05, 5.976184e-05, 5.976194e-05, 
    5.976203e-05, 5.976201e-05, 5.976192e-05, 5.976175e-05, 5.97616e-05, 
    5.976163e-05, 5.976152e-05, 5.976182e-05, 5.976169e-05, 5.976174e-05, 
    5.976162e-05, 5.97619e-05, 5.976166e-05, 5.976195e-05, 5.976193e-05, 
    5.976185e-05, 5.976169e-05, 5.976165e-05, 5.976161e-05, 5.976163e-05, 
    5.976175e-05, 5.976177e-05, 5.976185e-05, 5.976187e-05, 5.976194e-05, 
    5.976199e-05, 5.976194e-05, 5.976189e-05, 5.976175e-05, 5.976162e-05, 
    5.976149e-05, 5.976145e-05, 5.976129e-05, 5.976142e-05, 5.976121e-05, 
    5.976139e-05, 5.976107e-05, 5.976164e-05, 5.976139e-05, 5.976185e-05, 
    5.976179e-05, 5.976171e-05, 5.976151e-05, 5.976162e-05, 5.976149e-05, 
    5.976177e-05, 5.976191e-05, 5.976195e-05, 5.976202e-05, 5.976195e-05, 
    5.976196e-05, 5.976189e-05, 5.976191e-05, 5.976174e-05, 5.976183e-05, 
    5.976158e-05, 5.976149e-05, 5.976123e-05, 5.976107e-05, 5.976091e-05, 
    5.976084e-05, 5.976082e-05, 5.976081e-05 ;

 TOTLITN =
  1.375944e-06, 1.37594e-06, 1.375941e-06, 1.375937e-06, 1.375939e-06, 
    1.375937e-06, 1.375943e-06, 1.37594e-06, 1.375942e-06, 1.375943e-06, 
    1.375931e-06, 1.375937e-06, 1.375924e-06, 1.375928e-06, 1.375918e-06, 
    1.375925e-06, 1.375917e-06, 1.375918e-06, 1.375914e-06, 1.375915e-06, 
    1.375909e-06, 1.375913e-06, 1.375906e-06, 1.37591e-06, 1.375909e-06, 
    1.375913e-06, 1.375936e-06, 1.375931e-06, 1.375936e-06, 1.375935e-06, 
    1.375936e-06, 1.375939e-06, 1.375941e-06, 1.375944e-06, 1.375944e-06, 
    1.375941e-06, 1.375935e-06, 1.375937e-06, 1.375932e-06, 1.375932e-06, 
    1.375927e-06, 1.375929e-06, 1.37592e-06, 1.375922e-06, 1.375915e-06, 
    1.375917e-06, 1.375915e-06, 1.375916e-06, 1.375915e-06, 1.375918e-06, 
    1.375917e-06, 1.375919e-06, 1.375929e-06, 1.375926e-06, 1.375934e-06, 
    1.37594e-06, 1.375943e-06, 1.375945e-06, 1.375945e-06, 1.375944e-06, 
    1.375941e-06, 1.375938e-06, 1.375935e-06, 1.375934e-06, 1.375932e-06, 
    1.375927e-06, 1.375925e-06, 1.375919e-06, 1.37592e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375915e-06, 1.375913e-06, 1.375919e-06, 
    1.375915e-06, 1.375921e-06, 1.375919e-06, 1.375932e-06, 1.375937e-06, 
    1.375939e-06, 1.37594e-06, 1.375945e-06, 1.375942e-06, 1.375943e-06, 
    1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375934e-06, 1.375936e-06, 
    1.375925e-06, 1.37593e-06, 1.375917e-06, 1.37592e-06, 1.375916e-06, 
    1.375918e-06, 1.375915e-06, 1.375918e-06, 1.375913e-06, 1.375912e-06, 
    1.375913e-06, 1.37591e-06, 1.375918e-06, 1.375915e-06, 1.375939e-06, 
    1.375939e-06, 1.375938e-06, 1.375941e-06, 1.375942e-06, 1.375944e-06, 
    1.375942e-06, 1.375941e-06, 1.375938e-06, 1.375937e-06, 1.375935e-06, 
    1.375932e-06, 1.375928e-06, 1.375923e-06, 1.37592e-06, 1.375918e-06, 
    1.375919e-06, 1.375918e-06, 1.375919e-06, 1.37592e-06, 1.375912e-06, 
    1.375917e-06, 1.37591e-06, 1.375911e-06, 1.375913e-06, 1.375911e-06, 
    1.375939e-06, 1.37594e-06, 1.375943e-06, 1.37594e-06, 1.375945e-06, 
    1.375942e-06, 1.375941e-06, 1.375936e-06, 1.375935e-06, 1.375934e-06, 
    1.375932e-06, 1.375929e-06, 1.375925e-06, 1.375921e-06, 1.375917e-06, 
    1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 1.375916e-06, 
    1.375916e-06, 1.375917e-06, 1.375911e-06, 1.375912e-06, 1.375911e-06, 
    1.375912e-06, 1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375937e-06, 
    1.375938e-06, 1.375934e-06, 1.375933e-06, 1.375927e-06, 1.375929e-06, 
    1.375925e-06, 1.375929e-06, 1.375928e-06, 1.375925e-06, 1.375928e-06, 
    1.375921e-06, 1.375926e-06, 1.375916e-06, 1.375921e-06, 1.375916e-06, 
    1.375917e-06, 1.375915e-06, 1.375914e-06, 1.375912e-06, 1.375908e-06, 
    1.375909e-06, 1.375906e-06, 1.375936e-06, 1.375934e-06, 1.375934e-06, 
    1.375933e-06, 1.375931e-06, 1.375928e-06, 1.375923e-06, 1.375925e-06, 
    1.375922e-06, 1.375921e-06, 1.375926e-06, 1.375923e-06, 1.375933e-06, 
    1.375931e-06, 1.375932e-06, 1.375936e-06, 1.375925e-06, 1.375931e-06, 
    1.37592e-06, 1.375923e-06, 1.375914e-06, 1.375918e-06, 1.37591e-06, 
    1.375906e-06, 1.375902e-06, 1.375898e-06, 1.375933e-06, 1.375935e-06, 
    1.375932e-06, 1.375929e-06, 1.375927e-06, 1.375923e-06, 1.375922e-06, 
    1.375922e-06, 1.37592e-06, 1.375918e-06, 1.375921e-06, 1.375918e-06, 
    1.375931e-06, 1.375924e-06, 1.375935e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.375925e-06, 1.375924e-06, 1.375919e-06, 1.375922e-06, 
    1.375907e-06, 1.375913e-06, 1.375895e-06, 1.3759e-06, 1.375935e-06, 
    1.375933e-06, 1.375928e-06, 1.37593e-06, 1.375923e-06, 1.375921e-06, 
    1.375919e-06, 1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 
    1.375916e-06, 1.375923e-06, 1.37592e-06, 1.375928e-06, 1.375926e-06, 
    1.375927e-06, 1.375928e-06, 1.375925e-06, 1.375921e-06, 1.375921e-06, 
    1.37592e-06, 1.375917e-06, 1.375922e-06, 1.375906e-06, 1.375916e-06, 
    1.375932e-06, 1.375928e-06, 1.375928e-06, 1.375929e-06, 1.375921e-06, 
    1.375924e-06, 1.375916e-06, 1.375918e-06, 1.375914e-06, 1.375916e-06, 
    1.375916e-06, 1.375919e-06, 1.37592e-06, 1.375924e-06, 1.375927e-06, 
    1.375929e-06, 1.375928e-06, 1.375926e-06, 1.375921e-06, 1.375917e-06, 
    1.375918e-06, 1.375915e-06, 1.375923e-06, 1.37592e-06, 1.375921e-06, 
    1.375917e-06, 1.375925e-06, 1.375918e-06, 1.375927e-06, 1.375926e-06, 
    1.375924e-06, 1.375919e-06, 1.375918e-06, 1.375917e-06, 1.375918e-06, 
    1.375921e-06, 1.375922e-06, 1.375924e-06, 1.375925e-06, 1.375926e-06, 
    1.375928e-06, 1.375926e-06, 1.375925e-06, 1.375921e-06, 1.375918e-06, 
    1.375914e-06, 1.375913e-06, 1.375908e-06, 1.375912e-06, 1.375906e-06, 
    1.375911e-06, 1.375902e-06, 1.375918e-06, 1.375911e-06, 1.375924e-06, 
    1.375922e-06, 1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375914e-06, 
    1.375922e-06, 1.375926e-06, 1.375927e-06, 1.375929e-06, 1.375927e-06, 
    1.375927e-06, 1.375925e-06, 1.375926e-06, 1.375921e-06, 1.375923e-06, 
    1.375916e-06, 1.375914e-06, 1.375907e-06, 1.375902e-06, 1.375898e-06, 
    1.375896e-06, 1.375895e-06, 1.375895e-06 ;

 TOTLITN_1m =
  1.375944e-06, 1.37594e-06, 1.375941e-06, 1.375937e-06, 1.375939e-06, 
    1.375937e-06, 1.375943e-06, 1.37594e-06, 1.375942e-06, 1.375943e-06, 
    1.375931e-06, 1.375937e-06, 1.375924e-06, 1.375928e-06, 1.375918e-06, 
    1.375925e-06, 1.375917e-06, 1.375918e-06, 1.375914e-06, 1.375915e-06, 
    1.375909e-06, 1.375913e-06, 1.375906e-06, 1.37591e-06, 1.375909e-06, 
    1.375913e-06, 1.375936e-06, 1.375931e-06, 1.375936e-06, 1.375935e-06, 
    1.375936e-06, 1.375939e-06, 1.375941e-06, 1.375944e-06, 1.375944e-06, 
    1.375941e-06, 1.375935e-06, 1.375937e-06, 1.375932e-06, 1.375932e-06, 
    1.375927e-06, 1.375929e-06, 1.37592e-06, 1.375922e-06, 1.375915e-06, 
    1.375917e-06, 1.375915e-06, 1.375916e-06, 1.375915e-06, 1.375918e-06, 
    1.375917e-06, 1.375919e-06, 1.375929e-06, 1.375926e-06, 1.375934e-06, 
    1.37594e-06, 1.375943e-06, 1.375945e-06, 1.375945e-06, 1.375944e-06, 
    1.375941e-06, 1.375938e-06, 1.375935e-06, 1.375934e-06, 1.375932e-06, 
    1.375927e-06, 1.375925e-06, 1.375919e-06, 1.37592e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375915e-06, 1.375913e-06, 1.375919e-06, 
    1.375915e-06, 1.375921e-06, 1.375919e-06, 1.375932e-06, 1.375937e-06, 
    1.375939e-06, 1.37594e-06, 1.375945e-06, 1.375942e-06, 1.375943e-06, 
    1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375934e-06, 1.375936e-06, 
    1.375925e-06, 1.37593e-06, 1.375917e-06, 1.37592e-06, 1.375916e-06, 
    1.375918e-06, 1.375915e-06, 1.375918e-06, 1.375913e-06, 1.375912e-06, 
    1.375913e-06, 1.37591e-06, 1.375918e-06, 1.375915e-06, 1.375939e-06, 
    1.375939e-06, 1.375938e-06, 1.375941e-06, 1.375942e-06, 1.375944e-06, 
    1.375942e-06, 1.375941e-06, 1.375938e-06, 1.375937e-06, 1.375935e-06, 
    1.375932e-06, 1.375928e-06, 1.375923e-06, 1.37592e-06, 1.375918e-06, 
    1.375919e-06, 1.375918e-06, 1.375919e-06, 1.37592e-06, 1.375912e-06, 
    1.375917e-06, 1.37591e-06, 1.375911e-06, 1.375913e-06, 1.375911e-06, 
    1.375939e-06, 1.37594e-06, 1.375943e-06, 1.37594e-06, 1.375945e-06, 
    1.375942e-06, 1.375941e-06, 1.375936e-06, 1.375935e-06, 1.375934e-06, 
    1.375932e-06, 1.375929e-06, 1.375925e-06, 1.375921e-06, 1.375917e-06, 
    1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 1.375916e-06, 
    1.375916e-06, 1.375917e-06, 1.375911e-06, 1.375912e-06, 1.375911e-06, 
    1.375912e-06, 1.37594e-06, 1.375938e-06, 1.375939e-06, 1.375937e-06, 
    1.375938e-06, 1.375934e-06, 1.375933e-06, 1.375927e-06, 1.375929e-06, 
    1.375925e-06, 1.375929e-06, 1.375928e-06, 1.375925e-06, 1.375928e-06, 
    1.375921e-06, 1.375926e-06, 1.375916e-06, 1.375921e-06, 1.375916e-06, 
    1.375917e-06, 1.375915e-06, 1.375914e-06, 1.375912e-06, 1.375908e-06, 
    1.375909e-06, 1.375906e-06, 1.375936e-06, 1.375934e-06, 1.375934e-06, 
    1.375933e-06, 1.375931e-06, 1.375928e-06, 1.375923e-06, 1.375925e-06, 
    1.375922e-06, 1.375921e-06, 1.375926e-06, 1.375923e-06, 1.375933e-06, 
    1.375931e-06, 1.375932e-06, 1.375936e-06, 1.375925e-06, 1.375931e-06, 
    1.37592e-06, 1.375923e-06, 1.375914e-06, 1.375918e-06, 1.37591e-06, 
    1.375906e-06, 1.375902e-06, 1.375898e-06, 1.375933e-06, 1.375935e-06, 
    1.375932e-06, 1.375929e-06, 1.375927e-06, 1.375923e-06, 1.375922e-06, 
    1.375922e-06, 1.37592e-06, 1.375918e-06, 1.375921e-06, 1.375918e-06, 
    1.375931e-06, 1.375924e-06, 1.375935e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.375925e-06, 1.375924e-06, 1.375919e-06, 1.375922e-06, 
    1.375907e-06, 1.375913e-06, 1.375895e-06, 1.3759e-06, 1.375935e-06, 
    1.375933e-06, 1.375928e-06, 1.37593e-06, 1.375923e-06, 1.375921e-06, 
    1.375919e-06, 1.375917e-06, 1.375917e-06, 1.375916e-06, 1.375918e-06, 
    1.375916e-06, 1.375923e-06, 1.37592e-06, 1.375928e-06, 1.375926e-06, 
    1.375927e-06, 1.375928e-06, 1.375925e-06, 1.375921e-06, 1.375921e-06, 
    1.37592e-06, 1.375917e-06, 1.375922e-06, 1.375906e-06, 1.375916e-06, 
    1.375932e-06, 1.375928e-06, 1.375928e-06, 1.375929e-06, 1.375921e-06, 
    1.375924e-06, 1.375916e-06, 1.375918e-06, 1.375914e-06, 1.375916e-06, 
    1.375916e-06, 1.375919e-06, 1.37592e-06, 1.375924e-06, 1.375927e-06, 
    1.375929e-06, 1.375928e-06, 1.375926e-06, 1.375921e-06, 1.375917e-06, 
    1.375918e-06, 1.375915e-06, 1.375923e-06, 1.37592e-06, 1.375921e-06, 
    1.375917e-06, 1.375925e-06, 1.375918e-06, 1.375927e-06, 1.375926e-06, 
    1.375924e-06, 1.375919e-06, 1.375918e-06, 1.375917e-06, 1.375918e-06, 
    1.375921e-06, 1.375922e-06, 1.375924e-06, 1.375925e-06, 1.375926e-06, 
    1.375928e-06, 1.375926e-06, 1.375925e-06, 1.375921e-06, 1.375918e-06, 
    1.375914e-06, 1.375913e-06, 1.375908e-06, 1.375912e-06, 1.375906e-06, 
    1.375911e-06, 1.375902e-06, 1.375918e-06, 1.375911e-06, 1.375924e-06, 
    1.375922e-06, 1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375914e-06, 
    1.375922e-06, 1.375926e-06, 1.375927e-06, 1.375929e-06, 1.375927e-06, 
    1.375927e-06, 1.375925e-06, 1.375926e-06, 1.375921e-06, 1.375923e-06, 
    1.375916e-06, 1.375914e-06, 1.375907e-06, 1.375902e-06, 1.375898e-06, 
    1.375896e-06, 1.375895e-06, 1.375895e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34481, 17.34479, 17.3448, 17.34479, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.34481, 17.34476, 17.34479, 17.34474, 17.34476, 
    17.34472, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34471, 17.34472, 17.34471, 17.34473, 17.34472, 17.34473, 
    17.34473, 17.34477, 17.34478, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.3448, 17.3448, 17.34479, 17.34479, 17.34477, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34472, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.3448, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.3447, 17.34471, 17.34479, 17.34479, 17.34479, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34475, 17.34476, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34476, 17.34473, 17.34475, 17.34472, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 17.3447, 17.34469, 
    17.34478, 17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 
    17.34475, 17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 
    17.34477, 17.34478, 17.34475, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34473, 17.3447, 17.34469, 17.34468, 17.34466, 17.34477, 17.34478, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34474, 17.34473, 
    17.34473, 17.34474, 17.34472, 17.34477, 17.34475, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 
    17.34471, 17.34465, 17.34467, 17.34478, 17.34477, 17.34476, 17.34476, 
    17.34474, 17.34473, 17.34473, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34474, 17.34473, 17.34476, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 
    17.34472, 17.34477, 17.34476, 17.34476, 17.34476, 17.34473, 17.34474, 
    17.34472, 17.34472, 17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34474, 17.34473, 17.34473, 17.34472, 17.34475, 
    17.34473, 17.34475, 17.34475, 17.34474, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34469, 17.3447, 17.34468, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34474, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34475, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 TOTSOMC_1m =
  17.34481, 17.34479, 17.3448, 17.34479, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.34481, 17.34476, 17.34479, 17.34474, 17.34476, 
    17.34472, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34471, 17.34472, 17.34471, 17.34473, 17.34472, 17.34473, 
    17.34473, 17.34477, 17.34478, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.3448, 17.3448, 17.34479, 17.34479, 17.34477, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34472, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.3448, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 
    17.3447, 17.34471, 17.34479, 17.34479, 17.34479, 17.34479, 17.34479, 
    17.34478, 17.34477, 17.34475, 17.34476, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34476, 17.34473, 17.34475, 17.34472, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 17.3447, 17.34469, 
    17.34478, 17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 
    17.34475, 17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 
    17.34477, 17.34478, 17.34475, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34473, 17.3447, 17.34469, 17.34468, 17.34466, 17.34477, 17.34478, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34474, 17.34473, 
    17.34473, 17.34474, 17.34472, 17.34477, 17.34475, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 
    17.34471, 17.34465, 17.34467, 17.34478, 17.34477, 17.34476, 17.34476, 
    17.34474, 17.34473, 17.34473, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34474, 17.34473, 17.34476, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 
    17.34472, 17.34477, 17.34476, 17.34476, 17.34476, 17.34473, 17.34474, 
    17.34472, 17.34472, 17.34471, 17.34472, 17.34472, 17.34473, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 
    17.34472, 17.34472, 17.34474, 17.34473, 17.34473, 17.34472, 17.34475, 
    17.34473, 17.34475, 17.34475, 17.34474, 17.34473, 17.34473, 17.34472, 
    17.34472, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 17.34476, 
    17.34475, 17.34475, 17.34473, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34469, 17.3447, 17.34468, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34474, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34475, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 TOTSOMN =
  1.773786, 1.773784, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773784, 1.773785, 1.773786, 1.77378, 1.773783, 1.773777, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773773, 1.773771, 
    1.773772, 1.773769, 1.773771, 1.773771, 1.773772, 1.773782, 1.773781, 
    1.773783, 1.773782, 1.773782, 1.773784, 1.773785, 1.773786, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773778, 1.77378, 
    1.773775, 1.773777, 1.773773, 1.773774, 1.773773, 1.773773, 1.773773, 
    1.773775, 1.773774, 1.773775, 1.773779, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.773775, 1.773773, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773786, 1.773785, 
    1.773786, 1.773784, 1.773784, 1.773784, 1.773782, 1.773782, 1.773778, 
    1.77378, 1.773774, 1.773775, 1.773774, 1.773775, 1.773773, 1.773775, 
    1.773772, 1.773772, 1.773772, 1.773771, 1.773775, 1.773773, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773786, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773782, 1.773781, 1.773779, 1.773777, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773775, 1.773775, 1.773772, 1.773774, 
    1.773771, 1.773771, 1.773772, 1.773771, 1.773784, 1.773784, 1.773786, 
    1.773785, 1.773786, 1.773785, 1.773785, 1.773782, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773777, 1.773776, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773775, 1.773774, 1.773773, 1.773774, 1.773771, 1.773772, 
    1.773771, 1.773772, 1.773784, 1.773784, 1.773784, 1.773783, 1.773784, 
    1.773782, 1.773781, 1.773778, 1.77378, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773779, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.77377, 1.773771, 1.773769, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.77378, 1.773779, 1.773777, 
    1.773778, 1.773776, 1.773776, 1.773778, 1.773777, 1.773781, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773775, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773767, 1.773766, 1.773781, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773777, 1.773777, 1.773776, 1.773775, 
    1.773775, 1.773776, 1.773775, 1.77378, 1.773777, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773777, 1.773775, 1.773776, 1.773769, 
    1.773772, 1.773764, 1.773767, 1.773782, 1.773781, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773777, 1.773775, 1.773779, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773774, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.773779, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773775, 
    1.773777, 1.773778, 1.77378, 1.773779, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773775, 1.773776, 1.773774, 1.773778, 
    1.773775, 1.773779, 1.773778, 1.773777, 1.773775, 1.773775, 1.773774, 
    1.773775, 1.773776, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 
    1.773778, 1.773778, 1.773776, 1.773774, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773771, 1.773767, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773775, 1.773773, 1.773774, 1.773773, 1.773776, 1.773778, 
    1.773779, 1.773779, 1.773778, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.773769, 1.773767, 1.773765, 1.773764, 
    1.773764, 1.773764 ;

 TOTSOMN_1m =
  1.773786, 1.773784, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773784, 1.773785, 1.773786, 1.77378, 1.773783, 1.773777, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773773, 1.773771, 
    1.773772, 1.773769, 1.773771, 1.773771, 1.773772, 1.773782, 1.773781, 
    1.773783, 1.773782, 1.773782, 1.773784, 1.773785, 1.773786, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773778, 1.77378, 
    1.773775, 1.773777, 1.773773, 1.773774, 1.773773, 1.773773, 1.773773, 
    1.773775, 1.773774, 1.773775, 1.773779, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.773775, 1.773773, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773786, 1.773785, 
    1.773786, 1.773784, 1.773784, 1.773784, 1.773782, 1.773782, 1.773778, 
    1.77378, 1.773774, 1.773775, 1.773774, 1.773775, 1.773773, 1.773775, 
    1.773772, 1.773772, 1.773772, 1.773771, 1.773775, 1.773773, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773786, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773782, 1.773781, 1.773779, 1.773777, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773775, 1.773775, 1.773772, 1.773774, 
    1.773771, 1.773771, 1.773772, 1.773771, 1.773784, 1.773784, 1.773786, 
    1.773785, 1.773786, 1.773785, 1.773785, 1.773782, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773777, 1.773776, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773775, 1.773774, 1.773773, 1.773774, 1.773771, 1.773772, 
    1.773771, 1.773772, 1.773784, 1.773784, 1.773784, 1.773783, 1.773784, 
    1.773782, 1.773781, 1.773778, 1.77378, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773779, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773773, 1.773773, 1.773772, 1.77377, 1.773771, 1.773769, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.77378, 1.773779, 1.773777, 
    1.773778, 1.773776, 1.773776, 1.773778, 1.773777, 1.773781, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773775, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773767, 1.773766, 1.773781, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773777, 1.773777, 1.773776, 1.773775, 
    1.773775, 1.773776, 1.773775, 1.77378, 1.773777, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773777, 1.773775, 1.773776, 1.773769, 
    1.773772, 1.773764, 1.773767, 1.773782, 1.773781, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773774, 1.773777, 1.773775, 1.773779, 1.773778, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773774, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.773779, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773775, 
    1.773777, 1.773778, 1.77378, 1.773779, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773775, 1.773776, 1.773774, 1.773778, 
    1.773775, 1.773779, 1.773778, 1.773777, 1.773775, 1.773775, 1.773774, 
    1.773775, 1.773776, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 
    1.773778, 1.773778, 1.773776, 1.773774, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773771, 1.773767, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773775, 1.773773, 1.773774, 1.773773, 1.773776, 1.773778, 
    1.773779, 1.773779, 1.773778, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.773769, 1.773767, 1.773765, 1.773764, 
    1.773764, 1.773764 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9696, 249.9699, 249.9698, 249.9701, 249.9699, 249.9701, 249.9697, 
    249.9699, 249.9698, 249.9697, 249.9704, 249.9701, 249.9709, 249.9706, 
    249.9713, 249.9708, 249.9713, 249.9713, 249.9715, 249.9715, 249.9718, 
    249.9716, 249.972, 249.9718, 249.9718, 249.9716, 249.9702, 249.9704, 
    249.9701, 249.9702, 249.9702, 249.9699, 249.9698, 249.9696, 249.9697, 
    249.9698, 249.9702, 249.9701, 249.9704, 249.9704, 249.9707, 249.9706, 
    249.9711, 249.971, 249.9715, 249.9713, 249.9715, 249.9714, 249.9715, 
    249.9713, 249.9714, 249.9712, 249.9706, 249.9708, 249.9702, 249.9699, 
    249.9697, 249.9696, 249.9696, 249.9696, 249.9698, 249.97, 249.9702, 
    249.9703, 249.9704, 249.9707, 249.9708, 249.9712, 249.9711, 249.9712, 
    249.9713, 249.9715, 249.9715, 249.9716, 249.9712, 249.9714, 249.9711, 
    249.9712, 249.9704, 249.9701, 249.97, 249.9699, 249.9696, 249.9698, 
    249.9697, 249.9699, 249.97, 249.9699, 249.9703, 249.9701, 249.9708, 
    249.9705, 249.9713, 249.9711, 249.9714, 249.9713, 249.9715, 249.9713, 
    249.9716, 249.9716, 249.9716, 249.9718, 249.9713, 249.9715, 249.9699, 
    249.9699, 249.97, 249.9698, 249.9698, 249.9696, 249.9698, 249.9698, 
    249.97, 249.9701, 249.9702, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9713, 249.9712, 249.9713, 249.9712, 249.9711, 249.9716, 249.9714, 
    249.9718, 249.9717, 249.9716, 249.9717, 249.9699, 249.9699, 249.9697, 
    249.9699, 249.9696, 249.9697, 249.9698, 249.9701, 249.9702, 249.9703, 
    249.9704, 249.9706, 249.9709, 249.9711, 249.9713, 249.9713, 249.9713, 
    249.9714, 249.9713, 249.9714, 249.9714, 249.9714, 249.9717, 249.9716, 
    249.9717, 249.9717, 249.9699, 249.97, 249.97, 249.97, 249.97, 249.9702, 
    249.9703, 249.9707, 249.9706, 249.9708, 249.9706, 249.9706, 249.9708, 
    249.9706, 249.9711, 249.9707, 249.9714, 249.971, 249.9714, 249.9713, 
    249.9715, 249.9715, 249.9717, 249.9719, 249.9718, 249.972, 249.9701, 
    249.9702, 249.9702, 249.9704, 249.9704, 249.9706, 249.9709, 249.9708, 
    249.971, 249.9711, 249.9707, 249.9709, 249.9703, 249.9704, 249.9704, 
    249.9701, 249.9708, 249.9705, 249.9711, 249.9709, 249.9715, 249.9712, 
    249.9718, 249.972, 249.9723, 249.9725, 249.9703, 249.9702, 249.9704, 
    249.9706, 249.9707, 249.971, 249.971, 249.971, 249.9711, 249.9712, 
    249.971, 249.9713, 249.9704, 249.9709, 249.9702, 249.9704, 249.9705, 
    249.9705, 249.9708, 249.9709, 249.9712, 249.971, 249.972, 249.9716, 
    249.9727, 249.9724, 249.9702, 249.9703, 249.9707, 249.9705, 249.971, 
    249.9711, 249.9712, 249.9713, 249.9713, 249.9714, 249.9713, 249.9714, 
    249.971, 249.9712, 249.9706, 249.9707, 249.9707, 249.9706, 249.9708, 
    249.971, 249.9711, 249.9711, 249.9713, 249.971, 249.972, 249.9714, 
    249.9704, 249.9706, 249.9706, 249.9706, 249.9711, 249.9709, 249.9714, 
    249.9713, 249.9715, 249.9714, 249.9714, 249.9712, 249.9711, 249.9709, 
    249.9707, 249.9706, 249.9706, 249.9708, 249.9711, 249.9713, 249.9713, 
    249.9715, 249.9709, 249.9712, 249.9711, 249.9713, 249.9708, 249.9712, 
    249.9707, 249.9707, 249.9709, 249.9712, 249.9713, 249.9713, 249.9713, 
    249.9711, 249.971, 249.9709, 249.9709, 249.9707, 249.9707, 249.9707, 
    249.9708, 249.9711, 249.9713, 249.9715, 249.9716, 249.9719, 249.9716, 
    249.972, 249.9717, 249.9723, 249.9713, 249.9717, 249.9709, 249.971, 
    249.9711, 249.9715, 249.9713, 249.9715, 249.971, 249.9708, 249.9707, 
    249.9706, 249.9707, 249.9707, 249.9708, 249.9708, 249.9711, 249.9709, 
    249.9714, 249.9715, 249.972, 249.9723, 249.9726, 249.9727, 249.9727, 
    249.9727 ;

 TREFMNAV_R =
  249.9696, 249.9699, 249.9698, 249.9701, 249.9699, 249.9701, 249.9697, 
    249.9699, 249.9698, 249.9697, 249.9704, 249.9701, 249.9709, 249.9706, 
    249.9713, 249.9708, 249.9713, 249.9713, 249.9715, 249.9715, 249.9718, 
    249.9716, 249.972, 249.9718, 249.9718, 249.9716, 249.9702, 249.9704, 
    249.9701, 249.9702, 249.9702, 249.9699, 249.9698, 249.9696, 249.9697, 
    249.9698, 249.9702, 249.9701, 249.9704, 249.9704, 249.9707, 249.9706, 
    249.9711, 249.971, 249.9715, 249.9713, 249.9715, 249.9714, 249.9715, 
    249.9713, 249.9714, 249.9712, 249.9706, 249.9708, 249.9702, 249.9699, 
    249.9697, 249.9696, 249.9696, 249.9696, 249.9698, 249.97, 249.9702, 
    249.9703, 249.9704, 249.9707, 249.9708, 249.9712, 249.9711, 249.9712, 
    249.9713, 249.9715, 249.9715, 249.9716, 249.9712, 249.9714, 249.9711, 
    249.9712, 249.9704, 249.9701, 249.97, 249.9699, 249.9696, 249.9698, 
    249.9697, 249.9699, 249.97, 249.9699, 249.9703, 249.9701, 249.9708, 
    249.9705, 249.9713, 249.9711, 249.9714, 249.9713, 249.9715, 249.9713, 
    249.9716, 249.9716, 249.9716, 249.9718, 249.9713, 249.9715, 249.9699, 
    249.9699, 249.97, 249.9698, 249.9698, 249.9696, 249.9698, 249.9698, 
    249.97, 249.9701, 249.9702, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9713, 249.9712, 249.9713, 249.9712, 249.9711, 249.9716, 249.9714, 
    249.9718, 249.9717, 249.9716, 249.9717, 249.9699, 249.9699, 249.9697, 
    249.9699, 249.9696, 249.9697, 249.9698, 249.9701, 249.9702, 249.9703, 
    249.9704, 249.9706, 249.9709, 249.9711, 249.9713, 249.9713, 249.9713, 
    249.9714, 249.9713, 249.9714, 249.9714, 249.9714, 249.9717, 249.9716, 
    249.9717, 249.9717, 249.9699, 249.97, 249.97, 249.97, 249.97, 249.9702, 
    249.9703, 249.9707, 249.9706, 249.9708, 249.9706, 249.9706, 249.9708, 
    249.9706, 249.9711, 249.9707, 249.9714, 249.971, 249.9714, 249.9713, 
    249.9715, 249.9715, 249.9717, 249.9719, 249.9718, 249.972, 249.9701, 
    249.9702, 249.9702, 249.9704, 249.9704, 249.9706, 249.9709, 249.9708, 
    249.971, 249.9711, 249.9707, 249.9709, 249.9703, 249.9704, 249.9704, 
    249.9701, 249.9708, 249.9705, 249.9711, 249.9709, 249.9715, 249.9712, 
    249.9718, 249.972, 249.9723, 249.9725, 249.9703, 249.9702, 249.9704, 
    249.9706, 249.9707, 249.971, 249.971, 249.971, 249.9711, 249.9712, 
    249.971, 249.9713, 249.9704, 249.9709, 249.9702, 249.9704, 249.9705, 
    249.9705, 249.9708, 249.9709, 249.9712, 249.971, 249.972, 249.9716, 
    249.9727, 249.9724, 249.9702, 249.9703, 249.9707, 249.9705, 249.971, 
    249.9711, 249.9712, 249.9713, 249.9713, 249.9714, 249.9713, 249.9714, 
    249.971, 249.9712, 249.9706, 249.9707, 249.9707, 249.9706, 249.9708, 
    249.971, 249.9711, 249.9711, 249.9713, 249.971, 249.972, 249.9714, 
    249.9704, 249.9706, 249.9706, 249.9706, 249.9711, 249.9709, 249.9714, 
    249.9713, 249.9715, 249.9714, 249.9714, 249.9712, 249.9711, 249.9709, 
    249.9707, 249.9706, 249.9706, 249.9708, 249.9711, 249.9713, 249.9713, 
    249.9715, 249.9709, 249.9712, 249.9711, 249.9713, 249.9708, 249.9712, 
    249.9707, 249.9707, 249.9709, 249.9712, 249.9713, 249.9713, 249.9713, 
    249.9711, 249.971, 249.9709, 249.9709, 249.9707, 249.9707, 249.9707, 
    249.9708, 249.9711, 249.9713, 249.9715, 249.9716, 249.9719, 249.9716, 
    249.972, 249.9717, 249.9723, 249.9713, 249.9717, 249.9709, 249.971, 
    249.9711, 249.9715, 249.9713, 249.9715, 249.971, 249.9708, 249.9707, 
    249.9706, 249.9707, 249.9707, 249.9708, 249.9708, 249.9711, 249.9709, 
    249.9714, 249.9715, 249.972, 249.9723, 249.9726, 249.9727, 249.9727, 
    249.9727 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.5157, 258.5161, 258.516, 258.5164, 258.5162, 258.5164, 258.5158, 
    258.5161, 258.5159, 258.5157, 258.517, 258.5164, 258.5176, 258.5172, 
    258.5182, 258.5175, 258.5184, 258.5182, 258.5187, 258.5186, 258.5191, 
    258.5187, 258.5194, 258.519, 258.5191, 258.5187, 258.5165, 258.5169, 
    258.5165, 258.5165, 258.5165, 258.5162, 258.516, 258.5157, 258.5157, 
    258.516, 258.5165, 258.5164, 258.5168, 258.5168, 258.5174, 258.5172, 
    258.5181, 258.5178, 258.5186, 258.5184, 258.5186, 258.5185, 258.5186, 
    258.5182, 258.5184, 258.5181, 258.5172, 258.5175, 258.5166, 258.5161, 
    258.5158, 258.5156, 258.5156, 258.5157, 258.516, 258.5163, 258.5165, 
    258.5167, 258.5168, 258.5173, 258.5175, 258.5181, 258.518, 258.5182, 
    258.5183, 258.5186, 258.5186, 258.5187, 258.5182, 258.5185, 258.5179, 
    258.5181, 258.5168, 258.5164, 258.5162, 258.5161, 258.5156, 258.5159, 
    258.5158, 258.5161, 258.5162, 258.5162, 258.5167, 258.5165, 258.5175, 
    258.5171, 258.5183, 258.518, 258.5184, 258.5182, 258.5185, 258.5182, 
    258.5187, 258.5188, 258.5188, 258.519, 258.5182, 258.5185, 258.5161, 
    258.5162, 258.5162, 258.516, 258.5159, 258.5157, 258.5159, 258.516, 
    258.5163, 258.5164, 258.5165, 258.5168, 258.5172, 258.5177, 258.518, 
    258.5183, 258.5181, 258.5183, 258.5181, 258.5181, 258.5188, 258.5184, 
    258.519, 258.519, 258.5187, 258.519, 258.5162, 258.5161, 258.5158, 
    258.5161, 258.5157, 258.5159, 258.516, 258.5165, 258.5166, 258.5167, 
    258.5169, 258.5172, 258.5176, 258.518, 258.5183, 258.5183, 258.5183, 
    258.5184, 258.5182, 258.5184, 258.5185, 258.5184, 258.519, 258.5188, 
    258.519, 258.5189, 258.5161, 258.5163, 258.5162, 258.5163, 258.5162, 
    258.5167, 258.5168, 258.5174, 258.5172, 258.5175, 258.5172, 258.5172, 
    258.5175, 258.5172, 258.518, 258.5175, 258.5184, 258.5179, 258.5185, 
    258.5183, 258.5185, 258.5187, 258.5189, 258.5192, 258.5191, 258.5194, 
    258.5165, 258.5166, 258.5166, 258.5168, 258.5169, 258.5172, 258.5177, 
    258.5175, 258.5179, 258.5179, 258.5174, 258.5177, 258.5168, 258.5169, 
    258.5168, 258.5165, 258.5176, 258.517, 258.5181, 258.5178, 258.5186, 
    258.5182, 258.5191, 258.5194, 258.5198, 258.5202, 258.5167, 258.5166, 
    258.5168, 258.5171, 258.5174, 258.5178, 258.5178, 258.5179, 258.5181, 
    258.5182, 258.5179, 258.5182, 258.5169, 258.5176, 258.5166, 258.5169, 
    258.5171, 258.517, 258.5175, 258.5176, 258.5181, 258.5179, 258.5193, 
    258.5187, 258.5205, 258.52, 258.5166, 258.5167, 258.5173, 258.517, 
    258.5178, 258.518, 258.5181, 258.5183, 258.5183, 258.5185, 258.5183, 
    258.5185, 258.5178, 258.5181, 258.5172, 258.5174, 258.5173, 258.5172, 
    258.5175, 258.5179, 258.5179, 258.518, 258.5183, 258.5178, 258.5194, 
    258.5184, 258.5169, 258.5172, 258.5173, 258.5172, 258.5179, 258.5177, 
    258.5185, 258.5182, 258.5186, 258.5184, 258.5184, 258.5182, 258.518, 
    258.5177, 258.5174, 258.5172, 258.5172, 258.5175, 258.5179, 258.5183, 
    258.5182, 258.5186, 258.5177, 258.5181, 258.5179, 258.5183, 258.5175, 
    258.5182, 258.5174, 258.5174, 258.5177, 258.5181, 258.5182, 258.5183, 
    258.5182, 258.5179, 258.5179, 258.5176, 258.5176, 258.5174, 258.5173, 
    258.5174, 258.5175, 258.5179, 258.5183, 258.5187, 258.5188, 258.5192, 
    258.5188, 258.5194, 258.5189, 258.5198, 258.5182, 258.5189, 258.5177, 
    258.5178, 258.518, 258.5186, 258.5183, 258.5186, 258.5179, 258.5175, 
    258.5174, 258.5172, 258.5174, 258.5174, 258.5175, 258.5175, 258.5179, 
    258.5177, 258.5184, 258.5186, 258.5194, 258.5198, 258.5203, 258.5205, 
    258.5205, 258.5205 ;

 TREFMXAV_R =
  258.5157, 258.5161, 258.516, 258.5164, 258.5162, 258.5164, 258.5158, 
    258.5161, 258.5159, 258.5157, 258.517, 258.5164, 258.5176, 258.5172, 
    258.5182, 258.5175, 258.5184, 258.5182, 258.5187, 258.5186, 258.5191, 
    258.5187, 258.5194, 258.519, 258.5191, 258.5187, 258.5165, 258.5169, 
    258.5165, 258.5165, 258.5165, 258.5162, 258.516, 258.5157, 258.5157, 
    258.516, 258.5165, 258.5164, 258.5168, 258.5168, 258.5174, 258.5172, 
    258.5181, 258.5178, 258.5186, 258.5184, 258.5186, 258.5185, 258.5186, 
    258.5182, 258.5184, 258.5181, 258.5172, 258.5175, 258.5166, 258.5161, 
    258.5158, 258.5156, 258.5156, 258.5157, 258.516, 258.5163, 258.5165, 
    258.5167, 258.5168, 258.5173, 258.5175, 258.5181, 258.518, 258.5182, 
    258.5183, 258.5186, 258.5186, 258.5187, 258.5182, 258.5185, 258.5179, 
    258.5181, 258.5168, 258.5164, 258.5162, 258.5161, 258.5156, 258.5159, 
    258.5158, 258.5161, 258.5162, 258.5162, 258.5167, 258.5165, 258.5175, 
    258.5171, 258.5183, 258.518, 258.5184, 258.5182, 258.5185, 258.5182, 
    258.5187, 258.5188, 258.5188, 258.519, 258.5182, 258.5185, 258.5161, 
    258.5162, 258.5162, 258.516, 258.5159, 258.5157, 258.5159, 258.516, 
    258.5163, 258.5164, 258.5165, 258.5168, 258.5172, 258.5177, 258.518, 
    258.5183, 258.5181, 258.5183, 258.5181, 258.5181, 258.5188, 258.5184, 
    258.519, 258.519, 258.5187, 258.519, 258.5162, 258.5161, 258.5158, 
    258.5161, 258.5157, 258.5159, 258.516, 258.5165, 258.5166, 258.5167, 
    258.5169, 258.5172, 258.5176, 258.518, 258.5183, 258.5183, 258.5183, 
    258.5184, 258.5182, 258.5184, 258.5185, 258.5184, 258.519, 258.5188, 
    258.519, 258.5189, 258.5161, 258.5163, 258.5162, 258.5163, 258.5162, 
    258.5167, 258.5168, 258.5174, 258.5172, 258.5175, 258.5172, 258.5172, 
    258.5175, 258.5172, 258.518, 258.5175, 258.5184, 258.5179, 258.5185, 
    258.5183, 258.5185, 258.5187, 258.5189, 258.5192, 258.5191, 258.5194, 
    258.5165, 258.5166, 258.5166, 258.5168, 258.5169, 258.5172, 258.5177, 
    258.5175, 258.5179, 258.5179, 258.5174, 258.5177, 258.5168, 258.5169, 
    258.5168, 258.5165, 258.5176, 258.517, 258.5181, 258.5178, 258.5186, 
    258.5182, 258.5191, 258.5194, 258.5198, 258.5202, 258.5167, 258.5166, 
    258.5168, 258.5171, 258.5174, 258.5178, 258.5178, 258.5179, 258.5181, 
    258.5182, 258.5179, 258.5182, 258.5169, 258.5176, 258.5166, 258.5169, 
    258.5171, 258.517, 258.5175, 258.5176, 258.5181, 258.5179, 258.5193, 
    258.5187, 258.5205, 258.52, 258.5166, 258.5167, 258.5173, 258.517, 
    258.5178, 258.518, 258.5181, 258.5183, 258.5183, 258.5185, 258.5183, 
    258.5185, 258.5178, 258.5181, 258.5172, 258.5174, 258.5173, 258.5172, 
    258.5175, 258.5179, 258.5179, 258.518, 258.5183, 258.5178, 258.5194, 
    258.5184, 258.5169, 258.5172, 258.5173, 258.5172, 258.5179, 258.5177, 
    258.5185, 258.5182, 258.5186, 258.5184, 258.5184, 258.5182, 258.518, 
    258.5177, 258.5174, 258.5172, 258.5172, 258.5175, 258.5179, 258.5183, 
    258.5182, 258.5186, 258.5177, 258.5181, 258.5179, 258.5183, 258.5175, 
    258.5182, 258.5174, 258.5174, 258.5177, 258.5181, 258.5182, 258.5183, 
    258.5182, 258.5179, 258.5179, 258.5176, 258.5176, 258.5174, 258.5173, 
    258.5174, 258.5175, 258.5179, 258.5183, 258.5187, 258.5188, 258.5192, 
    258.5188, 258.5194, 258.5189, 258.5198, 258.5182, 258.5189, 258.5177, 
    258.5178, 258.518, 258.5186, 258.5183, 258.5186, 258.5179, 258.5175, 
    258.5174, 258.5172, 258.5174, 258.5174, 258.5175, 258.5175, 258.5179, 
    258.5177, 258.5184, 258.5186, 258.5194, 258.5198, 258.5203, 258.5205, 
    258.5205, 258.5205 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9562, 253.9564, 253.9564, 253.9565, 253.9565, 253.9565, 253.9563, 
    253.9564, 253.9563, 253.9563, 253.9568, 253.9565, 253.9571, 253.9569, 
    253.9573, 253.957, 253.9574, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9576, 253.9579, 253.9577, 253.9577, 253.9576, 253.9566, 253.9568, 
    253.9566, 253.9566, 253.9566, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9564, 253.9566, 253.9565, 253.9567, 253.9567, 253.957, 253.9569, 
    253.9573, 253.9571, 253.9575, 253.9574, 253.9575, 253.9574, 253.9575, 
    253.9574, 253.9574, 253.9573, 253.9569, 253.957, 253.9566, 253.9564, 
    253.9563, 253.9562, 253.9562, 253.9562, 253.9564, 253.9565, 253.9566, 
    253.9567, 253.9567, 253.9569, 253.957, 253.9573, 253.9572, 253.9573, 
    253.9574, 253.9575, 253.9575, 253.9575, 253.9573, 253.9575, 253.9572, 
    253.9573, 253.9567, 253.9565, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9563, 253.9564, 253.9565, 253.9564, 253.9567, 253.9566, 253.957, 
    253.9568, 253.9574, 253.9572, 253.9574, 253.9573, 253.9575, 253.9573, 
    253.9576, 253.9576, 253.9576, 253.9577, 253.9573, 253.9575, 253.9564, 
    253.9565, 253.9565, 253.9563, 253.9563, 253.9562, 253.9563, 253.9564, 
    253.9565, 253.9565, 253.9566, 253.9567, 253.9569, 253.9571, 253.9572, 
    253.9574, 253.9573, 253.9574, 253.9573, 253.9573, 253.9576, 253.9574, 
    253.9577, 253.9577, 253.9575, 253.9577, 253.9565, 253.9564, 253.9563, 
    253.9564, 253.9562, 253.9563, 253.9564, 253.9566, 253.9566, 253.9567, 
    253.9568, 253.9569, 253.9571, 253.9572, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9577, 253.9576, 
    253.9577, 253.9576, 253.9564, 253.9565, 253.9565, 253.9565, 253.9565, 
    253.9566, 253.9567, 253.957, 253.9569, 253.957, 253.9569, 253.9569, 
    253.957, 253.9569, 253.9572, 253.957, 253.9574, 253.9572, 253.9574, 
    253.9574, 253.9575, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9566, 253.9566, 253.9566, 253.9567, 253.9568, 253.9569, 253.9571, 
    253.957, 253.9572, 253.9572, 253.957, 253.9571, 253.9567, 253.9568, 
    253.9567, 253.9566, 253.957, 253.9568, 253.9573, 253.9571, 253.9575, 
    253.9573, 253.9577, 253.9579, 253.958, 253.9582, 253.9567, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9571, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9572, 253.9573, 253.9568, 253.9571, 253.9566, 253.9568, 
    253.9568, 253.9568, 253.957, 253.9571, 253.9573, 253.9572, 253.9578, 
    253.9575, 253.9583, 253.9581, 253.9566, 253.9567, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9573, 253.9574, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9571, 253.9573, 253.9569, 253.957, 253.957, 253.9569, 
    253.957, 253.9572, 253.9572, 253.9572, 253.9574, 253.9571, 253.9578, 
    253.9574, 253.9568, 253.9569, 253.9569, 253.9569, 253.9572, 253.9571, 
    253.9574, 253.9573, 253.9575, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.9571, 253.957, 253.9569, 253.9569, 253.957, 253.9572, 253.9574, 
    253.9573, 253.9575, 253.9571, 253.9573, 253.9572, 253.9574, 253.957, 
    253.9573, 253.957, 253.957, 253.9571, 253.9573, 253.9573, 253.9574, 
    253.9573, 253.9572, 253.9572, 253.9571, 253.9571, 253.957, 253.9569, 
    253.957, 253.957, 253.9572, 253.9574, 253.9575, 253.9576, 253.9577, 
    253.9576, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.9571, 
    253.9572, 253.9572, 253.9575, 253.9574, 253.9575, 253.9572, 253.957, 
    253.957, 253.9569, 253.957, 253.957, 253.957, 253.957, 253.9572, 
    253.9571, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9562, 253.9564, 253.9564, 253.9565, 253.9565, 253.9565, 253.9563, 
    253.9564, 253.9563, 253.9563, 253.9568, 253.9565, 253.9571, 253.9569, 
    253.9573, 253.957, 253.9574, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9576, 253.9579, 253.9577, 253.9577, 253.9576, 253.9566, 253.9568, 
    253.9566, 253.9566, 253.9566, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9564, 253.9566, 253.9565, 253.9567, 253.9567, 253.957, 253.9569, 
    253.9573, 253.9571, 253.9575, 253.9574, 253.9575, 253.9574, 253.9575, 
    253.9574, 253.9574, 253.9573, 253.9569, 253.957, 253.9566, 253.9564, 
    253.9563, 253.9562, 253.9562, 253.9562, 253.9564, 253.9565, 253.9566, 
    253.9567, 253.9567, 253.9569, 253.957, 253.9573, 253.9572, 253.9573, 
    253.9574, 253.9575, 253.9575, 253.9575, 253.9573, 253.9575, 253.9572, 
    253.9573, 253.9567, 253.9565, 253.9565, 253.9564, 253.9562, 253.9563, 
    253.9563, 253.9564, 253.9565, 253.9564, 253.9567, 253.9566, 253.957, 
    253.9568, 253.9574, 253.9572, 253.9574, 253.9573, 253.9575, 253.9573, 
    253.9576, 253.9576, 253.9576, 253.9577, 253.9573, 253.9575, 253.9564, 
    253.9565, 253.9565, 253.9563, 253.9563, 253.9562, 253.9563, 253.9564, 
    253.9565, 253.9565, 253.9566, 253.9567, 253.9569, 253.9571, 253.9572, 
    253.9574, 253.9573, 253.9574, 253.9573, 253.9573, 253.9576, 253.9574, 
    253.9577, 253.9577, 253.9575, 253.9577, 253.9565, 253.9564, 253.9563, 
    253.9564, 253.9562, 253.9563, 253.9564, 253.9566, 253.9566, 253.9567, 
    253.9568, 253.9569, 253.9571, 253.9572, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9577, 253.9576, 
    253.9577, 253.9576, 253.9564, 253.9565, 253.9565, 253.9565, 253.9565, 
    253.9566, 253.9567, 253.957, 253.9569, 253.957, 253.9569, 253.9569, 
    253.957, 253.9569, 253.9572, 253.957, 253.9574, 253.9572, 253.9574, 
    253.9574, 253.9575, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9566, 253.9566, 253.9566, 253.9567, 253.9568, 253.9569, 253.9571, 
    253.957, 253.9572, 253.9572, 253.957, 253.9571, 253.9567, 253.9568, 
    253.9567, 253.9566, 253.957, 253.9568, 253.9573, 253.9571, 253.9575, 
    253.9573, 253.9577, 253.9579, 253.958, 253.9582, 253.9567, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9571, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9572, 253.9573, 253.9568, 253.9571, 253.9566, 253.9568, 
    253.9568, 253.9568, 253.957, 253.9571, 253.9573, 253.9572, 253.9578, 
    253.9575, 253.9583, 253.9581, 253.9566, 253.9567, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9573, 253.9574, 253.9574, 253.9574, 253.9574, 
    253.9574, 253.9571, 253.9573, 253.9569, 253.957, 253.957, 253.9569, 
    253.957, 253.9572, 253.9572, 253.9572, 253.9574, 253.9571, 253.9578, 
    253.9574, 253.9568, 253.9569, 253.9569, 253.9569, 253.9572, 253.9571, 
    253.9574, 253.9573, 253.9575, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.9571, 253.957, 253.9569, 253.9569, 253.957, 253.9572, 253.9574, 
    253.9573, 253.9575, 253.9571, 253.9573, 253.9572, 253.9574, 253.957, 
    253.9573, 253.957, 253.957, 253.9571, 253.9573, 253.9573, 253.9574, 
    253.9573, 253.9572, 253.9572, 253.9571, 253.9571, 253.957, 253.9569, 
    253.957, 253.957, 253.9572, 253.9574, 253.9575, 253.9576, 253.9577, 
    253.9576, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.9571, 
    253.9572, 253.9572, 253.9575, 253.9574, 253.9575, 253.9572, 253.957, 
    253.957, 253.9569, 253.957, 253.957, 253.957, 253.957, 253.9572, 
    253.9571, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.3913, 254.3927, 254.3925, 254.3936, 254.393, 254.3937, 254.3916, 
    254.3928, 254.392, 254.3914, 254.3958, 254.3937, 254.3982, 254.3968, 
    254.4003, 254.3979, 254.4008, 254.4003, 254.4019, 254.4014, 254.4035, 
    254.4021, 254.4046, 254.4032, 254.4034, 254.4021, 254.3941, 254.3955, 
    254.394, 254.3942, 254.3941, 254.393, 254.3924, 254.3912, 254.3914, 
    254.3923, 254.3943, 254.3937, 254.3954, 254.3954, 254.3973, 254.3964, 
    254.3997, 254.3988, 254.4015, 254.4008, 254.4014, 254.4012, 254.4014, 
    254.4004, 254.4009, 254.4, 254.3966, 254.3976, 254.3946, 254.3928, 
    254.3916, 254.3908, 254.3909, 254.3912, 254.3923, 254.3934, 254.3943, 
    254.3948, 254.3954, 254.397, 254.3979, 254.3999, 254.3995, 254.4001, 
    254.4007, 254.4017, 254.4015, 254.402, 254.4001, 254.4013, 254.3993, 
    254.3999, 254.3954, 254.3938, 254.3931, 254.3925, 254.391, 254.3921, 
    254.3916, 254.3926, 254.3932, 254.3929, 254.3948, 254.3941, 254.3979, 
    254.3963, 254.4007, 254.3996, 254.4009, 254.4002, 254.4014, 254.4004, 
    254.4021, 254.4025, 254.4022, 254.4033, 254.4003, 254.4014, 254.3929, 
    254.393, 254.3932, 254.3922, 254.3921, 254.3912, 254.392, 254.3924, 
    254.3933, 254.3938, 254.3943, 254.3954, 254.3967, 254.3984, 254.3997, 
    254.4005, 254.4, 254.4005, 254.3999, 254.3997, 254.4023, 254.4008, 
    254.4031, 254.403, 254.402, 254.403, 254.393, 254.3927, 254.3917, 
    254.3925, 254.3911, 254.3919, 254.3923, 254.3941, 254.3945, 254.3948, 
    254.3956, 254.3965, 254.3981, 254.3995, 254.4008, 254.4007, 254.4007, 
    254.401, 254.4003, 254.4011, 254.4012, 254.4009, 254.403, 254.4024, 
    254.403, 254.4026, 254.3928, 254.3933, 254.3931, 254.3935, 254.3932, 
    254.3947, 254.3951, 254.3973, 254.3964, 254.3978, 254.3966, 254.3968, 
    254.3978, 254.3967, 254.3994, 254.3975, 254.401, 254.3991, 254.4011, 
    254.4007, 254.4013, 254.4019, 254.4025, 254.4038, 254.4035, 254.4045, 
    254.394, 254.3946, 254.3946, 254.3952, 254.3957, 254.3968, 254.3985, 
    254.3978, 254.399, 254.3992, 254.3975, 254.3985, 254.3951, 254.3956, 
    254.3953, 254.3941, 254.3979, 254.3959, 254.3997, 254.3986, 254.4018, 
    254.4002, 254.4033, 254.4046, 254.4059, 254.4074, 254.395, 254.3946, 
    254.3953, 254.3963, 254.3974, 254.3987, 254.3988, 254.399, 254.3997, 
    254.4002, 254.3991, 254.4003, 254.3957, 254.3981, 254.3944, 254.3955, 
    254.3963, 254.396, 254.3978, 254.3982, 254.3999, 254.399, 254.4043, 
    254.4019, 254.4086, 254.4067, 254.3944, 254.395, 254.397, 254.396, 
    254.3988, 254.3994, 254.4, 254.4007, 254.4007, 254.4012, 254.4005, 
    254.4011, 254.3987, 254.3998, 254.3968, 254.3975, 254.3972, 254.3968, 
    254.3979, 254.3991, 254.3992, 254.3995, 254.4005, 254.3988, 254.4045, 
    254.4009, 254.3956, 254.3967, 254.3969, 254.3965, 254.3994, 254.3983, 
    254.4012, 254.4004, 254.4016, 254.401, 254.4009, 254.4001, 254.3996, 
    254.3983, 254.3973, 254.3965, 254.3967, 254.3976, 254.3992, 254.4007, 
    254.4004, 254.4016, 254.3986, 254.3998, 254.3993, 254.4006, 254.3978, 
    254.4001, 254.3972, 254.3975, 254.3983, 254.3999, 254.4003, 254.4006, 
    254.4004, 254.3992, 254.3991, 254.3983, 254.398, 254.3974, 254.3969, 
    254.3974, 254.3978, 254.3992, 254.4005, 254.4019, 254.4022, 254.4037, 
    254.4025, 254.4046, 254.4027, 254.4059, 254.4003, 254.4027, 254.3983, 
    254.3988, 254.3996, 254.4016, 254.4006, 254.4018, 254.399, 254.3976, 
    254.3972, 254.3966, 254.3973, 254.3972, 254.3979, 254.3977, 254.3993, 
    254.3984, 254.4009, 254.4018, 254.4044, 254.406, 254.4076, 254.4084, 
    254.4086, 254.4087,
  255.5014, 255.5029, 255.5026, 255.5038, 255.5031, 255.5039, 255.5017, 
    255.5029, 255.5021, 255.5015, 255.506, 255.5038, 255.5084, 255.507, 
    255.5107, 255.5082, 255.5112, 255.5106, 255.5123, 255.5118, 255.514, 
    255.5126, 255.5152, 255.5137, 255.5139, 255.5125, 255.5043, 255.5057, 
    255.5042, 255.5044, 255.5043, 255.5031, 255.5025, 255.5013, 255.5015, 
    255.5024, 255.5045, 255.5038, 255.5056, 255.5056, 255.5076, 255.5067, 
    255.51, 255.5091, 255.5119, 255.5112, 255.5118, 255.5116, 255.5118, 
    255.5108, 255.5112, 255.5103, 255.5068, 255.5078, 255.5048, 255.5029, 
    255.5017, 255.5009, 255.501, 255.5012, 255.5024, 255.5036, 255.5044, 
    255.505, 255.5056, 255.5072, 255.5081, 255.5102, 255.5099, 255.5105, 
    255.5111, 255.5121, 255.5119, 255.5124, 255.5105, 255.5117, 255.5097, 
    255.5102, 255.5056, 255.504, 255.5032, 255.5026, 255.5011, 255.5022, 
    255.5017, 255.5027, 255.5034, 255.5031, 255.505, 255.5042, 255.5082, 
    255.5065, 255.511, 255.5099, 255.5113, 255.5106, 255.5118, 255.5107, 
    255.5125, 255.5129, 255.5127, 255.5137, 255.5107, 255.5118, 255.5031, 
    255.5031, 255.5033, 255.5023, 255.5022, 255.5013, 255.5021, 255.5025, 
    255.5034, 255.504, 255.5045, 255.5056, 255.5069, 255.5087, 255.51, 
    255.5109, 255.5103, 255.5108, 255.5103, 255.51, 255.5128, 255.5112, 
    255.5136, 255.5134, 255.5124, 255.5135, 255.5031, 255.5029, 255.5018, 
    255.5026, 255.5012, 255.502, 255.5024, 255.5042, 255.5047, 255.505, 
    255.5058, 255.5067, 255.5083, 255.5098, 255.5111, 255.511, 255.5111, 
    255.5114, 255.5106, 255.5115, 255.5116, 255.5112, 255.5134, 255.5128, 
    255.5134, 255.513, 255.5029, 255.5034, 255.5032, 255.5037, 255.5033, 
    255.5049, 255.5053, 255.5076, 255.5067, 255.5081, 255.5068, 255.507, 
    255.5081, 255.5069, 255.5097, 255.5078, 255.5114, 255.5094, 255.5115, 
    255.5111, 255.5117, 255.5123, 255.513, 255.5143, 255.514, 255.515, 
    255.5042, 255.5048, 255.5048, 255.5054, 255.5059, 255.507, 255.5088, 
    255.5081, 255.5093, 255.5096, 255.5077, 255.5088, 255.5052, 255.5058, 
    255.5055, 255.5042, 255.5082, 255.5061, 255.51, 255.5089, 255.5122, 
    255.5105, 255.5138, 255.5152, 255.5165, 255.518, 255.5052, 255.5047, 
    255.5055, 255.5066, 255.5076, 255.509, 255.5091, 255.5094, 255.51, 
    255.5106, 255.5094, 255.5107, 255.5059, 255.5084, 255.5046, 255.5057, 
    255.5065, 255.5062, 255.508, 255.5085, 255.5102, 255.5093, 255.5148, 
    255.5124, 255.5192, 255.5173, 255.5046, 255.5052, 255.5072, 255.5062, 
    255.509, 255.5098, 255.5103, 255.511, 255.5111, 255.5115, 255.5108, 
    255.5115, 255.509, 255.5101, 255.507, 255.5077, 255.5074, 255.507, 
    255.5082, 255.5094, 255.5095, 255.5099, 255.5109, 255.5091, 255.5151, 
    255.5113, 255.5058, 255.5069, 255.5071, 255.5067, 255.5097, 255.5086, 
    255.5115, 255.5107, 255.5121, 255.5114, 255.5113, 255.5105, 255.5099, 
    255.5086, 255.5076, 255.5067, 255.5069, 255.5078, 255.5095, 255.5111, 
    255.5108, 255.5119, 255.5089, 255.5101, 255.5096, 255.511, 255.5081, 
    255.5104, 255.5075, 255.5077, 255.5086, 255.5102, 255.5106, 255.511, 
    255.5108, 255.5096, 255.5094, 255.5085, 255.5083, 255.5077, 255.5072, 
    255.5076, 255.5081, 255.5096, 255.5109, 255.5123, 255.5126, 255.5143, 
    255.5129, 255.5151, 255.5132, 255.5165, 255.5106, 255.5132, 255.5086, 
    255.5091, 255.51, 255.512, 255.5109, 255.5122, 255.5094, 255.5079, 
    255.5075, 255.5068, 255.5075, 255.5075, 255.5082, 255.5079, 255.5096, 
    255.5087, 255.5113, 255.5122, 255.5149, 255.5166, 255.5183, 255.519, 
    255.5193, 255.5194,
  257.1078, 257.1091, 257.1089, 257.1099, 257.1093, 257.11, 257.1081, 
    257.1091, 257.1085, 257.1079, 257.112, 257.11, 257.1142, 257.1129, 
    257.1162, 257.114, 257.1167, 257.1162, 257.1177, 257.1173, 257.1193, 
    257.118, 257.1203, 257.119, 257.1192, 257.1179, 257.1104, 257.1117, 
    257.1103, 257.1105, 257.1104, 257.1093, 257.1088, 257.1077, 257.1079, 
    257.1087, 257.1106, 257.11, 257.1116, 257.1115, 257.1134, 257.1125, 
    257.1156, 257.1147, 257.1173, 257.1167, 257.1173, 257.1171, 257.1173, 
    257.1163, 257.1167, 257.1159, 257.1127, 257.1136, 257.1108, 257.1092, 
    257.1081, 257.1073, 257.1074, 257.1076, 257.1087, 257.1097, 257.1105, 
    257.111, 257.1115, 257.113, 257.1139, 257.1158, 257.1155, 257.116, 
    257.1166, 257.1175, 257.1174, 257.1178, 257.116, 257.1172, 257.1153, 
    257.1158, 257.1116, 257.1101, 257.1094, 257.1089, 257.1075, 257.1085, 
    257.1081, 257.109, 257.1096, 257.1093, 257.1111, 257.1104, 257.114, 
    257.1124, 257.1165, 257.1155, 257.1168, 257.1161, 257.1172, 257.1162, 
    257.1179, 257.1183, 257.118, 257.119, 257.1162, 257.1173, 257.1093, 
    257.1093, 257.1095, 257.1086, 257.1085, 257.1077, 257.1084, 257.1088, 
    257.1096, 257.1101, 257.1106, 257.1116, 257.1128, 257.1144, 257.1156, 
    257.1164, 257.1159, 257.1163, 257.1159, 257.1156, 257.1182, 257.1167, 
    257.1189, 257.1188, 257.1178, 257.1188, 257.1093, 257.1091, 257.1082, 
    257.1089, 257.1076, 257.1083, 257.1087, 257.1104, 257.1107, 257.1111, 
    257.1117, 257.1126, 257.1141, 257.1154, 257.1166, 257.1165, 257.1166, 
    257.1169, 257.1162, 257.1169, 257.1171, 257.1167, 257.1187, 257.1182, 
    257.1188, 257.1184, 257.1092, 257.1096, 257.1094, 257.1098, 257.1095, 
    257.1109, 257.1114, 257.1134, 257.1125, 257.1139, 257.1127, 257.1129, 
    257.1139, 257.1128, 257.1153, 257.1136, 257.1169, 257.1151, 257.117, 
    257.1166, 257.1172, 257.1177, 257.1183, 257.1195, 257.1192, 257.1202, 
    257.1103, 257.1109, 257.1108, 257.1115, 257.1119, 257.1129, 257.1145, 
    257.1139, 257.115, 257.1152, 257.1135, 257.1145, 257.1113, 257.1118, 
    257.1115, 257.1103, 257.114, 257.1121, 257.1156, 257.1146, 257.1176, 
    257.1161, 257.1191, 257.1203, 257.1216, 257.123, 257.1112, 257.1108, 
    257.1115, 257.1125, 257.1134, 257.1147, 257.1148, 257.115, 257.1156, 
    257.1161, 257.1151, 257.1162, 257.1118, 257.1142, 257.1106, 257.1117, 
    257.1124, 257.1121, 257.1138, 257.1142, 257.1158, 257.115, 257.12, 
    257.1178, 257.1241, 257.1223, 257.1107, 257.1112, 257.113, 257.1122, 
    257.1147, 257.1154, 257.1159, 257.1165, 257.1166, 257.117, 257.1164, 
    257.117, 257.1147, 257.1157, 257.1129, 257.1135, 257.1132, 257.1129, 
    257.114, 257.1151, 257.1151, 257.1155, 257.1165, 257.1147, 257.1203, 
    257.1168, 257.1118, 257.1128, 257.1129, 257.1125, 257.1153, 257.1143, 
    257.117, 257.1163, 257.1175, 257.1169, 257.1168, 257.116, 257.1155, 
    257.1143, 257.1134, 257.1126, 257.1128, 257.1136, 257.1151, 257.1166, 
    257.1163, 257.1174, 257.1145, 257.1157, 257.1153, 257.1165, 257.1139, 
    257.116, 257.1133, 257.1135, 257.1143, 257.1158, 257.1161, 257.1165, 
    257.1163, 257.1152, 257.115, 257.1143, 257.114, 257.1135, 257.113, 
    257.1134, 257.1139, 257.1152, 257.1164, 257.1177, 257.118, 257.1195, 
    257.1183, 257.1203, 257.1185, 257.1216, 257.1162, 257.1185, 257.1143, 
    257.1148, 257.1156, 257.1175, 257.1165, 257.1176, 257.115, 257.1136, 
    257.1133, 257.1127, 257.1133, 257.1133, 257.1139, 257.1137, 257.1152, 
    257.1144, 257.1168, 257.1176, 257.1201, 257.1216, 257.1232, 257.1239, 
    257.1241, 257.1242,
  259.2219, 259.2228, 259.2226, 259.2234, 259.223, 259.2235, 259.222, 
    259.2228, 259.2224, 259.222, 259.2249, 259.2234, 259.2265, 259.2256, 
    259.228, 259.2263, 259.2284, 259.228, 259.2292, 259.2288, 259.2303, 
    259.2293, 259.2311, 259.23, 259.2302, 259.2292, 259.2238, 259.2247, 
    259.2237, 259.2238, 259.2238, 259.223, 259.2226, 259.2218, 259.2219, 
    259.2225, 259.2239, 259.2234, 259.2246, 259.2246, 259.2259, 259.2253, 
    259.2276, 259.2269, 259.2288, 259.2283, 259.2288, 259.2287, 259.2288, 
    259.2281, 259.2284, 259.2278, 259.2254, 259.2261, 259.2241, 259.2228, 
    259.2221, 259.2215, 259.2216, 259.2218, 259.2225, 259.2233, 259.2238, 
    259.2242, 259.2246, 259.2257, 259.2263, 259.2277, 259.2274, 259.2279, 
    259.2283, 259.229, 259.2289, 259.2292, 259.2279, 259.2287, 259.2273, 
    259.2277, 259.2246, 259.2236, 259.2231, 259.2227, 259.2217, 259.2224, 
    259.2221, 259.2227, 259.2231, 259.223, 259.2242, 259.2237, 259.2263, 
    259.2252, 259.2282, 259.2275, 259.2284, 259.228, 259.2288, 259.228, 
    259.2293, 259.2296, 259.2294, 259.2301, 259.228, 259.2288, 259.2229, 
    259.223, 259.2231, 259.2224, 259.2224, 259.2218, 259.2224, 259.2226, 
    259.2232, 259.2235, 259.2239, 259.2246, 259.2255, 259.2267, 259.2276, 
    259.2281, 259.2278, 259.2281, 259.2278, 259.2276, 259.2295, 259.2284, 
    259.23, 259.2299, 259.2292, 259.2299, 259.223, 259.2228, 259.2221, 
    259.2227, 259.2217, 259.2222, 259.2225, 259.2237, 259.224, 259.2242, 
    259.2247, 259.2253, 259.2264, 259.2274, 259.2283, 259.2282, 259.2283, 
    259.2285, 259.228, 259.2285, 259.2286, 259.2284, 259.2299, 259.2295, 
    259.2299, 259.2296, 259.2229, 259.2232, 259.223, 259.2233, 259.2231, 
    259.2241, 259.2245, 259.2259, 259.2253, 259.2263, 259.2254, 259.2256, 
    259.2263, 259.2255, 259.2274, 259.226, 259.2285, 259.2271, 259.2286, 
    259.2283, 259.2287, 259.2291, 259.2296, 259.2305, 259.2303, 259.231, 
    259.2237, 259.2241, 259.2241, 259.2245, 259.2248, 259.2256, 259.2267, 
    259.2263, 259.2271, 259.2273, 259.226, 259.2268, 259.2244, 259.2248, 
    259.2245, 259.2237, 259.2264, 259.225, 259.2276, 259.2268, 259.229, 
    259.2279, 259.2301, 259.2311, 259.232, 259.2331, 259.2243, 259.2241, 
    259.2246, 259.2253, 259.226, 259.2269, 259.227, 259.2271, 259.2276, 
    259.2279, 259.2272, 259.228, 259.2248, 259.2265, 259.2239, 259.2247, 
    259.2252, 259.225, 259.2262, 259.2265, 259.2277, 259.2271, 259.2308, 
    259.2292, 259.2339, 259.2326, 259.2239, 259.2243, 259.2257, 259.225, 
    259.2269, 259.2274, 259.2278, 259.2282, 259.2283, 259.2286, 259.2281, 
    259.2286, 259.2269, 259.2276, 259.2256, 259.226, 259.2258, 259.2256, 
    259.2263, 259.2272, 259.2272, 259.2275, 259.2282, 259.2269, 259.231, 
    259.2285, 259.2248, 259.2255, 259.2256, 259.2253, 259.2273, 259.2266, 
    259.2286, 259.2281, 259.2289, 259.2285, 259.2284, 259.2279, 259.2275, 
    259.2266, 259.2259, 259.2254, 259.2255, 259.2261, 259.2272, 259.2283, 
    259.2281, 259.2289, 259.2268, 259.2277, 259.2273, 259.2282, 259.2263, 
    259.2278, 259.2259, 259.226, 259.2266, 259.2277, 259.228, 259.2282, 
    259.2281, 259.2273, 259.2271, 259.2266, 259.2264, 259.226, 259.2256, 
    259.226, 259.2263, 259.2273, 259.2281, 259.2291, 259.2293, 259.2304, 
    259.2295, 259.231, 259.2297, 259.232, 259.228, 259.2297, 259.2266, 
    259.227, 259.2275, 259.2289, 259.2282, 259.2291, 259.2271, 259.2261, 
    259.2259, 259.2254, 259.2259, 259.2259, 259.2263, 259.2262, 259.2273, 
    259.2267, 259.2284, 259.2291, 259.2309, 259.2321, 259.2332, 259.2338, 
    259.2339, 259.234,
  261.4064, 261.4069, 261.4068, 261.4071, 261.407, 261.4072, 261.4065, 
    261.4069, 261.4066, 261.4065, 261.4078, 261.4072, 261.4086, 261.4081, 
    261.4094, 261.4085, 261.4095, 261.4093, 261.4099, 261.4097, 261.4105, 
    261.41, 261.4109, 261.4104, 261.4104, 261.41, 261.4073, 261.4077, 
    261.4073, 261.4073, 261.4073, 261.407, 261.4067, 261.4064, 261.4065, 
    261.4067, 261.4073, 261.4071, 261.4077, 261.4077, 261.4083, 261.4081, 
    261.4091, 261.4088, 261.4098, 261.4095, 261.4097, 261.4097, 261.4097, 
    261.4094, 261.4095, 261.4092, 261.4081, 261.4084, 261.4074, 261.4069, 
    261.4065, 261.4063, 261.4063, 261.4064, 261.4067, 261.4071, 261.4073, 
    261.4075, 261.4077, 261.4082, 261.4085, 261.4092, 261.4091, 261.4093, 
    261.4095, 261.4098, 261.4098, 261.4099, 261.4093, 261.4097, 261.409, 
    261.4092, 261.4077, 261.4072, 261.407, 261.4068, 261.4063, 261.4066, 
    261.4065, 261.4068, 261.407, 261.4069, 261.4075, 261.4073, 261.4085, 
    261.408, 261.4095, 261.4091, 261.4095, 261.4093, 261.4097, 261.4094, 
    261.41, 261.4101, 261.41, 261.4104, 261.4093, 261.4097, 261.4069, 
    261.4069, 261.407, 261.4067, 261.4067, 261.4064, 261.4066, 261.4067, 
    261.407, 261.4072, 261.4073, 261.4077, 261.4081, 261.4087, 261.4091, 
    261.4094, 261.4092, 261.4094, 261.4092, 261.4091, 261.4101, 261.4095, 
    261.4103, 261.4103, 261.4099, 261.4103, 261.407, 261.4069, 261.4066, 
    261.4068, 261.4063, 261.4066, 261.4067, 261.4073, 261.4074, 261.4075, 
    261.4077, 261.4081, 261.4086, 261.4091, 261.4095, 261.4095, 261.4095, 
    261.4096, 261.4093, 261.4096, 261.4097, 261.4095, 261.4103, 261.4101, 
    261.4103, 261.4102, 261.4069, 261.407, 261.407, 261.4071, 261.407, 
    261.4075, 261.4076, 261.4083, 261.4081, 261.4085, 261.4081, 261.4082, 
    261.4085, 261.4081, 261.409, 261.4084, 261.4096, 261.4089, 261.4096, 
    261.4095, 261.4097, 261.4099, 261.4101, 261.4106, 261.4105, 261.4108, 
    261.4073, 261.4075, 261.4074, 261.4077, 261.4078, 261.4082, 261.4087, 
    261.4085, 261.4089, 261.409, 261.4084, 261.4088, 261.4076, 261.4078, 
    261.4077, 261.4073, 261.4085, 261.4079, 261.4091, 261.4088, 261.4099, 
    261.4093, 261.4104, 261.4109, 261.4113, 261.4119, 261.4076, 261.4074, 
    261.4077, 261.408, 261.4084, 261.4088, 261.4088, 261.4089, 261.4091, 
    261.4093, 261.4089, 261.4094, 261.4078, 261.4086, 261.4074, 261.4077, 
    261.408, 261.4079, 261.4085, 261.4086, 261.4092, 261.4089, 261.4108, 
    261.4099, 261.4123, 261.4116, 261.4074, 261.4076, 261.4082, 261.4079, 
    261.4088, 261.4091, 261.4092, 261.4095, 261.4095, 261.4096, 261.4094, 
    261.4096, 261.4088, 261.4091, 261.4081, 261.4084, 261.4083, 261.4082, 
    261.4085, 261.4089, 261.409, 261.4091, 261.4094, 261.4088, 261.4109, 
    261.4096, 261.4078, 261.4081, 261.4082, 261.4081, 261.409, 261.4087, 
    261.4096, 261.4094, 261.4098, 261.4096, 261.4095, 261.4093, 261.4091, 
    261.4087, 261.4083, 261.4081, 261.4081, 261.4084, 261.409, 261.4095, 
    261.4094, 261.4098, 261.4088, 261.4092, 261.409, 261.4095, 261.4085, 
    261.4093, 261.4083, 261.4084, 261.4087, 261.4092, 261.4093, 261.4095, 
    261.4094, 261.409, 261.4089, 261.4087, 261.4086, 261.4084, 261.4082, 
    261.4084, 261.4085, 261.409, 261.4094, 261.4099, 261.41, 261.4106, 
    261.4101, 261.4109, 261.4102, 261.4113, 261.4093, 261.4102, 261.4087, 
    261.4088, 261.4091, 261.4098, 261.4095, 261.4099, 261.4089, 261.4084, 
    261.4083, 261.4081, 261.4083, 261.4083, 261.4085, 261.4084, 261.409, 
    261.4087, 261.4095, 261.4099, 261.4108, 261.4114, 261.412, 261.4122, 
    261.4123, 261.4124,
  262.7626, 262.7627, 262.7627, 262.7628, 262.7627, 262.7628, 262.7626, 
    262.7627, 262.7627, 262.7626, 262.7629, 262.7628, 262.7631, 262.763, 
    262.7633, 262.7631, 262.7633, 262.7633, 262.7635, 262.7634, 262.7636, 
    262.7635, 262.7637, 262.7635, 262.7636, 262.7635, 262.7628, 262.7629, 
    262.7628, 262.7628, 262.7628, 262.7627, 262.7627, 262.7626, 262.7626, 
    262.7627, 262.7628, 262.7628, 262.7629, 262.7629, 262.7631, 262.763, 
    262.7632, 262.7632, 262.7634, 262.7633, 262.7634, 262.7634, 262.7634, 
    262.7633, 262.7634, 262.7633, 262.763, 262.7631, 262.7628, 262.7627, 
    262.7626, 262.7626, 262.7626, 262.7626, 262.7627, 262.7628, 262.7628, 
    262.7629, 262.7629, 262.763, 262.7631, 262.7633, 262.7632, 262.7633, 
    262.7633, 262.7634, 262.7634, 262.7635, 262.7633, 262.7634, 262.7632, 
    262.7633, 262.7629, 262.7628, 262.7628, 262.7627, 262.7626, 262.7627, 
    262.7626, 262.7627, 262.7628, 262.7627, 262.7629, 262.7628, 262.7631, 
    262.763, 262.7633, 262.7632, 262.7634, 262.7633, 262.7634, 262.7633, 
    262.7635, 262.7635, 262.7635, 262.7635, 262.7633, 262.7634, 262.7627, 
    262.7627, 262.7628, 262.7627, 262.7627, 262.7626, 262.7627, 262.7627, 
    262.7628, 262.7628, 262.7628, 262.7629, 262.763, 262.7632, 262.7632, 
    262.7633, 262.7633, 262.7633, 262.7633, 262.7632, 262.7635, 262.7634, 
    262.7635, 262.7635, 262.7635, 262.7635, 262.7627, 262.7627, 262.7626, 
    262.7627, 262.7626, 262.7627, 262.7627, 262.7628, 262.7628, 262.7629, 
    262.7629, 262.763, 262.7631, 262.7632, 262.7633, 262.7633, 262.7633, 
    262.7634, 262.7633, 262.7634, 262.7634, 262.7634, 262.7635, 262.7635, 
    262.7635, 262.7635, 262.7627, 262.7628, 262.7627, 262.7628, 262.7628, 
    262.7628, 262.7629, 262.7631, 262.763, 262.7631, 262.763, 262.763, 
    262.7631, 262.763, 262.7632, 262.7631, 262.7634, 262.7632, 262.7634, 
    262.7633, 262.7634, 262.7634, 262.7635, 262.7636, 262.7636, 262.7637, 
    262.7628, 262.7628, 262.7628, 262.7629, 262.7629, 262.763, 262.7632, 
    262.7631, 262.7632, 262.7632, 262.7631, 262.7632, 262.7629, 262.7629, 
    262.7629, 262.7628, 262.7631, 262.763, 262.7632, 262.7632, 262.7634, 
    262.7633, 262.7636, 262.7637, 262.7638, 262.7639, 262.7629, 262.7628, 
    262.7629, 262.763, 262.7631, 262.7632, 262.7632, 262.7632, 262.7632, 
    262.7633, 262.7632, 262.7633, 262.7629, 262.7631, 262.7628, 262.7629, 
    262.763, 262.763, 262.7631, 262.7631, 262.7633, 262.7632, 262.7637, 
    262.7635, 262.7641, 262.7639, 262.7628, 262.7629, 262.763, 262.763, 
    262.7632, 262.7632, 262.7633, 262.7633, 262.7633, 262.7634, 262.7633, 
    262.7634, 262.7632, 262.7633, 262.763, 262.7631, 262.7631, 262.763, 
    262.7631, 262.7632, 262.7632, 262.7632, 262.7633, 262.7632, 262.7637, 
    262.7634, 262.7629, 262.763, 262.763, 262.763, 262.7632, 262.7632, 
    262.7634, 262.7633, 262.7634, 262.7634, 262.7634, 262.7633, 262.7632, 
    262.7632, 262.7631, 262.763, 262.763, 262.7631, 262.7632, 262.7633, 
    262.7633, 262.7634, 262.7632, 262.7633, 262.7632, 262.7633, 262.7631, 
    262.7633, 262.7631, 262.7631, 262.7632, 262.7633, 262.7633, 262.7633, 
    262.7633, 262.7632, 262.7632, 262.7631, 262.7631, 262.7631, 262.763, 
    262.7631, 262.7631, 262.7632, 262.7633, 262.7634, 262.7635, 262.7636, 
    262.7635, 262.7637, 262.7635, 262.7638, 262.7633, 262.7635, 262.7632, 
    262.7632, 262.7632, 262.7634, 262.7633, 262.7634, 262.7632, 262.7631, 
    262.7631, 262.763, 262.7631, 262.7631, 262.7631, 262.7631, 262.7632, 
    262.7632, 262.7634, 262.7634, 262.7637, 262.7638, 262.764, 262.764, 
    262.7641, 262.7641,
  263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 
    263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1179, 263.1179, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1177, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1179, 263.1177, 263.1177, 263.1178, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1178, 263.1178, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1179, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 
    263.1179, 263.1179,
  263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  262.9297, 262.9442, 262.9414, 262.9531, 262.9466, 262.9542, 262.9327, 
    262.9448, 262.9371, 262.9311, 262.9756, 262.9536, 262.9984, 262.9844, 
    263.0195, 262.9962, 263.0242, 263.0188, 263.0349, 263.0303, 263.0509, 
    263.0371, 263.0615, 263.0476, 263.0498, 263.0366, 262.958, 262.9728, 
    262.9572, 262.9593, 262.9583, 262.9467, 262.9409, 262.9287, 262.9309, 
    262.9399, 262.9602, 262.9533, 262.9707, 262.9703, 262.9896, 262.9809, 
    263.0132, 263.0041, 263.0305, 263.0239, 263.0302, 263.0283, 263.0302, 
    263.0205, 263.0247, 263.0161, 262.9825, 262.9924, 262.9629, 262.9451, 
    262.9332, 262.9248, 262.926, 262.9283, 262.9399, 262.9509, 262.9592, 
    262.9648, 262.9702, 262.9868, 262.9955, 263.015, 263.0115, 263.0175, 
    263.0232, 263.0328, 263.0312, 263.0354, 263.0174, 263.0294, 263.0096, 
    263.015, 262.9716, 262.9552, 262.9481, 262.942, 262.9269, 262.9373, 
    262.9332, 262.943, 262.9492, 262.9461, 262.9649, 262.9576, 262.996, 
    262.9795, 263.0226, 263.0123, 263.025, 263.0185, 263.0296, 263.0196, 
    263.037, 263.0407, 263.0381, 263.0481, 263.0191, 263.0302, 262.946, 
    262.9465, 262.9488, 262.9386, 262.938, 262.9286, 262.937, 262.9405, 
    262.9495, 262.9548, 262.9599, 262.9709, 262.9833, 263.0005, 263.0129, 
    263.0212, 263.0161, 263.0206, 263.0156, 263.0133, 263.0393, 263.0247, 
    263.0466, 263.0454, 263.0355, 263.0456, 262.9469, 262.944, 262.934, 
    262.9418, 262.9276, 262.9355, 262.9401, 262.9577, 262.9616, 262.9652, 
    262.9723, 262.9813, 262.9972, 263.011, 263.0236, 263.0226, 263.0229, 
    263.0258, 263.0188, 263.0269, 263.0282, 263.0247, 263.0453, 263.0394, 
    263.0454, 263.0416, 262.9449, 262.9497, 262.9471, 262.952, 262.9486, 
    262.9639, 262.9685, 262.9899, 262.9811, 262.9951, 262.9826, 262.9848, 
    262.9955, 262.9832, 263.0102, 262.9919, 263.0258, 263.0076, 263.027, 
    263.0235, 263.0293, 263.0345, 263.041, 263.0531, 263.0503, 263.0604, 
    262.9569, 262.9632, 262.9626, 262.9691, 262.974, 262.9844, 263.0011, 
    262.9949, 263.0064, 263.0087, 262.9912, 263.0019, 262.9673, 262.9729, 
    262.9696, 262.9574, 262.9963, 262.9763, 263.0132, 263.0024, 263.0338, 
    263.0182, 263.0488, 263.0618, 263.074, 263.0882, 262.9666, 262.9623, 
    262.9699, 262.9804, 262.9901, 263.003, 263.0044, 263.0068, 263.013, 
    263.0183, 263.0075, 263.0196, 262.9742, 262.998, 262.9607, 262.972, 
    262.9798, 262.9763, 262.9941, 262.9983, 263.0153, 263.0065, 263.0586, 
    263.0356, 263.099, 263.0814, 262.9608, 262.9666, 262.9864, 262.977, 
    263.0039, 263.0105, 263.0159, 263.0227, 263.0235, 263.0276, 263.0209, 
    263.0273, 263.0031, 263.0139, 262.9841, 262.9914, 262.988, 262.9844, 
    262.9957, 263.0077, 263.008, 263.0118, 263.0226, 263.004, 263.0615, 
    263.026, 262.9728, 262.9837, 262.9853, 262.9811, 263.0098, 262.9994, 
    263.0274, 263.0199, 263.0323, 263.0261, 263.0252, 263.0173, 263.0124, 
    262.9999, 262.9897, 262.9817, 262.9836, 262.9924, 263.0084, 263.0236, 
    263.0202, 263.0313, 263.002, 263.0143, 263.0095, 263.0219, 262.9947, 
    263.0178, 262.9888, 262.9913, 262.9992, 263.0151, 263.0186, 263.0224, 
    263.0201, 263.0088, 263.007, 262.999, 262.9968, 262.9908, 262.9857, 
    262.9903, 262.9951, 263.0089, 263.0211, 263.0346, 263.0379, 263.0534, 
    263.0407, 263.0617, 263.0438, 263.0746, 263.0192, 263.0433, 262.9996, 
    263.0043, 263.0128, 263.0324, 263.0219, 263.0342, 263.0069, 262.9927, 
    262.989, 262.9822, 262.9892, 262.9886, 262.9954, 262.9932, 263.0093, 
    263.0006, 263.0252, 263.0341, 263.0593, 263.0746, 263.0902, 263.097, 
    263.0991, 263.1 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9051, 253.9059, 253.9058, 253.9064, 253.9061, 253.9065, 253.9053, 
    253.906, 253.9055, 253.9052, 253.9077, 253.9065, 253.9091, 253.9083, 
    253.9104, 253.909, 253.9107, 253.9104, 253.9113, 253.911, 253.9122, 
    253.9115, 253.9129, 253.9121, 253.9122, 253.9114, 253.9067, 253.9076, 
    253.9067, 253.9068, 253.9068, 253.9061, 253.9057, 253.905, 253.9052, 
    253.9057, 253.9069, 253.9065, 253.9075, 253.9075, 253.9086, 253.9081, 
    253.91, 253.9095, 253.9111, 253.9107, 253.911, 253.9109, 253.911, 
    253.9104, 253.9107, 253.9102, 253.9082, 253.9088, 253.907, 253.906, 
    253.9053, 253.9048, 253.9049, 253.905, 253.9057, 253.9063, 253.9068, 
    253.9072, 253.9075, 253.9084, 253.909, 253.9101, 253.9099, 253.9103, 
    253.9106, 253.9112, 253.9111, 253.9113, 253.9103, 253.911, 253.9098, 
    253.9101, 253.9075, 253.9066, 253.9061, 253.9058, 253.9049, 253.9055, 
    253.9053, 253.9059, 253.9062, 253.9061, 253.9072, 253.9067, 253.909, 
    253.908, 253.9106, 253.91, 253.9107, 253.9103, 253.911, 253.9104, 
    253.9114, 253.9117, 253.9115, 253.9121, 253.9104, 253.911, 253.906, 
    253.9061, 253.9062, 253.9056, 253.9056, 253.905, 253.9055, 253.9057, 
    253.9062, 253.9066, 253.9069, 253.9075, 253.9082, 253.9093, 253.91, 
    253.9105, 253.9102, 253.9105, 253.9102, 253.91, 253.9116, 253.9107, 
    253.912, 253.9119, 253.9113, 253.912, 253.9061, 253.9059, 253.9053, 
    253.9058, 253.905, 253.9054, 253.9057, 253.9067, 253.907, 253.9072, 
    253.9076, 253.9081, 253.9091, 253.9099, 253.9106, 253.9106, 253.9106, 
    253.9108, 253.9104, 253.9108, 253.9109, 253.9107, 253.9119, 253.9116, 
    253.9119, 253.9117, 253.906, 253.9063, 253.9061, 253.9064, 253.9062, 
    253.9071, 253.9073, 253.9086, 253.9081, 253.9089, 253.9082, 253.9083, 
    253.9089, 253.9082, 253.9098, 253.9087, 253.9108, 253.9097, 253.9108, 
    253.9106, 253.911, 253.9113, 253.9117, 253.9124, 253.9122, 253.9128, 
    253.9067, 253.907, 253.907, 253.9074, 253.9077, 253.9083, 253.9093, 
    253.9089, 253.9096, 253.9097, 253.9087, 253.9093, 253.9073, 253.9076, 
    253.9074, 253.9067, 253.909, 253.9078, 253.91, 253.9094, 253.9112, 
    253.9103, 253.9121, 253.9129, 253.9137, 253.9145, 253.9072, 253.907, 
    253.9075, 253.9081, 253.9086, 253.9094, 253.9095, 253.9096, 253.91, 
    253.9103, 253.9097, 253.9104, 253.9077, 253.9091, 253.9069, 253.9075, 
    253.908, 253.9078, 253.9089, 253.9091, 253.9101, 253.9096, 253.9127, 
    253.9113, 253.9152, 253.9141, 253.9069, 253.9073, 253.9084, 253.9079, 
    253.9095, 253.9099, 253.9102, 253.9106, 253.9106, 253.9109, 253.9105, 
    253.9109, 253.9094, 253.9101, 253.9083, 253.9087, 253.9085, 253.9083, 
    253.909, 253.9097, 253.9097, 253.9099, 253.9105, 253.9095, 253.9129, 
    253.9107, 253.9076, 253.9082, 253.9084, 253.9081, 253.9098, 253.9092, 
    253.9109, 253.9104, 253.9112, 253.9108, 253.9107, 253.9103, 253.91, 
    253.9092, 253.9086, 253.9081, 253.9083, 253.9088, 253.9097, 253.9106, 
    253.9104, 253.9111, 253.9093, 253.9101, 253.9098, 253.9105, 253.9089, 
    253.9102, 253.9086, 253.9087, 253.9092, 253.9101, 253.9103, 253.9106, 
    253.9104, 253.9097, 253.9096, 253.9092, 253.909, 253.9087, 253.9084, 
    253.9087, 253.9089, 253.9098, 253.9105, 253.9113, 253.9115, 253.9124, 
    253.9116, 253.9129, 253.9118, 253.9137, 253.9103, 253.9118, 253.9092, 
    253.9095, 253.91, 253.9111, 253.9105, 253.9113, 253.9096, 253.9088, 
    253.9086, 253.9082, 253.9086, 253.9086, 253.909, 253.9088, 253.9098, 
    253.9093, 253.9107, 253.9113, 253.9128, 253.9137, 253.9147, 253.9151, 
    253.9152, 253.9153 ;

 TWS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 T_SCALAR =
  0.1400014, 0.1400093, 0.1400078, 0.1400141, 0.1400107, 0.1400147, 
    0.1400031, 0.1400096, 0.1400055, 0.1400022, 0.1400261, 0.1400144, 
    0.140039, 0.1400314, 0.1400508, 0.1400377, 0.1400534, 0.1400505, 
    0.1400596, 0.140057, 0.1400684, 0.1400608, 0.1400745, 0.1400666, 
    0.1400678, 0.1400606, 0.1400169, 0.1400246, 0.1400164, 0.1400175, 
    0.140017, 0.1400107, 0.1400074, 0.1400009, 0.1400021, 0.1400069, 
    0.140018, 0.1400143, 0.1400239, 0.1400237, 0.1400342, 0.1400295, 
    0.1400474, 0.1400423, 0.1400571, 0.1400534, 0.1400569, 0.1400559, 
    0.140057, 0.1400515, 0.1400538, 0.140049, 0.1400303, 0.1400357, 
    0.1400195, 0.1400095, 0.1400033, 0.1399988, 0.1399995, 0.1400006, 
    0.1400069, 0.140013, 0.1400176, 0.1400206, 0.1400236, 0.1400324, 
    0.1400374, 0.1400483, 0.1400465, 0.1400497, 0.140053, 0.1400584, 
    0.1400575, 0.1400598, 0.1400497, 0.1400564, 0.1400454, 0.1400484, 
    0.1400239, 0.1400153, 0.1400112, 0.1400081, 0.1399999, 0.1400055, 
    0.1400033, 0.1400087, 0.140012, 0.1400104, 0.1400207, 0.1400167, 
    0.1400377, 0.1400286, 0.1400526, 0.1400469, 0.140054, 0.1400504, 
    0.1400566, 0.140051, 0.1400607, 0.1400628, 0.1400614, 0.140067, 
    0.1400507, 0.1400569, 0.1400103, 0.1400106, 0.1400119, 0.1400062, 
    0.1400059, 0.1400009, 0.1400054, 0.1400073, 0.1400123, 0.1400151, 
    0.1400179, 0.140024, 0.1400307, 0.1400403, 0.1400473, 0.1400519, 
    0.1400491, 0.1400516, 0.1400488, 0.1400475, 0.140062, 0.1400538, 
    0.1400662, 0.1400655, 0.1400599, 0.1400656, 0.1400108, 0.1400093, 
    0.1400038, 0.1400081, 0.1400003, 0.1400046, 0.140007, 0.1400166, 
    0.1400189, 0.1400208, 0.1400247, 0.1400297, 0.1400384, 0.1400461, 
    0.1400532, 0.1400527, 0.1400529, 0.1400544, 0.1400505, 0.1400551, 
    0.1400558, 0.1400539, 0.1400654, 0.1400621, 0.1400655, 0.1400634, 
    0.1400098, 0.1400124, 0.140011, 0.1400136, 0.1400117, 0.14002, 0.1400225, 
    0.1400343, 0.1400296, 0.1400373, 0.1400304, 0.1400316, 0.1400373, 
    0.1400308, 0.1400456, 0.1400353, 0.1400545, 0.140044, 0.1400551, 
    0.1400532, 0.1400565, 0.1400593, 0.140063, 0.1400697, 0.1400682, 
    0.1400739, 0.1400163, 0.1400196, 0.1400194, 0.140023, 0.1400256, 
    0.1400314, 0.1400407, 0.1400372, 0.1400436, 0.1400449, 0.1400352, 
    0.1400411, 0.140022, 0.1400249, 0.1400232, 0.1400165, 0.1400379, 
    0.1400268, 0.1400474, 0.1400414, 0.1400589, 0.1400501, 0.1400673, 
    0.1400745, 0.1400817, 0.1400897, 0.1400216, 0.1400193, 0.1400235, 
    0.1400291, 0.1400346, 0.1400417, 0.1400425, 0.1400438, 0.1400473, 
    0.1400503, 0.1400441, 0.140051, 0.1400254, 0.1400389, 0.1400183, 
    0.1400244, 0.1400288, 0.1400269, 0.1400369, 0.1400391, 0.1400485, 
    0.1400437, 0.1400726, 0.1400598, 0.1400961, 0.1400858, 0.1400185, 
    0.1400216, 0.1400324, 0.1400273, 0.1400422, 0.1400459, 0.140049, 
    0.1400527, 0.1400532, 0.1400554, 0.1400517, 0.1400553, 0.1400417, 
    0.1400478, 0.1400313, 0.1400352, 0.1400335, 0.1400314, 0.1400377, 
    0.1400442, 0.1400445, 0.1400466, 0.1400521, 0.1400423, 0.140074, 
    0.1400541, 0.140025, 0.1400309, 0.1400319, 0.1400296, 0.1400455, 
    0.1400397, 0.1400554, 0.1400512, 0.1400581, 0.1400547, 0.1400541, 
    0.1400497, 0.1400469, 0.14004, 0.1400343, 0.14003, 0.140031, 0.1400358, 
    0.1400446, 0.1400532, 0.1400513, 0.1400576, 0.1400411, 0.1400479, 
    0.1400453, 0.1400523, 0.1400371, 0.1400495, 0.1400339, 0.1400353, 
    0.1400396, 0.1400483, 0.1400505, 0.1400525, 0.1400513, 0.1400449, 
    0.1400439, 0.1400395, 0.1400383, 0.140035, 0.1400322, 0.1400347, 
    0.1400373, 0.140045, 0.1400518, 0.1400593, 0.1400613, 0.1400697, 
    0.1400626, 0.1400741, 0.140064, 0.1400817, 0.1400505, 0.140064, 
    0.1400399, 0.1400425, 0.1400471, 0.140058, 0.1400523, 0.140059, 
    0.1400439, 0.1400359, 0.140034, 0.1400302, 0.1400341, 0.1400338, 
    0.1400375, 0.1400363, 0.1400452, 0.1400404, 0.1400541, 0.140059, 
    0.1400733, 0.1400819, 0.140091, 0.140095, 0.1400962, 0.1400967,
  0.1463853, 0.146394, 0.1463923, 0.1463993, 0.1463955, 0.1464, 0.1463871, 
    0.1463943, 0.1463897, 0.1463861, 0.1464126, 0.1463996, 0.1464269, 
    0.1464184, 0.14644, 0.1464255, 0.146443, 0.1464398, 0.1464499, 0.146447, 
    0.1464596, 0.1464512, 0.1464665, 0.1464577, 0.146459, 0.1464509, 
    0.1464024, 0.1464109, 0.1464018, 0.1464031, 0.1464025, 0.1463955, 
    0.1463918, 0.1463847, 0.146386, 0.1463913, 0.1464036, 0.1463995, 
    0.1464101, 0.1464099, 0.1464216, 0.1464163, 0.1464363, 0.1464306, 
    0.1464471, 0.1464429, 0.1464469, 0.1464457, 0.1464469, 0.1464408, 
    0.1464434, 0.146438, 0.1464173, 0.1464233, 0.1464053, 0.1463943, 
    0.1463874, 0.1463824, 0.1463831, 0.1463844, 0.1463914, 0.1463981, 
    0.1464031, 0.1464065, 0.1464099, 0.1464196, 0.1464251, 0.1464373, 
    0.1464353, 0.1464389, 0.1464425, 0.1464485, 0.1464475, 0.1464501, 
    0.1464389, 0.1464463, 0.1464341, 0.1464374, 0.1464102, 0.1464007, 
    0.1463961, 0.1463926, 0.1463836, 0.1463898, 0.1463874, 0.1463933, 
    0.146397, 0.1463952, 0.1464066, 0.1464021, 0.1464255, 0.1464154, 
    0.1464421, 0.1464357, 0.1464436, 0.1464396, 0.1464465, 0.1464403, 
    0.1464511, 0.1464534, 0.1464518, 0.1464581, 0.1464399, 0.1464468, 
    0.1463951, 0.1463954, 0.1463968, 0.1463906, 0.1463902, 0.1463846, 
    0.1463896, 0.1463917, 0.1463973, 0.1464004, 0.1464035, 0.1464102, 
    0.1464177, 0.1464283, 0.1464361, 0.1464413, 0.1464381, 0.1464409, 
    0.1464378, 0.1464364, 0.1464525, 0.1464434, 0.1464572, 0.1464564, 
    0.1464501, 0.1464565, 0.1463956, 0.1463939, 0.1463879, 0.1463926, 
    0.146384, 0.1463888, 0.1463914, 0.1464021, 0.1464046, 0.1464067, 
    0.1464111, 0.1464166, 0.1464263, 0.1464348, 0.1464427, 0.1464422, 
    0.1464424, 0.1464441, 0.1464398, 0.1464448, 0.1464456, 0.1464434, 
    0.1464563, 0.1464527, 0.1464564, 0.146454, 0.1463945, 0.1463974, 
    0.1463958, 0.1463987, 0.1463966, 0.1464058, 0.1464086, 0.1464217, 
    0.1464165, 0.146425, 0.1464174, 0.1464187, 0.146425, 0.1464178, 
    0.1464342, 0.1464229, 0.1464442, 0.1464325, 0.1464449, 0.1464427, 
    0.1464463, 0.1464495, 0.1464537, 0.1464612, 0.1464594, 0.1464658, 
    0.1464017, 0.1464054, 0.1464052, 0.1464092, 0.1464121, 0.1464185, 
    0.1464288, 0.1464249, 0.1464321, 0.1464335, 0.1464227, 0.1464292, 
    0.146408, 0.1464113, 0.1464094, 0.146402, 0.1464257, 0.1464134, 
    0.1464362, 0.1464295, 0.1464491, 0.1464392, 0.1464585, 0.1464665, 
    0.1464746, 0.1464834, 0.1464076, 0.146405, 0.1464097, 0.1464159, 
    0.146422, 0.1464299, 0.1464308, 0.1464323, 0.1464362, 0.1464394, 
    0.1464326, 0.1464403, 0.1464119, 0.1464268, 0.146404, 0.1464107, 
    0.1464156, 0.1464135, 0.1464245, 0.1464271, 0.1464375, 0.1464322, 
    0.1464644, 0.1464501, 0.1464906, 0.1464791, 0.1464041, 0.1464076, 
    0.1464196, 0.1464139, 0.1464305, 0.1464346, 0.146438, 0.1464422, 
    0.1464427, 0.1464452, 0.1464411, 0.1464451, 0.1464299, 0.1464367, 
    0.1464184, 0.1464227, 0.1464208, 0.1464185, 0.1464255, 0.1464327, 
    0.146433, 0.1464353, 0.1464415, 0.1464306, 0.146466, 0.1464438, 
    0.1464114, 0.1464179, 0.146419, 0.1464165, 0.1464342, 0.1464277, 
    0.1464451, 0.1464405, 0.1464482, 0.1464443, 0.1464438, 0.1464389, 
    0.1464358, 0.146428, 0.1464217, 0.1464169, 0.146418, 0.1464234, 
    0.1464332, 0.1464427, 0.1464406, 0.1464476, 0.1464293, 0.1464369, 
    0.1464339, 0.1464417, 0.1464248, 0.1464387, 0.1464212, 0.1464228, 
    0.1464276, 0.1464373, 0.1464397, 0.1464419, 0.1464406, 0.1464335, 
    0.1464324, 0.1464275, 0.1464261, 0.1464224, 0.1464193, 0.1464221, 
    0.146425, 0.1464335, 0.1464412, 0.1464496, 0.1464517, 0.1464611, 
    0.1464532, 0.1464661, 0.1464548, 0.1464745, 0.1464397, 0.1464548, 
    0.1464279, 0.1464308, 0.1464359, 0.1464481, 0.1464417, 0.1464492, 
    0.1464324, 0.1464235, 0.1464214, 0.1464171, 0.1464215, 0.1464211, 
    0.1464253, 0.1464239, 0.1464338, 0.1464285, 0.1464437, 0.1464492, 
    0.1464651, 0.1464748, 0.146485, 0.1464894, 0.1464907, 0.1464913,
  0.1561714, 0.1561798, 0.1561782, 0.1561849, 0.1561813, 0.1561856, 
    0.1561732, 0.1561801, 0.1561757, 0.1561723, 0.1561978, 0.1561852, 
    0.1562117, 0.1562034, 0.1562244, 0.1562103, 0.1562273, 0.1562242, 
    0.156234, 0.1562312, 0.1562436, 0.1562353, 0.1562503, 0.1562417, 
    0.156243, 0.1562351, 0.1561879, 0.1561962, 0.1561874, 0.1561886, 
    0.1561881, 0.1561813, 0.1561778, 0.1561709, 0.1561722, 0.1561773, 
    0.1561891, 0.1561852, 0.1561954, 0.1561952, 0.1562065, 0.1562014, 
    0.1562207, 0.1562153, 0.1562313, 0.1562272, 0.1562311, 0.15623, 
    0.1562311, 0.1562252, 0.1562277, 0.1562225, 0.1562023, 0.1562082, 
    0.1561907, 0.1561801, 0.1561735, 0.1561687, 0.1561694, 0.1561706, 
    0.1561773, 0.1561837, 0.1561886, 0.1561919, 0.1561951, 0.1562046, 
    0.15621, 0.1562218, 0.1562198, 0.1562233, 0.1562268, 0.1562327, 
    0.1562317, 0.1562342, 0.1562233, 0.1562305, 0.1562186, 0.1562218, 
    0.1561955, 0.1561863, 0.1561819, 0.1561785, 0.1561699, 0.1561758, 
    0.1561734, 0.1561792, 0.1561827, 0.156181, 0.156192, 0.1561877, 
    0.1562103, 0.1562005, 0.1562264, 0.1562202, 0.1562279, 0.156224, 
    0.1562307, 0.1562247, 0.1562352, 0.1562375, 0.1562359, 0.1562421, 
    0.1562243, 0.1562311, 0.1561809, 0.1561812, 0.1561826, 0.1561765, 
    0.1561762, 0.1561708, 0.1561756, 0.1561777, 0.156183, 0.156186, 0.156189, 
    0.1561955, 0.1562027, 0.156213, 0.1562206, 0.1562257, 0.1562226, 
    0.1562253, 0.1562223, 0.1562209, 0.1562366, 0.1562277, 0.1562412, 
    0.1562405, 0.1562343, 0.1562405, 0.1561814, 0.1561798, 0.1561739, 
    0.1561785, 0.1561703, 0.1561748, 0.1561774, 0.1561877, 0.1561901, 
    0.1561921, 0.1561963, 0.1562017, 0.156211, 0.1562194, 0.1562271, 
    0.1562265, 0.1562267, 0.1562284, 0.1562242, 0.1562291, 0.1562299, 
    0.1562278, 0.1562404, 0.1562368, 0.1562404, 0.1562381, 0.1561803, 
    0.1561831, 0.1561816, 0.1561844, 0.1561824, 0.1561912, 0.1561939, 
    0.1562066, 0.1562015, 0.1562098, 0.1562024, 0.1562037, 0.1562098, 
    0.1562028, 0.1562188, 0.1562078, 0.1562285, 0.1562171, 0.1562292, 
    0.156227, 0.1562306, 0.1562337, 0.1562378, 0.1562451, 0.1562434, 
    0.1562496, 0.1561873, 0.1561909, 0.1561906, 0.1561945, 0.1561973, 
    0.1562035, 0.1562135, 0.1562097, 0.1562167, 0.1562181, 0.1562076, 
    0.1562139, 0.1561933, 0.1561965, 0.1561947, 0.1561875, 0.1562105, 
    0.1561986, 0.1562207, 0.1562142, 0.1562333, 0.1562237, 0.1562425, 
    0.1562503, 0.1562582, 0.156267, 0.1561929, 0.1561905, 0.156195, 0.156201, 
    0.1562069, 0.1562146, 0.1562154, 0.1562169, 0.1562207, 0.1562239, 
    0.1562172, 0.1562247, 0.1561971, 0.1562115, 0.1561895, 0.1561959, 
    0.1562007, 0.1561987, 0.1562093, 0.1562118, 0.156222, 0.1562168, 
    0.1562483, 0.1562342, 0.156274, 0.1562627, 0.1561896, 0.156193, 
    0.1562046, 0.1561991, 0.1562152, 0.1562191, 0.1562224, 0.1562265, 
    0.156227, 0.1562295, 0.1562255, 0.1562293, 0.1562146, 0.1562212, 
    0.1562034, 0.1562076, 0.1562057, 0.1562035, 0.1562103, 0.1562173, 
    0.1562176, 0.1562199, 0.1562259, 0.1562152, 0.1562498, 0.1562281, 
    0.1561966, 0.1562029, 0.156204, 0.1562015, 0.1562187, 0.1562124, 
    0.1562294, 0.1562248, 0.1562324, 0.1562286, 0.1562281, 0.1562233, 
    0.1562203, 0.1562127, 0.1562066, 0.1562019, 0.156203, 0.1562082, 
    0.1562178, 0.156227, 0.156225, 0.1562318, 0.156214, 0.1562214, 0.1562185, 
    0.1562261, 0.1562096, 0.1562231, 0.1562061, 0.1562076, 0.1562123, 
    0.1562217, 0.1562241, 0.1562263, 0.156225, 0.1562181, 0.156217, 
    0.1562123, 0.1562109, 0.1562073, 0.1562043, 0.156207, 0.1562098, 
    0.1562181, 0.1562255, 0.1562337, 0.1562358, 0.1562451, 0.1562373, 
    0.1562499, 0.1562389, 0.1562582, 0.1562242, 0.1562389, 0.1562126, 
    0.1562154, 0.1562204, 0.1562323, 0.156226, 0.1562334, 0.156217, 
    0.1562083, 0.1562063, 0.1562022, 0.1562064, 0.156206, 0.1562101, 
    0.1562088, 0.1562184, 0.1562132, 0.156228, 0.1562334, 0.1562489, 
    0.1562584, 0.1562685, 0.1562728, 0.1562742, 0.1562747,
  0.1699164, 0.1699228, 0.1699216, 0.1699268, 0.1699239, 0.1699273, 
    0.1699177, 0.169923, 0.1699197, 0.169917, 0.1699368, 0.169927, 0.1699477, 
    0.1699412, 0.1699577, 0.1699466, 0.16996, 0.1699575, 0.1699654, 
    0.1699631, 0.169973, 0.1699664, 0.1699784, 0.1699715, 0.1699725, 
    0.1699662, 0.1699291, 0.1699356, 0.1699287, 0.1699296, 0.1699292, 
    0.169924, 0.1699212, 0.169916, 0.1699169, 0.1699209, 0.16993, 0.169927, 
    0.1699349, 0.1699348, 0.1699436, 0.1699396, 0.1699549, 0.1699505, 
    0.1699632, 0.16996, 0.1699631, 0.1699621, 0.1699631, 0.1699583, 
    0.1699603, 0.1699562, 0.1699404, 0.1699449, 0.1699313, 0.1699231, 
    0.1699179, 0.1699142, 0.1699148, 0.1699157, 0.1699209, 0.1699259, 
    0.1699297, 0.1699322, 0.1699347, 0.1699421, 0.1699463, 0.1699557, 
    0.1699541, 0.1699569, 0.1699597, 0.1699643, 0.1699635, 0.1699656, 
    0.1699569, 0.1699626, 0.1699532, 0.1699557, 0.169935, 0.1699278, 
    0.1699245, 0.1699218, 0.1699152, 0.1699197, 0.1699179, 0.1699223, 
    0.1699251, 0.1699237, 0.1699323, 0.1699289, 0.1699466, 0.1699389, 
    0.1699593, 0.1699544, 0.1699605, 0.1699574, 0.1699627, 0.169958, 
    0.1699663, 0.1699681, 0.1699669, 0.1699718, 0.1699577, 0.169963, 
    0.1699237, 0.1699239, 0.169925, 0.1699203, 0.16992, 0.1699159, 0.1699196, 
    0.1699212, 0.1699253, 0.1699277, 0.16993, 0.169935, 0.1699407, 0.1699488, 
    0.1699547, 0.1699587, 0.1699563, 0.1699584, 0.169956, 0.1699549, 
    0.1699674, 0.1699603, 0.1699711, 0.1699705, 0.1699656, 0.1699706, 
    0.1699241, 0.1699228, 0.1699183, 0.1699218, 0.1699155, 0.169919, 
    0.169921, 0.1699289, 0.1699308, 0.1699324, 0.1699356, 0.1699398, 
    0.1699472, 0.1699537, 0.1699599, 0.1699594, 0.1699596, 0.1699609, 
    0.1699575, 0.1699614, 0.1699621, 0.1699604, 0.1699704, 0.1699675, 
    0.1699705, 0.1699686, 0.1699232, 0.1699254, 0.1699242, 0.1699264, 
    0.1699248, 0.1699317, 0.1699338, 0.1699437, 0.1699397, 0.1699462, 
    0.1699404, 0.1699414, 0.1699463, 0.1699408, 0.1699533, 0.1699446, 
    0.1699609, 0.169952, 0.1699615, 0.1699598, 0.1699626, 0.1699651, 
    0.1699683, 0.1699742, 0.1699729, 0.1699778, 0.1699286, 0.1699314, 
    0.1699312, 0.1699342, 0.1699364, 0.1699413, 0.1699491, 0.1699462, 
    0.1699516, 0.1699527, 0.1699445, 0.1699494, 0.1699333, 0.1699358, 
    0.1699344, 0.1699288, 0.1699467, 0.1699374, 0.1699548, 0.1699497, 
    0.1699648, 0.1699571, 0.1699721, 0.1699784, 0.1699847, 0.1699918, 
    0.169933, 0.1699311, 0.1699346, 0.1699393, 0.1699439, 0.16995, 0.1699507, 
    0.1699518, 0.1699548, 0.1699573, 0.1699521, 0.1699579, 0.1699363, 
    0.1699476, 0.1699303, 0.1699354, 0.1699391, 0.1699375, 0.1699459, 
    0.1699478, 0.1699558, 0.1699517, 0.1699768, 0.1699656, 0.1699975, 
    0.1699884, 0.1699304, 0.169933, 0.1699421, 0.1699378, 0.1699504, 
    0.1699536, 0.1699562, 0.1699594, 0.1699598, 0.1699618, 0.1699586, 
    0.1699616, 0.16995, 0.1699552, 0.1699412, 0.1699445, 0.169943, 0.1699413, 
    0.1699466, 0.1699521, 0.1699524, 0.1699542, 0.1699589, 0.1699505, 
    0.169978, 0.1699607, 0.1699359, 0.1699408, 0.1699417, 0.1699397, 
    0.1699532, 0.1699483, 0.1699617, 0.1699581, 0.1699641, 0.1699611, 
    0.1699606, 0.1699568, 0.1699545, 0.1699485, 0.1699437, 0.16994, 
    0.1699409, 0.169945, 0.1699525, 0.1699598, 0.1699582, 0.1699636, 
    0.1699495, 0.1699553, 0.169953, 0.1699591, 0.1699461, 0.1699567, 
    0.1699433, 0.1699445, 0.1699482, 0.1699556, 0.1699575, 0.1699592, 
    0.1699582, 0.1699527, 0.1699519, 0.1699481, 0.1699471, 0.1699443, 
    0.1699419, 0.169944, 0.1699463, 0.1699528, 0.1699586, 0.1699651, 
    0.1699668, 0.1699742, 0.169968, 0.1699781, 0.1699693, 0.1699847, 
    0.1699575, 0.1699692, 0.1699484, 0.1699506, 0.1699546, 0.169964, 
    0.169959, 0.1699649, 0.1699519, 0.1699451, 0.1699435, 0.1699402, 
    0.1699435, 0.1699433, 0.1699464, 0.1699454, 0.169953, 0.1699489, 
    0.1699606, 0.1699649, 0.1699773, 0.1699849, 0.169993, 0.1699965, 
    0.1699976, 0.169998,
  0.1852159, 0.1852192, 0.1852185, 0.1852212, 0.1852197, 0.1852214, 
    0.1852166, 0.1852193, 0.1852176, 0.1852162, 0.1852263, 0.1852213, 
    0.185232, 0.1852286, 0.1852373, 0.1852314, 0.1852386, 0.1852372, 
    0.1852414, 0.1852402, 0.1852455, 0.185242, 0.1852484, 0.1852447, 
    0.1852453, 0.1852418, 0.1852224, 0.1852257, 0.1852222, 0.1852226, 
    0.1852224, 0.1852197, 0.1852183, 0.1852157, 0.1852162, 0.1852182, 
    0.1852228, 0.1852213, 0.1852254, 0.1852253, 0.1852299, 0.1852278, 
    0.1852358, 0.1852335, 0.1852403, 0.1852385, 0.1852402, 0.1852397, 
    0.1852402, 0.1852376, 0.1852387, 0.1852365, 0.1852282, 0.1852306, 
    0.1852235, 0.1852193, 0.1852167, 0.1852148, 0.1852151, 0.1852156, 
    0.1852182, 0.1852207, 0.1852227, 0.185224, 0.1852253, 0.1852291, 
    0.1852313, 0.1852362, 0.1852354, 0.1852369, 0.1852384, 0.1852408, 
    0.1852404, 0.1852415, 0.1852369, 0.1852399, 0.1852349, 0.1852362, 
    0.1852254, 0.1852217, 0.18522, 0.1852186, 0.1852153, 0.1852176, 
    0.1852167, 0.1852189, 0.1852203, 0.1852196, 0.185224, 0.1852223, 
    0.1852314, 0.1852274, 0.1852382, 0.1852356, 0.1852388, 0.1852372, 
    0.18524, 0.1852375, 0.1852419, 0.1852429, 0.1852422, 0.1852449, 
    0.1852373, 0.1852401, 0.1852196, 0.1852197, 0.1852202, 0.1852179, 
    0.1852177, 0.1852157, 0.1852175, 0.1852183, 0.1852204, 0.1852216, 
    0.1852228, 0.1852254, 0.1852283, 0.1852326, 0.1852357, 0.1852379, 
    0.1852366, 0.1852377, 0.1852364, 0.1852358, 0.1852425, 0.1852387, 
    0.1852445, 0.1852442, 0.1852415, 0.1852442, 0.1852198, 0.1852192, 
    0.1852169, 0.1852186, 0.1852154, 0.1852172, 0.1852182, 0.1852223, 
    0.1852232, 0.185224, 0.1852257, 0.1852279, 0.1852318, 0.1852352, 
    0.1852385, 0.1852382, 0.1852383, 0.185239, 0.1852372, 0.1852393, 
    0.1852396, 0.1852387, 0.1852441, 0.1852426, 0.1852442, 0.1852432, 
    0.1852194, 0.1852205, 0.1852199, 0.185221, 0.1852202, 0.1852237, 
    0.1852248, 0.1852299, 0.1852279, 0.1852312, 0.1852282, 0.1852287, 
    0.1852313, 0.1852284, 0.185235, 0.1852304, 0.185239, 0.1852343, 
    0.1852393, 0.1852384, 0.1852399, 0.1852413, 0.185243, 0.1852462, 
    0.1852455, 0.1852482, 0.1852221, 0.1852235, 0.1852235, 0.185225, 
    0.1852261, 0.1852287, 0.1852328, 0.1852312, 0.1852341, 0.1852347, 
    0.1852303, 0.1852329, 0.1852245, 0.1852258, 0.1852251, 0.1852222, 
    0.1852315, 0.1852267, 0.1852358, 0.1852331, 0.1852411, 0.185237, 
    0.185245, 0.1852485, 0.1852519, 0.1852558, 0.1852244, 0.1852234, 
    0.1852252, 0.1852276, 0.18523, 0.1852332, 0.1852336, 0.1852342, 
    0.1852358, 0.1852371, 0.1852343, 0.1852374, 0.1852261, 0.185232, 
    0.185223, 0.1852256, 0.1852275, 0.1852267, 0.1852311, 0.1852321, 
    0.1852363, 0.1852341, 0.1852476, 0.1852415, 0.185259, 0.1852539, 
    0.185223, 0.1852244, 0.1852291, 0.1852268, 0.1852335, 0.1852351, 
    0.1852365, 0.1852382, 0.1852384, 0.1852395, 0.1852378, 0.1852394, 
    0.1852332, 0.185236, 0.1852286, 0.1852303, 0.1852296, 0.1852287, 
    0.1852314, 0.1852344, 0.1852345, 0.1852354, 0.185238, 0.1852335, 
    0.1852482, 0.1852389, 0.1852259, 0.1852284, 0.1852289, 0.1852279, 
    0.1852349, 0.1852323, 0.1852394, 0.1852375, 0.1852407, 0.1852391, 
    0.1852389, 0.1852369, 0.1852356, 0.1852324, 0.1852299, 0.185228, 
    0.1852285, 0.1852306, 0.1852345, 0.1852384, 0.1852376, 0.1852405, 
    0.185233, 0.1852361, 0.1852348, 0.185238, 0.1852312, 0.1852368, 
    0.1852297, 0.1852303, 0.1852323, 0.1852362, 0.1852372, 0.1852381, 
    0.1852376, 0.1852347, 0.1852342, 0.1852323, 0.1852317, 0.1852302, 
    0.185229, 0.1852301, 0.1852313, 0.1852347, 0.1852378, 0.1852413, 
    0.1852422, 0.1852462, 0.1852428, 0.1852483, 0.1852435, 0.1852519, 
    0.1852372, 0.1852435, 0.1852324, 0.1852336, 0.1852357, 0.1852407, 
    0.185238, 0.1852411, 0.1852342, 0.1852306, 0.1852298, 0.1852281, 
    0.1852298, 0.1852297, 0.1852313, 0.1852308, 0.1852348, 0.1852327, 
    0.1852389, 0.1852411, 0.1852479, 0.185252, 0.1852565, 0.1852584, 
    0.185259, 0.1852593,
  0.1954502, 0.1954509, 0.1954508, 0.1954514, 0.1954511, 0.1954515, 
    0.1954503, 0.195451, 0.1954506, 0.1954502, 0.1954527, 0.1954515, 
    0.1954542, 0.1954533, 0.1954556, 0.195454, 0.1954559, 0.1954555, 
    0.1954566, 0.1954563, 0.1954578, 0.1954568, 0.1954586, 0.1954575, 
    0.1954577, 0.1954568, 0.1954517, 0.1954526, 0.1954517, 0.1954518, 
    0.1954518, 0.1954511, 0.1954508, 0.1954501, 0.1954502, 0.1954507, 
    0.1954519, 0.1954515, 0.1954525, 0.1954525, 0.1954536, 0.1954531, 
    0.1954551, 0.1954546, 0.1954563, 0.1954559, 0.1954563, 0.1954562, 
    0.1954563, 0.1954556, 0.1954559, 0.1954553, 0.1954532, 0.1954538, 
    0.195452, 0.195451, 0.1954504, 0.1954499, 0.19545, 0.1954501, 0.1954507, 
    0.1954513, 0.1954518, 0.1954521, 0.1954525, 0.1954534, 0.195454, 
    0.1954553, 0.195455, 0.1954554, 0.1954558, 0.1954565, 0.1954564, 
    0.1954567, 0.1954554, 0.1954562, 0.1954549, 0.1954553, 0.1954525, 
    0.1954516, 0.1954512, 0.1954508, 0.19545, 0.1954506, 0.1954504, 
    0.1954509, 0.1954512, 0.1954511, 0.1954521, 0.1954517, 0.195454, 
    0.195453, 0.1954558, 0.1954551, 0.195456, 0.1954555, 0.1954563, 
    0.1954556, 0.1954568, 0.195457, 0.1954569, 0.1954576, 0.1954556, 
    0.1954563, 0.1954511, 0.1954511, 0.1954512, 0.1954506, 0.1954506, 
    0.1954501, 0.1954506, 0.1954508, 0.1954513, 0.1954516, 0.1954518, 
    0.1954525, 0.1954532, 0.1954543, 0.1954551, 0.1954557, 0.1954554, 
    0.1954557, 0.1954553, 0.1954552, 0.1954569, 0.1954559, 0.1954575, 
    0.1954574, 0.1954567, 0.1954574, 0.1954511, 0.1954509, 0.1954504, 
    0.1954508, 0.1954501, 0.1954505, 0.1954507, 0.1954517, 0.1954519, 
    0.1954522, 0.1954526, 0.1954531, 0.1954541, 0.195455, 0.1954558, 
    0.1954558, 0.1954558, 0.195456, 0.1954555, 0.1954561, 0.1954562, 
    0.1954559, 0.1954574, 0.195457, 0.1954574, 0.1954571, 0.195451, 
    0.1954513, 0.1954511, 0.1954514, 0.1954512, 0.1954521, 0.1954523, 
    0.1954536, 0.1954531, 0.195454, 0.1954532, 0.1954533, 0.195454, 
    0.1954532, 0.1954549, 0.1954537, 0.195456, 0.1954547, 0.1954561, 
    0.1954558, 0.1954563, 0.1954566, 0.1954571, 0.1954579, 0.1954577, 
    0.1954585, 0.1954517, 0.195452, 0.195452, 0.1954524, 0.1954527, 
    0.1954533, 0.1954544, 0.195454, 0.1954547, 0.1954549, 0.1954537, 
    0.1954544, 0.1954523, 0.1954526, 0.1954524, 0.1954517, 0.195454, 
    0.1954528, 0.1954551, 0.1954544, 0.1954565, 0.1954555, 0.1954576, 
    0.1954586, 0.1954595, 0.1954606, 0.1954522, 0.195452, 0.1954524, 
    0.195453, 0.1954537, 0.1954545, 0.1954546, 0.1954547, 0.1954551, 
    0.1954555, 0.1954548, 0.1954556, 0.1954526, 0.1954542, 0.1954519, 
    0.1954525, 0.195453, 0.1954528, 0.1954539, 0.1954542, 0.1954553, 
    0.1954547, 0.1954583, 0.1954567, 0.1954615, 0.1954601, 0.1954519, 
    0.1954522, 0.1954534, 0.1954529, 0.1954545, 0.195455, 0.1954553, 
    0.1954558, 0.1954558, 0.1954561, 0.1954557, 0.1954561, 0.1954545, 
    0.1954552, 0.1954533, 0.1954537, 0.1954535, 0.1954533, 0.195454, 
    0.1954548, 0.1954548, 0.195455, 0.1954557, 0.1954546, 0.1954585, 
    0.195456, 0.1954526, 0.1954532, 0.1954534, 0.1954531, 0.1954549, 
    0.1954543, 0.1954561, 0.1954556, 0.1954564, 0.195456, 0.195456, 
    0.1954554, 0.1954551, 0.1954543, 0.1954536, 0.1954531, 0.1954533, 
    0.1954538, 0.1954548, 0.1954558, 0.1954556, 0.1954564, 0.1954544, 
    0.1954552, 0.1954549, 0.1954557, 0.1954539, 0.1954554, 0.1954536, 
    0.1954537, 0.1954542, 0.1954553, 0.1954555, 0.1954558, 0.1954556, 
    0.1954549, 0.1954547, 0.1954542, 0.1954541, 0.1954537, 0.1954534, 
    0.1954537, 0.195454, 0.1954549, 0.1954557, 0.1954566, 0.1954568, 
    0.1954579, 0.195457, 0.1954585, 0.1954572, 0.1954595, 0.1954555, 
    0.1954572, 0.1954543, 0.1954546, 0.1954551, 0.1954564, 0.1954557, 
    0.1954566, 0.1954547, 0.1954538, 0.1954536, 0.1954532, 0.1954536, 
    0.1954536, 0.195454, 0.1954539, 0.1954549, 0.1954543, 0.195456, 
    0.1954566, 0.1954584, 0.1954596, 0.1954608, 0.1954614, 0.1954615, 
    0.1954616,
  0.1982628, 0.1982629, 0.1982629, 0.198263, 0.1982629, 0.198263, 0.1982629, 
    0.1982629, 0.1982629, 0.1982629, 0.1982631, 0.198263, 0.1982633, 
    0.1982632, 0.1982635, 0.1982633, 0.1982635, 0.1982635, 0.1982636, 
    0.1982636, 0.1982638, 0.1982637, 0.1982639, 0.1982637, 0.1982638, 
    0.1982637, 0.198263, 0.1982631, 0.198263, 0.198263, 0.198263, 0.1982629, 
    0.1982629, 0.1982628, 0.1982629, 0.1982629, 0.198263, 0.198263, 
    0.1982631, 0.1982631, 0.1982633, 0.1982632, 0.1982635, 0.1982634, 
    0.1982636, 0.1982635, 0.1982636, 0.1982636, 0.1982636, 0.1982635, 
    0.1982635, 0.1982635, 0.1982632, 0.1982633, 0.1982631, 0.1982629, 
    0.1982629, 0.1982628, 0.1982628, 0.1982628, 0.1982629, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982635, 
    0.1982634, 0.1982635, 0.1982635, 0.1982636, 0.1982636, 0.1982636, 
    0.1982635, 0.1982636, 0.1982634, 0.1982635, 0.1982631, 0.198263, 
    0.198263, 0.1982629, 0.1982628, 0.1982629, 0.1982629, 0.1982629, 
    0.198263, 0.1982629, 0.1982631, 0.198263, 0.1982633, 0.1982632, 
    0.1982635, 0.1982634, 0.1982635, 0.1982635, 0.1982636, 0.1982635, 
    0.1982637, 0.1982637, 0.1982637, 0.1982638, 0.1982635, 0.1982636, 
    0.1982629, 0.1982629, 0.198263, 0.1982629, 0.1982629, 0.1982628, 
    0.1982629, 0.1982629, 0.198263, 0.198263, 0.198263, 0.1982631, 0.1982632, 
    0.1982633, 0.1982634, 0.1982635, 0.1982635, 0.1982635, 0.1982635, 
    0.1982635, 0.1982637, 0.1982635, 0.1982637, 0.1982637, 0.1982636, 
    0.1982637, 0.198263, 0.1982629, 0.1982629, 0.1982629, 0.1982628, 
    0.1982629, 0.1982629, 0.198263, 0.198263, 0.1982631, 0.1982631, 
    0.1982632, 0.1982633, 0.1982634, 0.1982635, 0.1982635, 0.1982635, 
    0.1982636, 0.1982635, 0.1982636, 0.1982636, 0.1982635, 0.1982637, 
    0.1982637, 0.1982637, 0.1982637, 0.1982629, 0.198263, 0.198263, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982633, 0.1982632, 0.1982633, 
    0.1982632, 0.1982632, 0.1982633, 0.1982632, 0.1982634, 0.1982633, 
    0.1982636, 0.1982634, 0.1982636, 0.1982635, 0.1982636, 0.1982636, 
    0.1982637, 0.1982638, 0.1982638, 0.1982639, 0.198263, 0.1982631, 
    0.1982631, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982633, 
    0.1982634, 0.1982634, 0.1982633, 0.1982633, 0.1982631, 0.1982631, 
    0.1982631, 0.198263, 0.1982633, 0.1982632, 0.1982635, 0.1982634, 
    0.1982636, 0.1982635, 0.1982638, 0.1982639, 0.198264, 0.1982642, 
    0.1982631, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982634, 
    0.1982634, 0.1982634, 0.1982635, 0.1982635, 0.1982634, 0.1982635, 
    0.1982631, 0.1982633, 0.198263, 0.1982631, 0.1982632, 0.1982632, 
    0.1982633, 0.1982633, 0.1982635, 0.1982634, 0.1982639, 0.1982636, 
    0.1982643, 0.1982641, 0.198263, 0.1982631, 0.1982632, 0.1982632, 
    0.1982634, 0.1982634, 0.1982635, 0.1982635, 0.1982635, 0.1982636, 
    0.1982635, 0.1982636, 0.1982634, 0.1982635, 0.1982632, 0.1982633, 
    0.1982632, 0.1982632, 0.1982633, 0.1982634, 0.1982634, 0.1982634, 
    0.1982635, 0.1982634, 0.1982639, 0.1982636, 0.1982631, 0.1982632, 
    0.1982632, 0.1982632, 0.1982634, 0.1982633, 0.1982636, 0.1982635, 
    0.1982636, 0.1982636, 0.1982636, 0.1982635, 0.1982634, 0.1982633, 
    0.1982633, 0.1982632, 0.1982632, 0.1982633, 0.1982634, 0.1982635, 
    0.1982635, 0.1982636, 0.1982633, 0.1982635, 0.1982634, 0.1982635, 
    0.1982633, 0.1982635, 0.1982632, 0.1982633, 0.1982633, 0.1982635, 
    0.1982635, 0.1982635, 0.1982635, 0.1982634, 0.1982634, 0.1982633, 
    0.1982633, 0.1982633, 0.1982632, 0.1982633, 0.1982633, 0.1982634, 
    0.1982635, 0.1982636, 0.1982637, 0.1982638, 0.1982637, 0.1982639, 
    0.1982637, 0.198264, 0.1982635, 0.1982637, 0.1982633, 0.1982634, 
    0.1982634, 0.1982636, 0.1982635, 0.1982636, 0.1982634, 0.1982633, 
    0.1982633, 0.1982632, 0.1982633, 0.1982632, 0.1982633, 0.1982633, 
    0.1982634, 0.1982633, 0.1982636, 0.1982636, 0.1982639, 0.198264, 
    0.1982642, 0.1982643, 0.1982643, 0.1982643,
  0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.601481, 8.601533, 8.601523, 8.601563, 8.601542, 8.601567, 8.601493, 
    8.601534, 8.601508, 8.601487, 8.601641, 8.601565, 8.601724, 8.601675, 
    8.601799, 8.601716, 8.601816, 8.601798, 8.601856, 8.601839, 8.601912, 
    8.601864, 8.601951, 8.601901, 8.601908, 8.601862, 8.601582, 8.601631, 
    8.601579, 8.601585, 8.601583, 8.601542, 8.601521, 8.601479, 8.601486, 
    8.601517, 8.601589, 8.601565, 8.601627, 8.601625, 8.601693, 8.601663, 
    8.601778, 8.601746, 8.60184, 8.601816, 8.601839, 8.601832, 8.601839, 
    8.601804, 8.601819, 8.601789, 8.601668, 8.601704, 8.601599, 8.601534, 
    8.601494, 8.601465, 8.601469, 8.601477, 8.601518, 8.601557, 8.601586, 
    8.601605, 8.601625, 8.601682, 8.601714, 8.601784, 8.601772, 8.601793, 
    8.601814, 8.601848, 8.601843, 8.601857, 8.601793, 8.601835, 8.601766, 
    8.601785, 8.601627, 8.601572, 8.601545, 8.601524, 8.601472, 8.601508, 
    8.601494, 8.601529, 8.60155, 8.60154, 8.601606, 8.601581, 8.601716, 
    8.601657, 8.601811, 8.601774, 8.60182, 8.601797, 8.601836, 8.601801, 
    8.601863, 8.601876, 8.601867, 8.601903, 8.601799, 8.601838, 8.60154, 
    8.601542, 8.601549, 8.601513, 8.601511, 8.601478, 8.601507, 8.60152, 
    8.601552, 8.60157, 8.601588, 8.601627, 8.60167, 8.601732, 8.601777, 
    8.601807, 8.601789, 8.601805, 8.601787, 8.601779, 8.601871, 8.601819, 
    8.601898, 8.601893, 8.601857, 8.601894, 8.601542, 8.601532, 8.601497, 
    8.601524, 8.601475, 8.601502, 8.601518, 8.60158, 8.601595, 8.601607, 
    8.601632, 8.601665, 8.60172, 8.601769, 8.601815, 8.601812, 8.601813, 
    8.601823, 8.601798, 8.601827, 8.601831, 8.601819, 8.601893, 8.601872, 
    8.601893, 8.60188, 8.601536, 8.601553, 8.601543, 8.601561, 8.601548, 
    8.601602, 8.601618, 8.601694, 8.601664, 8.601713, 8.601668, 8.601676, 
    8.601713, 8.601671, 8.601767, 8.601701, 8.601823, 8.601756, 8.601828, 
    8.601815, 8.601836, 8.601854, 8.601878, 8.60192, 8.601911, 8.601947, 
    8.601578, 8.6016, 8.601599, 8.601622, 8.601638, 8.601675, 8.601735, 
    8.601712, 8.601754, 8.601762, 8.6017, 8.601737, 8.601614, 8.601633, 
    8.601623, 8.60158, 8.601717, 8.601645, 8.601778, 8.601739, 8.601851, 
    8.601795, 8.601905, 8.601951, 8.601996, 8.602047, 8.601612, 8.601597, 
    8.601624, 8.60166, 8.601695, 8.601742, 8.601747, 8.601755, 8.601778, 
    8.601796, 8.601757, 8.601801, 8.601637, 8.601724, 8.601591, 8.60163, 
    8.601659, 8.601646, 8.60171, 8.601725, 8.601785, 8.601754, 8.601939, 
    8.601857, 8.602088, 8.602022, 8.601592, 8.601612, 8.601682, 8.601648, 
    8.601745, 8.601768, 8.601788, 8.601811, 8.601815, 8.60183, 8.601806, 
    8.601829, 8.601742, 8.601781, 8.601675, 8.6017, 8.601688, 8.601676, 
    8.601716, 8.601757, 8.601759, 8.601772, 8.601808, 8.601746, 8.601948, 
    8.601821, 8.601634, 8.601672, 8.601679, 8.601664, 8.601766, 8.601728, 
    8.601829, 8.601802, 8.601847, 8.601825, 8.601821, 8.601793, 8.601775, 
    8.60173, 8.601694, 8.601666, 8.601672, 8.601704, 8.60176, 8.601814, 
    8.601803, 8.601843, 8.601738, 8.601782, 8.601765, 8.60181, 8.601712, 
    8.601791, 8.601691, 8.6017, 8.601728, 8.601784, 8.601797, 8.60181, 
    8.601803, 8.601762, 8.601756, 8.601727, 8.601719, 8.601698, 8.601681, 
    8.601696, 8.601713, 8.601763, 8.601806, 8.601854, 8.601867, 8.60192, 
    8.601875, 8.601948, 8.601884, 8.601996, 8.601798, 8.601884, 8.601729, 
    8.601747, 8.601776, 8.601846, 8.60181, 8.601852, 8.601755, 8.601704, 
    8.601692, 8.601667, 8.601692, 8.60169, 8.601714, 8.601707, 8.601764, 
    8.601733, 8.601821, 8.601852, 8.601943, 8.601998, 8.602056, 8.602081, 
    8.602089, 8.602092 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  3.955521e-15, 3.955926e-15, 3.955849e-15, 3.956172e-15, 3.955995e-15, 
    3.956205e-15, 3.955607e-15, 3.955939e-15, 3.955729e-15, 3.955563e-15, 
    3.956788e-15, 3.956187e-15, 3.957447e-15, 3.957057e-15, 3.958049e-15, 
    3.957382e-15, 3.958185e-15, 3.958037e-15, 3.9585e-15, 3.958368e-15, 
    3.958945e-15, 3.958562e-15, 3.959258e-15, 3.958858e-15, 3.958917e-15, 
    3.958548e-15, 3.956315e-15, 3.956711e-15, 3.95629e-15, 3.956347e-15, 
    3.956323e-15, 3.955996e-15, 3.955827e-15, 3.955496e-15, 3.955557e-15, 
    3.955803e-15, 3.956372e-15, 3.956184e-15, 3.956674e-15, 3.956663e-15, 
    3.957204e-15, 3.95696e-15, 3.957877e-15, 3.957618e-15, 3.958374e-15, 
    3.958182e-15, 3.958364e-15, 3.958309e-15, 3.958364e-15, 3.958084e-15, 
    3.958204e-15, 3.957959e-15, 3.957004e-15, 3.957282e-15, 3.95645e-15, 
    3.955939e-15, 3.95562e-15, 3.955388e-15, 3.95542e-15, 3.955481e-15, 
    3.955805e-15, 3.956116e-15, 3.956351e-15, 3.956507e-15, 3.956662e-15, 
    3.957111e-15, 3.957366e-15, 3.957925e-15, 3.957831e-15, 3.957996e-15, 
    3.958164e-15, 3.958436e-15, 3.958392e-15, 3.958511e-15, 3.957996e-15, 
    3.958336e-15, 3.957776e-15, 3.957928e-15, 3.956677e-15, 3.956236e-15, 
    3.956026e-15, 3.955863e-15, 3.955445e-15, 3.955732e-15, 3.955618e-15, 
    3.955895e-15, 3.956067e-15, 3.955983e-15, 3.956511e-15, 3.956305e-15, 
    3.957381e-15, 3.956917e-15, 3.958144e-15, 3.957851e-15, 3.958215e-15, 
    3.958031e-15, 3.958345e-15, 3.958062e-15, 3.958557e-15, 3.958661e-15, 
    3.958589e-15, 3.958876e-15, 3.958046e-15, 3.958361e-15, 3.955979e-15, 
    3.955992e-15, 3.956059e-15, 3.955768e-15, 3.955751e-15, 3.955493e-15, 
    3.955725e-15, 3.955822e-15, 3.956079e-15, 3.956226e-15, 3.956367e-15, 
    3.956679e-15, 3.957023e-15, 3.957513e-15, 3.957869e-15, 3.958108e-15, 
    3.957963e-15, 3.958091e-15, 3.957947e-15, 3.957882e-15, 3.95862e-15, 
    3.958203e-15, 3.958835e-15, 3.9588e-15, 3.958512e-15, 3.958805e-15, 
    3.956003e-15, 3.955924e-15, 3.955642e-15, 3.955863e-15, 3.955465e-15, 
    3.955684e-15, 3.955808e-15, 3.956303e-15, 3.956418e-15, 3.956517e-15, 
    3.956717e-15, 3.956972e-15, 3.957418e-15, 3.957811e-15, 3.958174e-15, 
    3.958149e-15, 3.958157e-15, 3.958236e-15, 3.958038e-15, 3.958268e-15, 
    3.958305e-15, 3.958206e-15, 3.958796e-15, 3.958628e-15, 3.9588e-15, 
    3.958691e-15, 3.95595e-15, 3.956084e-15, 3.956011e-15, 3.956146e-15, 
    3.956049e-15, 3.956474e-15, 3.956602e-15, 3.957208e-15, 3.956966e-15, 
    3.957359e-15, 3.957008e-15, 3.957069e-15, 3.95736e-15, 3.957028e-15, 
    3.957784e-15, 3.957262e-15, 3.958239e-15, 3.957705e-15, 3.958272e-15, 
    3.958173e-15, 3.958339e-15, 3.958485e-15, 3.958675e-15, 3.959015e-15, 
    3.958938e-15, 3.959228e-15, 3.956285e-15, 3.956457e-15, 3.956447e-15, 
    3.956629e-15, 3.956764e-15, 3.957061e-15, 3.957532e-15, 3.957357e-15, 
    3.957685e-15, 3.95775e-15, 3.957253e-15, 3.957553e-15, 3.956575e-15, 
    3.956728e-15, 3.95664e-15, 3.956296e-15, 3.95739e-15, 3.956825e-15, 
    3.957875e-15, 3.957569e-15, 3.958464e-15, 3.958013e-15, 3.958894e-15, 
    3.959258e-15, 3.959625e-15, 3.960027e-15, 3.956556e-15, 3.956439e-15, 
    3.956653e-15, 3.956939e-15, 3.957221e-15, 3.957587e-15, 3.957627e-15, 
    3.957694e-15, 3.957874e-15, 3.958023e-15, 3.95771e-15, 3.958061e-15, 
    3.956753e-15, 3.957442e-15, 3.95639e-15, 3.956699e-15, 3.956925e-15, 
    3.956831e-15, 3.957338e-15, 3.957456e-15, 3.957933e-15, 3.957689e-15, 
    3.959163e-15, 3.958509e-15, 3.960351e-15, 3.959831e-15, 3.956397e-15, 
    3.956558e-15, 3.957111e-15, 3.956848e-15, 3.957614e-15, 3.9578e-15, 
    3.957956e-15, 3.958147e-15, 3.958172e-15, 3.958286e-15, 3.958099e-15, 
    3.958281e-15, 3.957587e-15, 3.957897e-15, 3.957054e-15, 3.957256e-15, 
    3.957165e-15, 3.957061e-15, 3.957381e-15, 3.957714e-15, 3.957729e-15, 
    3.957834e-15, 3.958117e-15, 3.957617e-15, 3.959233e-15, 3.958219e-15, 
    3.956733e-15, 3.957032e-15, 3.957085e-15, 3.956967e-15, 3.957781e-15, 
    3.957485e-15, 3.958284e-15, 3.95807e-15, 3.958424e-15, 3.958247e-15, 
    3.958221e-15, 3.957996e-15, 3.957854e-15, 3.957497e-15, 3.957209e-15, 
    3.956985e-15, 3.957038e-15, 3.957284e-15, 3.957736e-15, 3.958171e-15, 
    3.958074e-15, 3.958397e-15, 3.957558e-15, 3.957905e-15, 3.957768e-15, 
    3.958127e-15, 3.95735e-15, 3.957987e-15, 3.957185e-15, 3.957257e-15, 
    3.957479e-15, 3.957923e-15, 3.958034e-15, 3.958137e-15, 3.958075e-15, 
    3.957749e-15, 3.957699e-15, 3.957476e-15, 3.95741e-15, 3.957242e-15, 
    3.957099e-15, 3.957227e-15, 3.957361e-15, 3.957753e-15, 3.958102e-15, 
    3.958486e-15, 3.958583e-15, 3.959013e-15, 3.958652e-15, 3.959237e-15, 
    3.958723e-15, 3.959622e-15, 3.958035e-15, 3.958724e-15, 3.957492e-15, 
    3.957626e-15, 3.957861e-15, 3.958417e-15, 3.958125e-15, 3.958471e-15, 
    3.957698e-15, 3.957288e-15, 3.957193e-15, 3.956997e-15, 3.957197e-15, 
    3.957181e-15, 3.957372e-15, 3.957311e-15, 3.957766e-15, 3.957522e-15, 
    3.958218e-15, 3.95847e-15, 3.959195e-15, 3.959635e-15, 3.960097e-15, 
    3.960297e-15, 3.960358e-15, 3.960384e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  9.912854, 9.961175, 9.951769, 9.990828, 9.969147, 9.994741, 9.922636, 
    9.963099, 9.937255, 9.917194, 10.0669, 9.992572, 10.14443, 10.09677, 
    10.21673, 10.13701, 10.23285, 10.21441, 10.26993, 10.254, 10.32522, 
    10.27728, 10.36223, 10.31375, 10.32133, 10.2757, 10.0075, 10.05763, 
    10.00453, 10.01167, 10.00846, 9.969597, 9.950049, 9.909162, 9.916575, 
    9.946607, 10.01488, 9.991668, 10.05022, 10.04889, 10.11432, 10.08479, 
    10.19512, 10.16369, 10.25467, 10.23174, 10.25359, 10.24696, 10.25368, 
    10.22007, 10.23446, 10.20491, 10.09031, 10.12392, 10.0239, 9.964057, 
    9.92441, 9.89634, 9.900306, 9.907869, 9.946783, 9.983447, 10.01145, 
    10.0302, 10.0487, 10.10485, 10.13462, 10.20149, 10.18939, 10.20988, 
    10.22946, 10.2624, 10.25698, 10.27151, 10.20933, 10.25063, 10.18251, 
    10.20112, 10.05376, 9.997926, 9.974274, 9.953577, 9.903356, 9.938023, 
    9.924349, 9.956893, 9.97761, 9.96736, 10.03071, 10.00606, 10.13639, 
    10.08012, 10.22718, 10.19187, 10.23565, 10.2133, 10.25162, 10.21713, 
    10.27692, 10.28996, 10.28105, 10.31532, 10.21522, 10.2536, 9.967073, 
    9.968745, 9.976531, 9.942333, 9.940242, 9.90896, 9.936789, 9.948656, 
    9.978809, 9.996676, 10.01368, 10.05112, 10.09303, 10.15181, 10.19416, 
    10.22261, 10.20516, 10.22056, 10.20334, 10.19528, 10.28508, 10.2346, 
    10.31038, 10.30618, 10.27185, 10.30665, 9.969918, 9.960302, 9.926968, 
    9.953049, 9.905557, 9.932127, 9.947426, 10.00658, 10.0196, 10.03168, 
    10.05558, 10.0863, 10.14032, 10.18746, 10.2306, 10.22744, 10.22855, 
    10.23821, 10.21431, 10.24213, 10.24681, 10.23459, 10.30562, 10.2853, 
    10.30609, 10.29286, 9.963427, 9.979612, 9.970864, 9.98732, 9.975727, 
    10.02734, 10.04285, 10.11559, 10.08569, 10.13329, 10.09052, 10.09809, 
    10.13486, 10.09283, 10.18486, 10.12242, 10.23858, 10.17604, 10.24251, 
    10.23042, 10.25044, 10.2684, 10.29101, 10.33281, 10.32312, 10.35813, 
    10.00377, 10.02482, 10.02296, 10.04501, 10.06134, 10.09678, 10.15378, 
    10.13232, 10.17173, 10.17966, 10.11979, 10.15653, 10.03892, 10.05787, 
    10.04658, 10.00543, 10.13727, 10.06948, 10.19486, 10.15798, 10.26584, 
    10.21212, 10.31779, 10.36317, 10.40534, 10.45475, 10.03631, 10.022, 
    10.04763, 10.08318, 10.11621, 10.16023, 10.16474, 10.173, 10.19442, 
    10.21245, 10.17562, 10.21697, 10.06228, 10.14317, 10.01659, 10.05461, 
    10.08108, 10.06946, 10.12987, 10.14414, 10.20226, 10.17219, 10.35196, 
    10.2722, 10.49245, 10.43101, 10.017, 10.03626, 10.10348, 10.07146, 
    10.16317, 10.18582, 10.20425, 10.22785, 10.2304, 10.2444, 10.22146, 
    10.24349, 10.16032, 10.19744, 10.09578, 10.12047, 10.1091, 10.09665, 
    10.13511, 10.1762, 10.17707, 10.19027, 10.22753, 10.16354, 10.3623, 
    10.2393, 10.05729, 10.09451, 10.09982, 10.08539, 10.18355, 10.14792, 
    10.24405, 10.21802, 10.2607, 10.23948, 10.23636, 10.20914, 10.19223, 
    10.14955, 10.11491, 10.08749, 10.09386, 10.124, 10.17871, 10.23063, 
    10.21925, 10.25745, 10.1565, 10.19876, 10.18242, 10.22507, 10.13175, 
    10.21121, 10.11151, 10.12022, 10.14721, 10.20164, 10.21369, 10.22659, 
    10.21863, 10.18011, 10.1738, 10.14656, 10.13905, 10.11832, 10.10119, 
    10.11685, 10.1333, 10.18012, 10.22242, 10.26865, 10.27998, 10.33421, 
    10.29007, 10.36299, 10.30099, 10.40778, 10.21581, 10.29915, 10.14844, 
    10.16461, 10.19391, 10.26128, 10.22487, 10.26745, 10.17355, 10.12504, 
    10.1125, 10.08915, 10.11304, 10.11109, 10.13398, 10.12662, 10.18167, 
    10.15208, 10.23628, 10.26711, 10.35446, 10.40757, 10.46163, 10.48555, 
    10.49284, 10.49589 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  1.67987e-09, 1.66068e-09, 1.664375e-09, 1.64916e-09, 1.657564e-09, 
    1.647653e-09, 1.675942e-09, 1.659928e-09, 1.670114e-09, 1.678124e-09, 
    1.620452e-09, 1.648488e-09, 1.592374e-09, 1.609493e-09, 1.567202e-09, 
    1.595012e-09, 1.561717e-09, 1.567991e-09, 1.549266e-09, 1.554583e-09, 
    1.531133e-09, 1.546825e-09, 1.519266e-09, 1.534851e-09, 1.532391e-09, 
    1.547349e-09, 1.642765e-09, 1.623887e-09, 1.643898e-09, 1.641174e-09, 
    1.642395e-09, 1.657389e-09, 1.665054e-09, 1.681357e-09, 1.678372e-09, 
    1.666411e-09, 1.639952e-09, 1.648834e-09, 1.626642e-09, 1.627136e-09, 
    1.60314e-09, 1.613866e-09, 1.574625e-09, 1.585574e-09, 1.55436e-09, 
    1.562089e-09, 1.554721e-09, 1.556948e-09, 1.554692e-09, 1.56606e-09, 
    1.561168e-09, 1.571249e-09, 1.611846e-09, 1.599688e-09, 1.636531e-09, 
    1.659555e-09, 1.675233e-09, 1.686549e-09, 1.684939e-09, 1.681879e-09, 
    1.666342e-09, 1.652008e-09, 1.641258e-09, 1.634149e-09, 1.627207e-09, 
    1.606565e-09, 1.595862e-09, 1.572429e-09, 1.576606e-09, 1.569545e-09, 
    1.562862e-09, 1.551773e-09, 1.553587e-09, 1.548742e-09, 1.569731e-09, 
    1.555716e-09, 1.578995e-09, 1.572556e-09, 1.625327e-09, 1.646428e-09, 
    1.65557e-09, 1.663663e-09, 1.683704e-09, 1.66981e-09, 1.675258e-09, 
    1.662359e-09, 1.65427e-09, 1.658261e-09, 1.633955e-09, 1.643315e-09, 
    1.595233e-09, 1.615576e-09, 1.563638e-09, 1.575747e-09, 1.560765e-09, 
    1.568373e-09, 1.555384e-09, 1.567064e-09, 1.546947e-09, 1.542637e-09, 
    1.545579e-09, 1.534341e-09, 1.567716e-09, 1.554721e-09, 1.658373e-09, 
    1.65772e-09, 1.654689e-09, 1.668101e-09, 1.66893e-09, 1.681439e-09, 
    1.670299e-09, 1.665602e-09, 1.653805e-09, 1.646908e-09, 1.640409e-09, 
    1.626307e-09, 1.610855e-09, 1.589759e-09, 1.574956e-09, 1.565194e-09, 
    1.571165e-09, 1.565891e-09, 1.571789e-09, 1.57457e-09, 1.544249e-09, 
    1.561123e-09, 1.535947e-09, 1.537318e-09, 1.548627e-09, 1.537163e-09, 
    1.657263e-09, 1.661021e-09, 1.674211e-09, 1.66387e-09, 1.682813e-09, 
    1.672153e-09, 1.666088e-09, 1.643117e-09, 1.63816e-09, 1.63359e-09, 
    1.624645e-09, 1.613314e-09, 1.593831e-09, 1.577277e-09, 1.562475e-09, 
    1.56355e-09, 1.563171e-09, 1.559901e-09, 1.568028e-09, 1.558575e-09, 
    1.557e-09, 1.561125e-09, 1.537502e-09, 1.544175e-09, 1.537347e-09, 
    1.541684e-09, 1.659798e-09, 1.653494e-09, 1.656894e-09, 1.650512e-09, 
    1.655002e-09, 1.63523e-09, 1.629398e-09, 1.602682e-09, 1.613535e-09, 
    1.596334e-09, 1.61177e-09, 1.609012e-09, 1.595778e-09, 1.610928e-09, 
    1.578179e-09, 1.600226e-09, 1.559774e-09, 1.581251e-09, 1.558448e-09, 
    1.562539e-09, 1.555779e-09, 1.549776e-09, 1.542293e-09, 1.52868e-09, 
    1.53181e-09, 1.520569e-09, 1.644189e-09, 1.636182e-09, 1.636885e-09, 
    1.628586e-09, 1.622505e-09, 1.609489e-09, 1.589062e-09, 1.59668e-09, 
    1.582754e-09, 1.579989e-09, 1.601169e-09, 1.588094e-09, 1.63087e-09, 
    1.623795e-09, 1.628e-09, 1.643554e-09, 1.594917e-09, 1.619494e-09, 
    1.574714e-09, 1.58758e-09, 1.550629e-09, 1.568778e-09, 1.533539e-09, 
    1.51897e-09, 1.505521e-09, 1.490109e-09, 1.631848e-09, 1.637249e-09, 
    1.627605e-09, 1.614457e-09, 1.602457e-09, 1.586789e-09, 1.585205e-09, 
    1.582311e-09, 1.574867e-09, 1.568664e-09, 1.581397e-09, 1.567117e-09, 
    1.622162e-09, 1.592821e-09, 1.6393e-09, 1.625006e-09, 1.615226e-09, 
    1.619502e-09, 1.597556e-09, 1.592473e-09, 1.572164e-09, 1.582595e-09, 
    1.522538e-09, 1.548513e-09, 1.478594e-09, 1.497466e-09, 1.639145e-09, 
    1.631867e-09, 1.607057e-09, 1.618762e-09, 1.585755e-09, 1.577845e-09, 
    1.571476e-09, 1.56341e-09, 1.562545e-09, 1.557813e-09, 1.565583e-09, 
    1.558118e-09, 1.586756e-09, 1.573824e-09, 1.609854e-09, 1.600926e-09, 
    1.60502e-09, 1.609536e-09, 1.595683e-09, 1.581195e-09, 1.58089e-09, 
    1.576304e-09, 1.563527e-09, 1.585624e-09, 1.519249e-09, 1.559537e-09, 
    1.624008e-09, 1.610316e-09, 1.608382e-09, 1.613643e-09, 1.578634e-09, 
    1.591134e-09, 1.557928e-09, 1.566759e-09, 1.552344e-09, 1.559472e-09, 
    1.560527e-09, 1.569796e-09, 1.575625e-09, 1.590556e-09, 1.602925e-09, 
    1.612878e-09, 1.610552e-09, 1.599659e-09, 1.580318e-09, 1.562466e-09, 
    1.566341e-09, 1.55343e-09, 1.588101e-09, 1.573367e-09, 1.579027e-09, 
    1.564357e-09, 1.596883e-09, 1.569094e-09, 1.604152e-09, 1.601013e-09, 
    1.591384e-09, 1.572377e-09, 1.568238e-09, 1.563841e-09, 1.566551e-09, 
    1.579833e-09, 1.582033e-09, 1.591617e-09, 1.594284e-09, 1.601695e-09, 
    1.607886e-09, 1.602228e-09, 1.59633e-09, 1.579828e-09, 1.565259e-09, 
    1.549691e-09, 1.54593e-09, 1.52823e-09, 1.542605e-09, 1.51903e-09, 
    1.539023e-09, 1.504754e-09, 1.567516e-09, 1.539621e-09, 1.590949e-09, 
    1.585249e-09, 1.575044e-09, 1.552152e-09, 1.564425e-09, 1.550092e-09, 
    1.582119e-09, 1.599285e-09, 1.603792e-09, 1.612269e-09, 1.603599e-09, 
    1.604301e-09, 1.596088e-09, 1.598717e-09, 1.579287e-09, 1.589662e-09, 
    1.560553e-09, 1.550205e-09, 1.521739e-09, 1.504817e-09, 1.487989e-09, 
    1.480683e-09, 1.478474e-09, 1.477552e-09 ;

 W_SCALAR =
  0.6251647, 0.6268236, 0.6265013, 0.6278382, 0.6270967, 0.6279719, 
    0.6255011, 0.6268895, 0.6260033, 0.625314, 0.6304291, 0.6278978, 
    0.6330526, 0.6314422, 0.6354835, 0.6328022, 0.6360235, 0.6354061, 
    0.6372628, 0.6367311, 0.6391034, 0.6375081, 0.6403309, 0.6387225, 
    0.6389743, 0.6374555, 0.6284074, 0.6301143, 0.6283063, 0.6285498, 
    0.6284405, 0.627112, 0.6264422, 0.6250377, 0.6252927, 0.6263242, 
    0.6286593, 0.627867, 0.6298626, 0.6298175, 0.6320359, 0.6310362, 
    0.6347587, 0.6337017, 0.6367534, 0.6359866, 0.6367174, 0.6364958, 
    0.6367203, 0.6355956, 0.6360776, 0.6350874, 0.6312234, 0.6323603, 
    0.6289667, 0.6269222, 0.6255621, 0.6245962, 0.6247327, 0.6249931, 
    0.6263303, 0.627586, 0.6285422, 0.6291815, 0.6298111, 0.6317154, 
    0.6327217, 0.6349724, 0.6345664, 0.635254, 0.6359103, 0.6370117, 
    0.6368305, 0.6373155, 0.6352357, 0.6366184, 0.634335, 0.63496, 0.6299828, 
    0.6280808, 0.627272, 0.6265633, 0.6248378, 0.6260296, 0.6255599, 
    0.626677, 0.6273863, 0.6270355, 0.629199, 0.6283583, 0.6327813, 0.630878, 
    0.6358338, 0.6346497, 0.6361175, 0.6353686, 0.6366514, 0.635497, 
    0.6374959, 0.6379308, 0.6376337, 0.6387746, 0.635433, 0.6367174, 
    0.6270257, 0.6270829, 0.6273494, 0.6261775, 0.6261058, 0.6250307, 
    0.6259873, 0.6263945, 0.6274274, 0.628038, 0.6286183, 0.6298931, 
    0.6313155, 0.6333016, 0.6347265, 0.6356807, 0.6350957, 0.6356122, 
    0.6350347, 0.634764, 0.637768, 0.6360821, 0.6386105, 0.6384708, 
    0.6373271, 0.6384865, 0.6271231, 0.6267938, 0.6256499, 0.6265452, 
    0.6249136, 0.6258272, 0.6263523, 0.6283761, 0.6288201, 0.6292319, 
    0.6300448, 0.6310873, 0.6329141, 0.6345014, 0.6359485, 0.6358425, 
    0.6358798, 0.6362029, 0.6354025, 0.6363343, 0.6364907, 0.6360819, 
    0.6384521, 0.6377754, 0.6384678, 0.6380273, 0.6269008, 0.6274548, 
    0.6271555, 0.6277183, 0.6273219, 0.6290841, 0.6296119, 0.6320789, 
    0.6310669, 0.632677, 0.6312305, 0.6314869, 0.6327297, 0.6313086, 
    0.634414, 0.6323097, 0.6362155, 0.6341174, 0.6363469, 0.6359422, 
    0.6366121, 0.6372117, 0.6379656, 0.6393555, 0.6390338, 0.6401951, 
    0.6282803, 0.6289981, 0.6289348, 0.6296856, 0.6302406, 0.6314425, 
    0.633368, 0.6326442, 0.6339725, 0.634239, 0.6322209, 0.6334605, 
    0.6294782, 0.6301226, 0.6297389, 0.628337, 0.6328112, 0.630517, 0.63475, 
    0.6335096, 0.6371263, 0.6353291, 0.6388566, 0.6403618, 0.6417761, 
    0.6434274, 0.6293896, 0.628902, 0.6297748, 0.6309816, 0.6320999, 
    0.6335853, 0.6337371, 0.6340152, 0.6347351, 0.6353402, 0.6341032, 
    0.6354917, 0.6302722, 0.6330101, 0.6287178, 0.6300119, 0.6309104, 
    0.6305162, 0.6325614, 0.6330431, 0.6349983, 0.6339878, 0.6399906, 
    0.6373385, 0.6446828, 0.642635, 0.6287317, 0.6293879, 0.6316692, 
    0.6305842, 0.6336843, 0.6344463, 0.6350653, 0.6358563, 0.6359416, 
    0.6364099, 0.6356423, 0.6363796, 0.6335885, 0.6348366, 0.6314085, 
    0.6322438, 0.6318595, 0.6314381, 0.6327385, 0.6341228, 0.6341521, 
    0.6345957, 0.6358451, 0.6336969, 0.6403329, 0.6362392, 0.6301031, 
    0.6313656, 0.6315456, 0.6310568, 0.63437, 0.6331705, 0.6363985, 
    0.6355269, 0.6369547, 0.6362454, 0.6361411, 0.6352293, 0.6346615, 
    0.6332256, 0.632056, 0.6311277, 0.6313435, 0.6323631, 0.6342074, 
    0.6359494, 0.635568, 0.6368462, 0.6334598, 0.634881, 0.634332, 0.635763, 
    0.632625, 0.6352983, 0.6319409, 0.6322356, 0.6331467, 0.6349775, 
    0.6353819, 0.6358139, 0.6355473, 0.6342541, 0.634042, 0.6331245, 
    0.6328712, 0.6321714, 0.6315919, 0.6321214, 0.6326774, 0.6342546, 
    0.6356743, 0.6372203, 0.6375982, 0.639402, 0.6379341, 0.6403556, 
    0.6382976, 0.6418577, 0.6354527, 0.6382366, 0.6331881, 0.6337329, 
    0.634718, 0.6369739, 0.6357563, 0.6371801, 0.6340337, 0.6323984, 
    0.6319746, 0.6311842, 0.6319927, 0.631927, 0.6327003, 0.6324518, 
    0.6343069, 0.6333107, 0.6361384, 0.6371688, 0.6400735, 0.6418509, 
    0.643657, 0.6444536, 0.6446959, 0.6447972,
  0.546157, 0.5482014, 0.5478041, 0.5494519, 0.5485379, 0.5496167, 0.5465716, 
    0.5482826, 0.5471904, 0.546341, 0.5526459, 0.5495253, 0.555881, 
    0.5538949, 0.5588794, 0.5555722, 0.5595455, 0.5587839, 0.5610747, 
    0.5604187, 0.563346, 0.5613773, 0.5648611, 0.5628759, 0.5631867, 
    0.5613124, 0.5501536, 0.5522578, 0.5500289, 0.550329, 0.5501943, 
    0.5485569, 0.5477313, 0.5460005, 0.5463148, 0.5475859, 0.550464, 
    0.5494874, 0.5519474, 0.5518919, 0.554627, 0.5533943, 0.5579852, 
    0.5566816, 0.5604461, 0.5595002, 0.5604017, 0.5601283, 0.5604053, 
    0.5590177, 0.5596123, 0.5583908, 0.5536253, 0.5550272, 0.550843, 
    0.5483229, 0.5466467, 0.5454565, 0.5456248, 0.5459456, 0.5475933, 
    0.549141, 0.5503197, 0.5511078, 0.5518839, 0.5542318, 0.5554729, 
    0.5582489, 0.557748, 0.5585963, 0.559406, 0.5607648, 0.5605412, 
    0.5611397, 0.5585737, 0.5602796, 0.5574627, 0.5582336, 0.5520956, 
    0.5497509, 0.548754, 0.5478805, 0.5457542, 0.5472229, 0.546644, 
    0.5480206, 0.5488949, 0.5484625, 0.5511293, 0.550093, 0.5555463, 
    0.5531994, 0.5593116, 0.5578508, 0.5596615, 0.5587378, 0.5603203, 
    0.5588961, 0.5613623, 0.561899, 0.5615323, 0.5629402, 0.5588171, 
    0.5604017, 0.5484505, 0.548521, 0.5488495, 0.5474051, 0.5473167, 
    0.5459919, 0.5471707, 0.5476725, 0.5489455, 0.5496982, 0.5504134, 
    0.551985, 0.5537388, 0.556188, 0.5579455, 0.5591227, 0.5584009, 
    0.5590382, 0.5583258, 0.5579918, 0.561698, 0.5596179, 0.5627378, 
    0.5625653, 0.5611539, 0.5625847, 0.5485705, 0.5481646, 0.546755, 
    0.5478582, 0.5458476, 0.5469734, 0.5476205, 0.5501148, 0.5506622, 
    0.5511699, 0.5521721, 0.5534574, 0.5557102, 0.5576679, 0.5594531, 
    0.5593223, 0.5593683, 0.559767, 0.5587795, 0.5599291, 0.560122, 
    0.5596176, 0.5625422, 0.5617071, 0.5625616, 0.5620179, 0.5482965, 
    0.5489793, 0.5486104, 0.5493042, 0.5488155, 0.5509876, 0.5516384, 
    0.5546801, 0.5534322, 0.5554177, 0.5536339, 0.5539501, 0.5554827, 
    0.5537303, 0.5575601, 0.5549648, 0.5597825, 0.5571942, 0.5599446, 
    0.5594453, 0.5602717, 0.5610116, 0.5619419, 0.5636572, 0.5632601, 
    0.5646935, 0.5499968, 0.5508817, 0.5508036, 0.5517291, 0.5524134, 
    0.5538954, 0.5562699, 0.5553773, 0.5570155, 0.5573443, 0.5548552, 
    0.556384, 0.5514736, 0.5522679, 0.5517949, 0.5500666, 0.5555832, 
    0.5527542, 0.5579746, 0.5564446, 0.5609062, 0.5586889, 0.5630415, 
    0.5648993, 0.5666452, 0.568684, 0.5513642, 0.5507632, 0.5518392, 
    0.553327, 0.554706, 0.556538, 0.5567252, 0.5570682, 0.5579562, 0.5587025, 
    0.5571768, 0.5588896, 0.5524524, 0.5558285, 0.5505361, 0.5521315, 
    0.5532393, 0.5527533, 0.5552752, 0.5558692, 0.5582808, 0.5570344, 
    0.5644411, 0.5611681, 0.5702342, 0.5677056, 0.5505532, 0.5513622, 
    0.554175, 0.5528371, 0.5566601, 0.5576, 0.5583635, 0.5593393, 0.5594445, 
    0.5600224, 0.5590754, 0.5599849, 0.5565419, 0.5580813, 0.5538535, 
    0.5548835, 0.5544097, 0.5538899, 0.5554936, 0.5572008, 0.5572371, 
    0.5577842, 0.5593255, 0.5566756, 0.5648635, 0.5598118, 0.5522438, 
    0.5538005, 0.5540225, 0.5534198, 0.5575058, 0.5560263, 0.5600083, 
    0.558933, 0.5606945, 0.5598193, 0.5596906, 0.5585659, 0.5578654, 
    0.5560943, 0.5546519, 0.5535071, 0.5537734, 0.5550306, 0.5573052, 
    0.5594542, 0.5589837, 0.5605606, 0.5563832, 0.5581362, 0.5574589, 
    0.5592243, 0.5553536, 0.558651, 0.5545099, 0.5548733, 0.555997, 
    0.5582552, 0.5587541, 0.559287, 0.5589581, 0.5573629, 0.5571012, 
    0.5559696, 0.5556571, 0.5547942, 0.5540795, 0.5547326, 0.5554181, 
    0.5573635, 0.5591148, 0.5610222, 0.5614886, 0.5637145, 0.5619031, 
    0.5648916, 0.5623516, 0.5667459, 0.5588415, 0.5622764, 0.556048, 0.55672, 
    0.5579351, 0.5607182, 0.559216, 0.5609726, 0.557091, 0.5550741, 
    0.5545516, 0.5535768, 0.5545738, 0.5544928, 0.5554464, 0.55514, 0.557428, 
    0.5561993, 0.5596874, 0.5609587, 0.5645434, 0.5667375, 0.5689675, 
    0.5699512, 0.5702505, 0.5703756,
  0.5139313, 0.5161815, 0.5157441, 0.5175582, 0.516552, 0.5177397, 0.5143875, 
    0.5162709, 0.5150687, 0.5141338, 0.5210757, 0.5176391, 0.5246401, 
    0.5224517, 0.5279453, 0.5242998, 0.5286797, 0.52784, 0.5303661, 
    0.5296426, 0.5328715, 0.5306999, 0.5345433, 0.5323529, 0.5326958, 
    0.5306283, 0.5183308, 0.5206482, 0.5181935, 0.5185241, 0.5183757, 
    0.5165728, 0.515664, 0.5137591, 0.514105, 0.515504, 0.5186727, 0.5175973, 
    0.5203063, 0.5202452, 0.5232583, 0.5219002, 0.5269595, 0.5255224, 
    0.5296728, 0.5286297, 0.5296239, 0.5293224, 0.5296278, 0.5280977, 
    0.5287534, 0.5274066, 0.5221546, 0.5236993, 0.51909, 0.5163153, 
    0.5144702, 0.5131604, 0.5133456, 0.5136987, 0.5155122, 0.517216, 
    0.5185137, 0.5193816, 0.5202364, 0.5228229, 0.5241903, 0.5272501, 
    0.5266979, 0.5276331, 0.5285259, 0.5300243, 0.5297777, 0.5304378, 
    0.5276083, 0.5294892, 0.5263835, 0.5272333, 0.5204695, 0.5178874, 
    0.5167899, 0.5158283, 0.513488, 0.5151044, 0.5144673, 0.5159825, 
    0.516945, 0.516469, 0.5194053, 0.5182641, 0.5242713, 0.5216854, 
    0.5284218, 0.5268112, 0.5288076, 0.5277891, 0.529534, 0.5279636, 
    0.5306833, 0.5312753, 0.5308708, 0.5324239, 0.5278766, 0.5296239, 
    0.5164557, 0.5165333, 0.5168949, 0.515305, 0.5152077, 0.5137497, 
    0.515047, 0.5155994, 0.5170007, 0.5178295, 0.518617, 0.5203478, 
    0.5222796, 0.5249785, 0.5269157, 0.5282135, 0.5274177, 0.5281203, 
    0.5273349, 0.5269667, 0.5310535, 0.5287595, 0.5322006, 0.5320103, 
    0.5304535, 0.5320317, 0.5165879, 0.516141, 0.5145894, 0.5158038, 
    0.5135908, 0.5148298, 0.515542, 0.5182882, 0.518891, 0.5194501, 
    0.5205538, 0.5219697, 0.5244519, 0.5266096, 0.5285777, 0.5284336, 
    0.5284843, 0.5289239, 0.5278351, 0.5291026, 0.5293154, 0.5287592, 
    0.5319847, 0.5310636, 0.5320062, 0.5314065, 0.5162863, 0.517038, 
    0.5166318, 0.5173956, 0.5168576, 0.5192493, 0.5199659, 0.5233168, 
    0.5219419, 0.5241295, 0.5221641, 0.5225125, 0.5242012, 0.5222703, 
    0.5264909, 0.5236305, 0.528941, 0.5260875, 0.5291197, 0.5285692, 
    0.5294805, 0.5302965, 0.5313225, 0.5332149, 0.5327768, 0.5343584, 
    0.5181582, 0.5191326, 0.5190467, 0.520066, 0.5208196, 0.5224522, 
    0.5250688, 0.524085, 0.5258905, 0.5262529, 0.5235097, 0.5251945, 
    0.5197845, 0.5206594, 0.5201384, 0.5182351, 0.524312, 0.5211951, 
    0.5269477, 0.5252612, 0.5301802, 0.5277352, 0.5325356, 0.5345855, 
    0.5365125, 0.5387634, 0.5196641, 0.5190022, 0.5201871, 0.521826, 
    0.5233454, 0.5253642, 0.5255706, 0.5259486, 0.5269275, 0.5277503, 
    0.5260683, 0.5279564, 0.5208626, 0.5245823, 0.518752, 0.5205091, 
    0.5217294, 0.521194, 0.5239726, 0.5246271, 0.5272853, 0.5259114, 
    0.5340798, 0.5304691, 0.5404754, 0.5376831, 0.5187709, 0.5196617, 
    0.5227602, 0.5212864, 0.5254988, 0.5265348, 0.5273765, 0.5284523, 
    0.5285684, 0.5292056, 0.5281613, 0.5291643, 0.5253685, 0.5270654, 
    0.522406, 0.5235409, 0.5230188, 0.5224462, 0.5242132, 0.5260948, 
    0.5261347, 0.5267379, 0.5284371, 0.5255159, 0.534546, 0.5289733, 
    0.5206329, 0.5223477, 0.5225922, 0.5219282, 0.5264309, 0.5248003, 
    0.52919, 0.5280043, 0.5299467, 0.5289817, 0.5288397, 0.5275996, 
    0.5268273, 0.5248752, 0.5232857, 0.5220245, 0.5223178, 0.523703, 
    0.5262098, 0.528579, 0.5280603, 0.5297992, 0.5251936, 0.5271259, 
    0.5263793, 0.5283255, 0.5240589, 0.5276934, 0.5231293, 0.5235297, 
    0.5247679, 0.5272571, 0.5278071, 0.5283946, 0.5280321, 0.5262734, 
    0.525985, 0.5247378, 0.5243934, 0.5234425, 0.5226551, 0.5233746, 0.52413, 
    0.526274, 0.5282048, 0.5303082, 0.5308225, 0.5332782, 0.5312797, 
    0.5345771, 0.5317745, 0.5366237, 0.5279034, 0.5316915, 0.5248242, 
    0.5255648, 0.5269042, 0.5299729, 0.5283164, 0.5302535, 0.5259737, 
    0.5237509, 0.5231752, 0.5221012, 0.5231997, 0.5231104, 0.5241612, 
    0.5238235, 0.5263452, 0.5249909, 0.5288362, 0.5302381, 0.5341928, 
    0.5366143, 0.5390764, 0.5401628, 0.5404934, 0.5406315,
  0.5071235, 0.5095142, 0.5090494, 0.5109773, 0.5099078, 0.5111702, 
    0.5076081, 0.5096092, 0.5083317, 0.5073386, 0.5147178, 0.5110633, 
    0.5185111, 0.5161818, 0.5220314, 0.5181488, 0.522814, 0.5219192, 
    0.5246115, 0.5238402, 0.5272833, 0.5249674, 0.529067, 0.5267302, 
    0.5270959, 0.524891, 0.5117986, 0.514263, 0.5116526, 0.5120041, 
    0.5118464, 0.50993, 0.5089643, 0.5069406, 0.507308, 0.5087942, 0.5121621, 
    0.5110189, 0.5138994, 0.5138344, 0.5170403, 0.515595, 0.5209812, 
    0.5194507, 0.5238724, 0.5227607, 0.5238203, 0.523499, 0.5238245, 
    0.5221938, 0.5228925, 0.5214575, 0.5158657, 0.5175096, 0.5126059, 
    0.5096563, 0.507696, 0.5063048, 0.5065015, 0.5068765, 0.5088029, 
    0.5106135, 0.5119932, 0.5129159, 0.513825, 0.5165768, 0.5180323, 
    0.5212908, 0.5207026, 0.5216988, 0.5226501, 0.5242472, 0.5239843, 
    0.5246879, 0.5216724, 0.5236768, 0.5203676, 0.5212729, 0.514073, 
    0.5113273, 0.5101607, 0.5091388, 0.5066527, 0.5083697, 0.5076929, 
    0.5093027, 0.5103256, 0.5098196, 0.5129412, 0.5117278, 0.5181186, 
    0.5153664, 0.5225391, 0.5208233, 0.5229503, 0.521865, 0.5237246, 
    0.522051, 0.5249497, 0.5255808, 0.5251496, 0.5268058, 0.5219582, 
    0.5238203, 0.5098055, 0.5098881, 0.5102723, 0.5085828, 0.5084794, 
    0.5069306, 0.5083087, 0.5088955, 0.5103848, 0.5112657, 0.512103, 
    0.5139435, 0.5159987, 0.5188715, 0.5209346, 0.5223172, 0.5214694, 
    0.5222179, 0.5213811, 0.5209889, 0.5253444, 0.5228991, 0.5265676, 
    0.5263647, 0.5247047, 0.5263875, 0.5099459, 0.5094711, 0.5078226, 
    0.5091127, 0.5067619, 0.508078, 0.5088347, 0.5117533, 0.5123942, 
    0.5129887, 0.5141626, 0.5156689, 0.5183108, 0.5206085, 0.5227054, 
    0.5225518, 0.5226058, 0.5230743, 0.521914, 0.5232648, 0.5234915, 
    0.5228987, 0.5263375, 0.5253552, 0.5263603, 0.5257208, 0.5096254, 
    0.5104244, 0.5099927, 0.5108045, 0.5102326, 0.5127752, 0.5135373, 
    0.5171025, 0.5156393, 0.5179676, 0.5158758, 0.5162466, 0.5180439, 
    0.5159888, 0.520482, 0.5174364, 0.5230925, 0.5200525, 0.5232829, 
    0.5226963, 0.5236675, 0.5245373, 0.5256313, 0.5276496, 0.5271823, 
    0.5288697, 0.5116151, 0.5126511, 0.5125598, 0.5136437, 0.5144454, 
    0.5161823, 0.5189676, 0.5179203, 0.5198427, 0.5202286, 0.5173079, 
    0.5191014, 0.5133443, 0.514275, 0.5137208, 0.5116969, 0.5181618, 
    0.5148448, 0.5209687, 0.5191725, 0.5244133, 0.5218076, 0.526925, 
    0.529112, 0.5311689, 0.5335729, 0.5132164, 0.5125125, 0.5137726, 
    0.515516, 0.5171329, 0.5192821, 0.5195019, 0.5199045, 0.5209471, 
    0.5218236, 0.520032, 0.5220433, 0.5144911, 0.5184496, 0.5122465, 
    0.5141151, 0.5154132, 0.5148436, 0.5178005, 0.5184973, 0.5213283, 
    0.5198649, 0.5285724, 0.5247213, 0.5354021, 0.532419, 0.5122666, 
    0.5132139, 0.5165101, 0.5149419, 0.5194255, 0.5205288, 0.5214254, 
    0.5225717, 0.5226954, 0.5233744, 0.5222617, 0.5233305, 0.5192867, 
    0.521094, 0.5161332, 0.517341, 0.5167854, 0.5161759, 0.5180567, 
    0.5200602, 0.5201027, 0.5207451, 0.5225555, 0.5194436, 0.5290699, 
    0.5231269, 0.5142467, 0.5160711, 0.5163314, 0.5156248, 0.5204182, 
    0.5186818, 0.5233579, 0.5220943, 0.5241644, 0.5231358, 0.5229845, 
    0.5216631, 0.5208404, 0.5187615, 0.5170694, 0.5157272, 0.5160393, 
    0.5175136, 0.5201827, 0.5227067, 0.5221539, 0.5240071, 0.5191005, 
    0.5211585, 0.5203632, 0.5224366, 0.5178925, 0.521763, 0.5169029, 
    0.5173291, 0.5186473, 0.5212982, 0.5218842, 0.5225103, 0.5221239, 
    0.5202504, 0.5199433, 0.5186152, 0.5182486, 0.5172363, 0.5163983, 
    0.5171641, 0.5179682, 0.5202511, 0.5223079, 0.5245497, 0.5250981, 
    0.5277171, 0.5255856, 0.529103, 0.5261132, 0.5312877, 0.5219868, 
    0.5260248, 0.5187072, 0.5194958, 0.5209222, 0.5241923, 0.5224268, 
    0.5244914, 0.5199313, 0.5175645, 0.5169517, 0.5158089, 0.5169779, 
    0.5168828, 0.5180013, 0.5176418, 0.5203269, 0.5188847, 0.5229808, 
    0.524475, 0.528693, 0.5312777, 0.5339073, 0.5350681, 0.5354213, 0.535569,
  0.5311409, 0.5336103, 0.53313, 0.5351228, 0.5340171, 0.5353222, 0.5316414, 
    0.5337085, 0.5323887, 0.531363, 0.5389929, 0.5352116, 0.5429236, 
    0.5405093, 0.5465766, 0.5425479, 0.5473894, 0.54646, 0.5492572, 
    0.5484556, 0.552036, 0.5496271, 0.553893, 0.5514605, 0.551841, 0.5495477, 
    0.5359721, 0.5385221, 0.5358211, 0.5361846, 0.5360214, 0.53404, 
    0.5330421, 0.5309521, 0.5313314, 0.5328664, 0.536348, 0.5351657, 
    0.5381457, 0.5380784, 0.5413988, 0.5399013, 0.5454862, 0.543898, 
    0.548489, 0.547334, 0.5484348, 0.5481009, 0.5484391, 0.5467452, 
    0.5474709, 0.5459806, 0.5401818, 0.5418853, 0.5368071, 0.5337572, 
    0.531732, 0.5302957, 0.5304988, 0.5308859, 0.5328754, 0.5347466, 
    0.5361732, 0.5371279, 0.5380687, 0.5409185, 0.5424271, 0.5458076, 
    0.5451971, 0.5462312, 0.5472191, 0.5488785, 0.5486053, 0.5493366, 
    0.5462037, 0.5482857, 0.5448494, 0.545789, 0.5383254, 0.5354846, 
    0.5342785, 0.5332224, 0.5306549, 0.5324278, 0.5317289, 0.5333918, 
    0.5344489, 0.533926, 0.537154, 0.5358987, 0.5425165, 0.5396647, 
    0.5471038, 0.5453224, 0.5475309, 0.5464038, 0.5483354, 0.5465969, 
    0.5496088, 0.550265, 0.5498165, 0.5515392, 0.5465006, 0.5484349, 
    0.5339114, 0.5339966, 0.5343939, 0.532648, 0.5325412, 0.5309417, 
    0.5323648, 0.5329711, 0.5345101, 0.5354209, 0.5362868, 0.5381913, 
    0.5403196, 0.5432973, 0.5454378, 0.5468734, 0.545993, 0.5467702, 
    0.5459014, 0.5454942, 0.5500191, 0.5474778, 0.5512914, 0.5510802, 
    0.5493541, 0.5511041, 0.5340565, 0.5335658, 0.5318628, 0.5331955, 
    0.5307676, 0.5321265, 0.5329082, 0.5359252, 0.5365881, 0.5372033, 
    0.5384182, 0.539978, 0.5427158, 0.5450994, 0.5472765, 0.5471169, 
    0.5471731, 0.5476598, 0.5464547, 0.5478576, 0.5480932, 0.5474774, 
    0.551052, 0.5500304, 0.5510758, 0.5504105, 0.5337253, 0.534551, 
    0.5341048, 0.534944, 0.5343528, 0.5369823, 0.537771, 0.5414633, 
    0.5399473, 0.5423601, 0.5401922, 0.5405763, 0.5424392, 0.5403093, 
    0.5449681, 0.5418093, 0.5476786, 0.5445224, 0.5478765, 0.5472671, 
    0.5482761, 0.5491801, 0.5503175, 0.5524173, 0.5519309, 0.5536875, 
    0.5357823, 0.536854, 0.5367594, 0.5378811, 0.5387109, 0.5405098, 
    0.5433969, 0.542311, 0.5443047, 0.5447052, 0.5416761, 0.5435358, 
    0.5375712, 0.5385344, 0.5379608, 0.5358669, 0.5425614, 0.5391244, 
    0.5454732, 0.5436096, 0.5490512, 0.5463442, 0.5516632, 0.5539398, 
    0.5560829, 0.5585899, 0.5374388, 0.5367104, 0.5380145, 0.5398196, 
    0.5414948, 0.5437232, 0.5439512, 0.5443689, 0.5454508, 0.5463608, 
    0.5445011, 0.546589, 0.5387582, 0.5428598, 0.5364353, 0.538369, 
    0.5397131, 0.5391232, 0.5421868, 0.5429093, 0.5458465, 0.5443277, 
    0.553378, 0.5493713, 0.5604994, 0.5573863, 0.536456, 0.5374362, 
    0.5408494, 0.539225, 0.5438719, 0.5450167, 0.5459474, 0.5471377, 
    0.5472661, 0.5479715, 0.5468157, 0.5479258, 0.5437279, 0.5456033, 
    0.5404589, 0.5417105, 0.5411347, 0.5405031, 0.5424524, 0.5445305, 
    0.5445746, 0.5452412, 0.5471208, 0.5438908, 0.553896, 0.5477144, 
    0.5385052, 0.5403947, 0.5406643, 0.5399323, 0.5449019, 0.5431005, 
    0.5479543, 0.5466419, 0.5487925, 0.5477237, 0.5475665, 0.5461941, 
    0.5453401, 0.5431831, 0.541429, 0.5400383, 0.5403616, 0.5418894, 
    0.5446575, 0.5472779, 0.5467038, 0.548629, 0.5435348, 0.5456702, 
    0.5448449, 0.5469973, 0.5422822, 0.5462978, 0.5412565, 0.5416982, 
    0.5430648, 0.5458153, 0.5464237, 0.5470738, 0.5466726, 0.5447278, 
    0.5444091, 0.5430315, 0.5426514, 0.541602, 0.5407336, 0.5415271, 
    0.5423606, 0.5447285, 0.5468637, 0.549193, 0.5497631, 0.5524875, 0.55027, 
    0.5539305, 0.5508187, 0.5562066, 0.5465303, 0.5507267, 0.5431269, 
    0.5439448, 0.5454251, 0.5488215, 0.5469872, 0.5491323, 0.5443966, 
    0.5419422, 0.5413071, 0.5401229, 0.5413342, 0.5412356, 0.5423949, 
    0.5420223, 0.5448071, 0.543311, 0.5475626, 0.5491154, 0.5535035, 
    0.5561963, 0.5589389, 0.5601506, 0.5605194, 0.5606736,
  0.5352592, 0.5381025, 0.5375492, 0.5398464, 0.5385715, 0.5400766, 0.535835, 
    0.5382156, 0.5366953, 0.5355148, 0.5443176, 0.539949, 0.5488714, 
    0.5460728, 0.5531155, 0.5484356, 0.5540615, 0.55298, 0.5562374, 
    0.5553033, 0.5594807, 0.5566688, 0.5616519, 0.5588084, 0.5592529, 
    0.5565763, 0.5408266, 0.5437729, 0.5406523, 0.541072, 0.5408835, 
    0.5385979, 0.5374479, 0.535042, 0.5354784, 0.5372455, 0.5412607, 
    0.539896, 0.5433377, 0.5432599, 0.5471033, 0.5453688, 0.5518475, 
    0.5500024, 0.5553422, 0.553997, 0.555279, 0.5548901, 0.5552841, 
    0.5533118, 0.5541564, 0.5524224, 0.5456935, 0.5476671, 0.5417908, 
    0.5382718, 0.5359394, 0.5342872, 0.5345206, 0.5349658, 0.5372558, 
    0.5394126, 0.5410588, 0.5421614, 0.5432487, 0.5465468, 0.5482955, 
    0.5522211, 0.5515115, 0.5527138, 0.5538632, 0.5557961, 0.5554777, 
    0.5563301, 0.5526819, 0.5551053, 0.5511075, 0.5521995, 0.5435455, 
    0.540264, 0.5388727, 0.5376556, 0.5347002, 0.5367404, 0.5359358, 
    0.5378507, 0.5390692, 0.5384664, 0.5421916, 0.540742, 0.5483992, 
    0.5450948, 0.5537291, 0.5516571, 0.5542263, 0.5529145, 0.5551632, 
    0.5531392, 0.5566474, 0.5574129, 0.5568898, 0.5589004, 0.5530271, 
    0.5552791, 0.5384496, 0.5385479, 0.5390058, 0.536994, 0.536871, 
    0.5350301, 0.5366679, 0.537366, 0.5391399, 0.5401905, 0.54119, 0.5433905, 
    0.5458531, 0.5493051, 0.5517913, 0.5534609, 0.5524367, 0.5533409, 
    0.5523303, 0.5518568, 0.5571261, 0.5541644, 0.5586109, 0.5583644, 
    0.5563504, 0.5583922, 0.5386169, 0.5380513, 0.5360899, 0.5376246, 
    0.5348298, 0.5363935, 0.5372936, 0.5407725, 0.5415379, 0.5422484, 
    0.5436527, 0.5454575, 0.5486304, 0.551398, 0.5539301, 0.5537444, 
    0.5538098, 0.5543762, 0.5529737, 0.5546067, 0.554881, 0.5541639, 
    0.5583314, 0.5571392, 0.5583591, 0.5575827, 0.5382351, 0.539187, 
    0.5386726, 0.5396402, 0.5389585, 0.5419931, 0.5429045, 0.547178, 
    0.545422, 0.5482177, 0.5457056, 0.5461504, 0.5483094, 0.5458412, 
    0.5512454, 0.5475792, 0.5543983, 0.5507275, 0.5546287, 0.5539191, 
    0.5550941, 0.5561476, 0.5574741, 0.5599262, 0.5593579, 0.5614115, 
    0.5406075, 0.5418449, 0.5417357, 0.5430318, 0.5439913, 0.5460734, 
    0.5494207, 0.5481608, 0.5504747, 0.5509398, 0.5474247, 0.5495819, 
    0.5426736, 0.5437872, 0.5431239, 0.5407052, 0.5484512, 0.5444697, 
    0.5518324, 0.5496675, 0.5559973, 0.5528452, 0.5590452, 0.5617067, 
    0.5642166, 0.5671582, 0.5425206, 0.5416792, 0.5431859, 0.5452742, 
    0.5472146, 0.5497994, 0.5500641, 0.5505492, 0.5518064, 0.5528646, 
    0.5507028, 0.55313, 0.544046, 0.5487974, 0.5413614, 0.5435959, 0.5451509, 
    0.5444683, 0.5480168, 0.5488548, 0.5522664, 0.5505014, 0.5610494, 
    0.5563705, 0.5694026, 0.5657451, 0.5413854, 0.5425176, 0.5464668, 
    0.5445861, 0.5499721, 0.5513018, 0.5523837, 0.5537686, 0.553918, 
    0.5547394, 0.5533938, 0.5546861, 0.5498049, 0.5519837, 0.5460144, 
    0.5474646, 0.5467972, 0.5460657, 0.5483248, 0.5507368, 0.5507881, 
    0.5515627, 0.5537488, 0.549994, 0.5616553, 0.5544399, 0.5437534, 0.54594, 
    0.5462523, 0.5454046, 0.5511684, 0.5490767, 0.5547193, 0.5531915, 
    0.5556958, 0.5544508, 0.5542676, 0.5526707, 0.5516777, 0.5491726, 
    0.5471383, 0.5455275, 0.5459018, 0.5476719, 0.5508845, 0.5539317, 
    0.5532635, 0.5555053, 0.5495808, 0.5520614, 0.5511021, 0.5536051, 
    0.5481274, 0.5527913, 0.5469384, 0.5474503, 0.5490353, 0.5522301, 
    0.5529377, 0.5536942, 0.5532272, 0.5509661, 0.5505959, 0.5489966, 
    0.5485556, 0.5473388, 0.5463325, 0.5472519, 0.5482184, 0.5509669, 
    0.5534497, 0.5561627, 0.5568274, 0.5600083, 0.5574187, 0.5616957, 
    0.558059, 0.5643616, 0.5530617, 0.5579516, 0.5491073, 0.5500568, 
    0.5517764, 0.5557296, 0.5535934, 0.556092, 0.5505814, 0.5477332, 
    0.546997, 0.5456254, 0.5470284, 0.5469142, 0.5482582, 0.5478261, 
    0.5510583, 0.549321, 0.5542632, 0.5560721, 0.5611962, 0.5643494, 
    0.5675681, 0.5689924, 0.5694262, 0.5696077,
  0.5840976, 0.5875086, 0.5868437, 0.5896073, 0.5880725, 0.5898846, 
    0.5847872, 0.5876446, 0.5858188, 0.5844036, 0.5950114, 0.5897309, 
    0.6005509, 0.5971422, 0.6057471, 0.6000192, 0.6069097, 0.6055806, 
    0.6095905, 0.6084385, 0.613603, 0.610123, 0.6163005, 0.6127695, 
    0.6133204, 0.6100087, 0.5907891, 0.5943512, 0.5905789, 0.5910851, 
    0.5908578, 0.5881042, 0.5867221, 0.5838375, 0.58436, 0.5864791, 
    0.5913129, 0.589667, 0.5938241, 0.5937299, 0.5983957, 0.596287, 
    0.6041912, 0.6019324, 0.6084865, 0.6068304, 0.6084087, 0.6079295, 
    0.6084149, 0.6059882, 0.6070265, 0.6048962, 0.5966813, 0.5990824, 
    0.5919532, 0.5877121, 0.5849124, 0.5829344, 0.5832136, 0.5837463, 
    0.5864915, 0.5890847, 0.5910693, 0.5924011, 0.5937164, 0.5977185, 
    0.5998483, 0.6046493, 0.6037793, 0.6052538, 0.6066659, 0.609046, 
    0.6086535, 0.6097049, 0.6052146, 0.6081945, 0.6032844, 0.6046228, 
    0.5940757, 0.5901105, 0.5884349, 0.5869715, 0.5834284, 0.5858728, 
    0.5849079, 0.587206, 0.5886714, 0.5879461, 0.5924375, 0.590687, 
    0.5999748, 0.5959544, 0.606501, 0.6039577, 0.6071125, 0.6055002, 
    0.6082659, 0.6057761, 0.6100966, 0.6110424, 0.6103959, 0.6128834, 
    0.6056384, 0.6084088, 0.5879259, 0.588044, 0.5885951, 0.5861772, 
    0.5860295, 0.5838232, 0.5857859, 0.5866238, 0.5887564, 0.5900219, 
    0.5912276, 0.593888, 0.5968752, 0.6010804, 0.6041222, 0.6061714, 
    0.6049138, 0.6060239, 0.6047831, 0.6042026, 0.6106879, 0.6070363, 
    0.6125249, 0.6122196, 0.6097299, 0.612254, 0.5881271, 0.587447, 
    0.5850927, 0.5869343, 0.5835835, 0.5854568, 0.5865368, 0.5907238, 
    0.5916477, 0.5925063, 0.5942057, 0.5963947, 0.6002568, 0.6036403, 
    0.6067482, 0.6065198, 0.6066002, 0.6072969, 0.6055729, 0.6075805, 
    0.6079184, 0.6070357, 0.6121787, 0.6107041, 0.6122131, 0.6112524, 
    0.5876679, 0.5888132, 0.5881941, 0.5893589, 0.5885381, 0.5921977, 
    0.5932998, 0.5984868, 0.5963516, 0.5997534, 0.5966961, 0.5972366, 
    0.5998653, 0.5968608, 0.6034534, 0.5989752, 0.6073241, 0.6028193, 
    0.6076077, 0.6067347, 0.6081808, 0.6094796, 0.6111181, 0.6141557, 
    0.6134506, 0.6160014, 0.5905248, 0.5920186, 0.5918867, 0.5934538, 
    0.5946159, 0.5971429, 0.6012216, 0.5996841, 0.60251, 0.6030792, 
    0.5987871, 0.6014184, 0.5930204, 0.5943686, 0.5935653, 0.5906426, 
    0.6000383, 0.5951958, 0.6041727, 0.601523, 0.6092943, 0.6054151, 
    0.613063, 0.6163687, 0.619499, 0.623184, 0.5928354, 0.5918184, 0.5936404, 
    0.5961721, 0.5985312, 0.6016843, 0.6020079, 0.6026012, 0.6041408, 
    0.6054389, 0.6027891, 0.6057648, 0.5946822, 0.6004606, 0.5914346, 
    0.5941368, 0.5960224, 0.5951942, 0.5995085, 0.6005306, 0.6047048, 
    0.6025427, 0.615551, 0.6097547, 0.6260078, 0.6214116, 0.5914636, 
    0.5928317, 0.5976212, 0.595337, 0.6018954, 0.6035225, 0.6048487, 
    0.6065495, 0.6067333, 0.607744, 0.6060889, 0.6076784, 0.6016911, 
    0.6043581, 0.5970713, 0.5988357, 0.5980232, 0.5971336, 0.5998841, 
    0.6028308, 0.6028935, 0.6038421, 0.6065252, 0.6019221, 0.6163048, 
    0.6073753, 0.5943276, 0.5969808, 0.5973604, 0.5963304, 0.6033591, 
    0.6008015, 0.6077192, 0.6058404, 0.6089224, 0.6073886, 0.6071634, 
    0.6052009, 0.603983, 0.6009186, 0.5984383, 0.5964796, 0.5969344, 
    0.5990883, 0.6030115, 0.6067501, 0.6059289, 0.6086875, 0.6014171, 
    0.6044534, 0.6032779, 0.6063486, 0.5996433, 0.6053489, 0.598195, 
    0.5988182, 0.6007509, 0.6046603, 0.6055287, 0.6064581, 0.6058843, 
    0.6031114, 0.6026583, 0.6007037, 0.6001655, 0.5986825, 0.5974579, 
    0.5985767, 0.5997543, 0.6031124, 0.6061576, 0.6094982, 0.6103189, 
    0.6142576, 0.6110495, 0.6163551, 0.6118417, 0.6196803, 0.6056809, 
    0.6117087, 0.6008388, 0.6019989, 0.604104, 0.6089641, 0.6063341, 
    0.609411, 0.6026406, 0.5991629, 0.5982664, 0.5965986, 0.5983046, 
    0.5981656, 0.5998029, 0.5992761, 0.6032243, 0.6010998, 0.6071578, 
    0.6093865, 0.6157336, 0.6196651, 0.623699, 0.6254908, 0.6260375, 0.6262662,
  0.6622251, 0.667787, 0.6666976, 0.6712429, 0.6687129, 0.6717016, 0.6633443, 
    0.6680101, 0.6650231, 0.6627214, 0.6802661, 0.6714472, 0.6897115, 
    0.6838751, 0.6987642, 0.6887959, 0.7008165, 0.6984711, 0.7055877, 
    0.7035307, 0.7128337, 0.7065421, 0.7177787, 0.711318, 0.7123192, 
    0.706337, 0.6732006, 0.679154, 0.6728517, 0.6736924, 0.6733148, 
    0.6687651, 0.6664985, 0.6618038, 0.6626507, 0.6661011, 0.6740712, 
    0.6713416, 0.6782681, 0.6781098, 0.6860123, 0.682423, 0.6960332, 
    0.6920996, 0.7036162, 0.7006762, 0.7034775, 0.7026251, 0.7034886, 
    0.6991889, 0.7010233, 0.6972684, 0.683092, 0.6871875, 0.6751375, 
    0.6681209, 0.6635476, 0.6603438, 0.6607947, 0.6616562, 0.6661214, 
    0.6703799, 0.6736662, 0.6758848, 0.6780871, 0.6848564, 0.688502, 
    0.6968355, 0.6953132, 0.6978964, 0.7003853, 0.7046142, 0.7039137, 
    0.7057924, 0.6978275, 0.7030964, 0.6944497, 0.696789, 0.6786907, 
    0.6720755, 0.669309, 0.6669068, 0.6611419, 0.6651114, 0.6635405, 
    0.6672908, 0.6696985, 0.6685052, 0.6759457, 0.6730312, 0.6887196, 
    0.6818596, 0.7000939, 0.6956249, 0.7011755, 0.6983296, 0.7032234, 
    0.6988153, 0.7064946, 0.7081949, 0.707032, 0.7115249, 0.6985729, 
    0.7034777, 0.6684719, 0.6686662, 0.6695728, 0.665608, 0.665367, 
    0.6617807, 0.6649695, 0.6663378, 0.6698384, 0.6719288, 0.6739292, 
    0.6783753, 0.6834213, 0.6906251, 0.6959125, 0.6995119, 0.6972994, 
    0.6992519, 0.6970701, 0.6960531, 0.7075568, 0.7010406, 0.7108743, 
    0.710321, 0.7058374, 0.7103833, 0.6688027, 0.6676859, 0.6638409, 
    0.6668458, 0.6613927, 0.6644333, 0.6661956, 0.6730922, 0.6746284, 
    0.6760606, 0.6789091, 0.6826057, 0.6892048, 0.6950704, 0.7005307, 
    0.7001271, 0.7002691, 0.7015024, 0.6984575, 0.7020053, 0.7026053, 
    0.7010396, 0.710247, 0.7075859, 0.7103093, 0.7085733, 0.6680484, 
    0.6699321, 0.6689128, 0.6708325, 0.6694789, 0.6755454, 0.6773884, 
    0.6861679, 0.6825325, 0.6883391, 0.683117, 0.6840357, 0.6885313, 
    0.6833967, 0.6947443, 0.6870038, 0.7015504, 0.6936398, 0.7020535, 
    0.7005069, 0.703072, 0.7053893, 0.7083312, 0.713842, 0.7125562, 
    0.7172273, 0.672762, 0.6752465, 0.6750265, 0.6776467, 0.6795995, 
    0.6838763, 0.6908692, 0.6882198, 0.6931019, 0.6940922, 0.6866817, 
    0.6912096, 0.6769205, 0.6791831, 0.6778337, 0.6729575, 0.6888287, 
    0.6805774, 0.6960008, 0.6913906, 0.7050577, 0.69818, 0.711851, 0.7179045, 
    0.7237219, 0.7306815, 0.6766108, 0.6749127, 0.6779597, 0.6822283, 
    0.6862438, 0.6916698, 0.6922304, 0.6932604, 0.6959449, 0.6982217, 
    0.6935872, 0.6987953, 0.6797112, 0.6895558, 0.6742736, 0.6787933, 
    0.6819748, 0.6805746, 0.6879184, 0.6896765, 0.6969327, 0.6931587, 
    0.7163987, 0.7058818, 0.7360995, 0.7273188, 0.6743218, 0.6766047, 
    0.6846905, 0.6808156, 0.6920354, 0.6948648, 0.6971852, 0.7001796, 
    0.7005044, 0.7022954, 0.6993665, 0.702179, 0.6916814, 0.6963252, 
    0.6837546, 0.6867649, 0.685376, 0.6838604, 0.6885635, 0.6936597, 
    0.6937689, 0.6954229, 0.7001367, 0.6920817, 0.7177866, 0.7016412, 
    0.6791143, 0.6836007, 0.6842464, 0.6824967, 0.6945799, 0.6901437, 
    0.7022516, 0.6989285, 0.7043934, 0.7016648, 0.7012656, 0.6978035, 
    0.6956691, 0.6903458, 0.6860851, 0.6827497, 0.6835218, 0.6871974, 
    0.6939742, 0.7005342, 0.6990844, 0.7039744, 0.6912072, 0.6964923, 
    0.6944383, 0.6998248, 0.6881498, 0.6980637, 0.6856694, 0.686735, 
    0.6900563, 0.6968548, 0.6983797, 0.7000182, 0.6990059, 0.6941482, 
    0.6933598, 0.689975, 0.6890477, 0.6865026, 0.6844125, 0.6863217, 
    0.6883404, 0.6941499, 0.6994876, 0.7054225, 0.7068936, 0.7140281, 
    0.7082077, 0.7178792, 0.7096372, 0.7240614, 0.6986477, 0.709397, 
    0.6902081, 0.6922148, 0.6958807, 0.7044679, 0.6997992, 0.7052665, 
    0.6933289, 0.6873254, 0.6857913, 0.6829515, 0.6858565, 0.6856191, 
    0.6884239, 0.6875196, 0.6943448, 0.6906587, 0.7012558, 0.7052227, 
    0.7167343, 0.7240329, 0.731664, 0.7351019, 0.7361569, 0.7365991,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.506774e-11, 3.522342e-11, 3.519307e-11, 3.531871e-11, 3.524898e-11, 
    3.533118e-11, 3.509911e-11, 3.522932e-11, 3.514615e-11, 3.508145e-11, 
    3.556242e-11, 3.532402e-11, 3.581065e-11, 3.565821e-11, 3.604128e-11, 
    3.578679e-11, 3.609261e-11, 3.603389e-11, 3.621064e-11, 3.615992e-11, 
    3.638605e-11, 3.623392e-11, 3.650343e-11, 3.634967e-11, 3.637364e-11, 
    3.622871e-11, 3.537228e-11, 3.553298e-11, 3.536268e-11, 3.53856e-11, 
    3.537528e-11, 3.525023e-11, 3.518724e-11, 3.505553e-11, 3.507938e-11, 
    3.517611e-11, 3.539562e-11, 3.532103e-11, 3.5509e-11, 3.550476e-11, 
    3.571422e-11, 3.561971e-11, 3.597232e-11, 3.587197e-11, 3.616199e-11, 
    3.608893e-11, 3.615848e-11, 3.613733e-11, 3.615864e-11, 3.605161e-11, 
    3.609737e-11, 3.600324e-11, 3.563785e-11, 3.574532e-11, 3.54248e-11, 
    3.523227e-11, 3.510466e-11, 3.501417e-11, 3.502687e-11, 3.505125e-11, 
    3.517659e-11, 3.529457e-11, 3.538455e-11, 3.544472e-11, 3.550403e-11, 
    3.568374e-11, 3.577902e-11, 3.59925e-11, 3.595397e-11, 3.601919e-11, 
    3.608163e-11, 3.618642e-11, 3.616915e-11, 3.621529e-11, 3.60173e-11, 
    3.614882e-11, 3.593168e-11, 3.599102e-11, 3.552038e-11, 3.534131e-11, 
    3.526512e-11, 3.519855e-11, 3.503667e-11, 3.514841e-11, 3.51043e-11, 
    3.520912e-11, 3.527575e-11, 3.524273e-11, 3.544632e-11, 3.536706e-11, 
    3.57846e-11, 3.560461e-11, 3.60744e-11, 3.596179e-11, 3.610128e-11, 
    3.603008e-11, 3.615201e-11, 3.60422e-11, 3.623242e-11, 3.627388e-11, 
    3.624546e-11, 3.635438e-11, 3.603587e-11, 3.615807e-11, 3.524202e-11, 
    3.524741e-11, 3.527242e-11, 3.516222e-11, 3.515548e-11, 3.505463e-11, 
    3.514428e-11, 3.518249e-11, 3.527953e-11, 3.533689e-11, 3.539146e-11, 
    3.551163e-11, 3.564585e-11, 3.583381e-11, 3.596904e-11, 3.605969e-11, 
    3.600405e-11, 3.605309e-11, 3.599818e-11, 3.597241e-11, 3.625822e-11, 
    3.609764e-11, 3.63386e-11, 3.632527e-11, 3.621608e-11, 3.632666e-11, 
    3.52511e-11, 3.522012e-11, 3.511271e-11, 3.519669e-11, 3.504359e-11, 
    3.512922e-11, 3.517842e-11, 3.536862e-11, 3.541045e-11, 3.544925e-11, 
    3.552588e-11, 3.562425e-11, 3.579706e-11, 3.594755e-11, 3.608512e-11, 
    3.607498e-11, 3.60785e-11, 3.610917e-11, 3.603302e-11, 3.61216e-11, 
    3.613642e-11, 3.609754e-11, 3.632336e-11, 3.62588e-11, 3.632483e-11, 
    3.628273e-11, 3.523013e-11, 3.528213e-11, 3.525395e-11, 3.530685e-11, 
    3.526949e-11, 3.54353e-11, 3.5485e-11, 3.571799e-11, 3.56223e-11, 
    3.577461e-11, 3.56377e-11, 3.566194e-11, 3.577937e-11, 3.5645e-11, 
    3.593909e-11, 3.573951e-11, 3.611033e-11, 3.591074e-11, 3.612276e-11, 
    3.608421e-11, 3.614791e-11, 3.620502e-11, 3.627683e-11, 3.640953e-11, 
    3.637872e-11, 3.648978e-11, 3.535975e-11, 3.542725e-11, 3.542132e-11, 
    3.549203e-11, 3.554432e-11, 3.565789e-11, 3.584011e-11, 3.57715e-11, 
    3.589736e-11, 3.592265e-11, 3.57313e-11, 3.584868e-11, 3.547212e-11, 
    3.553279e-11, 3.549664e-11, 3.536446e-11, 3.578692e-11, 3.556988e-11, 
    3.59708e-11, 3.585303e-11, 3.619676e-11, 3.602567e-11, 3.636177e-11, 
    3.65056e-11, 3.664118e-11, 3.679955e-11, 3.546414e-11, 3.541815e-11, 
    3.550037e-11, 3.561423e-11, 3.571994e-11, 3.586067e-11, 3.587504e-11, 
    3.590135e-11, 3.596966e-11, 3.602715e-11, 3.590956e-11, 3.604145e-11, 
    3.554676e-11, 3.580578e-11, 3.540025e-11, 3.55222e-11, 3.560699e-11, 
    3.556979e-11, 3.576317e-11, 3.580872e-11, 3.599414e-11, 3.589827e-11, 
    3.646994e-11, 3.621674e-11, 3.692032e-11, 3.672338e-11, 3.540205e-11, 
    3.546383e-11, 3.567914e-11, 3.557665e-11, 3.586997e-11, 3.594227e-11, 
    3.6001e-11, 3.607617e-11, 3.608423e-11, 3.61288e-11, 3.60557e-11, 
    3.612585e-11, 3.586055e-11, 3.597903e-11, 3.565413e-11, 3.573306e-11, 
    3.569671e-11, 3.565679e-11, 3.57798e-11, 3.591096e-11, 3.591378e-11, 
    3.595578e-11, 3.607427e-11, 3.587045e-11, 3.650239e-11, 3.611167e-11, 
    3.553124e-11, 3.565034e-11, 3.566739e-11, 3.562121e-11, 3.593491e-11, 
    3.582114e-11, 3.612772e-11, 3.604474e-11, 3.618058e-11, 3.611305e-11, 
    3.610302e-11, 3.601634e-11, 3.596229e-11, 3.582604e-11, 3.571519e-11, 
    3.562746e-11, 3.564778e-11, 3.574419e-11, 3.591889e-11, 3.608447e-11, 
    3.604812e-11, 3.616977e-11, 3.584789e-11, 3.598274e-11, 3.59305e-11, 
    3.606653e-11, 3.576951e-11, 3.602293e-11, 3.570473e-11, 3.573255e-11, 
    3.581877e-11, 3.599243e-11, 3.603088e-11, 3.607193e-11, 3.604653e-11, 
    3.592363e-11, 3.590347e-11, 3.581643e-11, 3.579235e-11, 3.572614e-11, 
    3.567123e-11, 3.572131e-11, 3.577382e-11, 3.59234e-11, 3.605822e-11, 
    3.620534e-11, 3.624139e-11, 3.641335e-11, 3.627321e-11, 3.650437e-11, 
    3.630763e-11, 3.664831e-11, 3.60376e-11, 3.630276e-11, 3.582273e-11, 
    3.587432e-11, 3.596772e-11, 3.618223e-11, 3.606637e-11, 3.620185e-11, 
    3.590267e-11, 3.574755e-11, 3.570748e-11, 3.563273e-11, 3.570911e-11, 
    3.57029e-11, 3.577605e-11, 3.575247e-11, 3.592825e-11, 3.583379e-11, 
    3.610224e-11, 3.620034e-11, 3.647767e-11, 3.664783e-11, 3.682134e-11, 
    3.689792e-11, 3.692124e-11, 3.693094e-11,
  1.781549e-11, 1.79512e-11, 1.79248e-11, 1.803447e-11, 1.797361e-11, 
    1.804547e-11, 1.784298e-11, 1.795659e-11, 1.788404e-11, 1.78277e-11, 
    1.824801e-11, 1.803938e-11, 1.846581e-11, 1.833202e-11, 1.866883e-11, 
    1.844495e-11, 1.87141e-11, 1.866239e-11, 1.881827e-11, 1.877357e-11, 
    1.897341e-11, 1.883892e-11, 1.907735e-11, 1.894127e-11, 1.896253e-11, 
    1.883448e-11, 1.808132e-11, 1.822198e-11, 1.807299e-11, 1.809302e-11, 
    1.808404e-11, 1.797486e-11, 1.791992e-11, 1.780515e-11, 1.782597e-11, 
    1.791028e-11, 1.810203e-11, 1.803687e-11, 1.820131e-11, 1.819759e-11, 
    1.83813e-11, 1.829838e-11, 1.860821e-11, 1.851996e-11, 1.877543e-11, 
    1.871106e-11, 1.87724e-11, 1.87538e-11, 1.877264e-11, 1.867827e-11, 
    1.871868e-11, 1.863572e-11, 1.83139e-11, 1.840825e-11, 1.812737e-11, 
    1.795923e-11, 1.784795e-11, 1.776913e-11, 1.778027e-11, 1.780149e-11, 
    1.791078e-11, 1.801378e-11, 1.809242e-11, 1.81451e-11, 1.819706e-11, 
    1.835461e-11, 1.843827e-11, 1.862606e-11, 1.859214e-11, 1.864964e-11, 
    1.870466e-11, 1.879714e-11, 1.878191e-11, 1.882269e-11, 1.864814e-11, 
    1.876407e-11, 1.857283e-11, 1.862506e-11, 1.82111e-11, 1.805445e-11, 
    1.798794e-11, 1.792987e-11, 1.778883e-11, 1.788618e-11, 1.784777e-11, 
    1.793921e-11, 1.799738e-11, 1.796861e-11, 1.814654e-11, 1.807728e-11, 
    1.844323e-11, 1.828526e-11, 1.869824e-11, 1.85991e-11, 1.872203e-11, 
    1.865927e-11, 1.876685e-11, 1.867002e-11, 1.883788e-11, 1.88745e-11, 
    1.884947e-11, 1.89457e-11, 1.866466e-11, 1.877239e-11, 1.79678e-11, 
    1.797249e-11, 1.799436e-11, 1.789828e-11, 1.789241e-11, 1.780457e-11, 
    1.788273e-11, 1.791605e-11, 1.800077e-11, 1.805093e-11, 1.809868e-11, 
    1.820382e-11, 1.83215e-11, 1.848657e-11, 1.860553e-11, 1.868541e-11, 
    1.863642e-11, 1.867967e-11, 1.863132e-11, 1.860868e-11, 1.886077e-11, 
    1.871905e-11, 1.893185e-11, 1.892005e-11, 1.882365e-11, 1.892138e-11, 
    1.797578e-11, 1.794879e-11, 1.785514e-11, 1.792841e-11, 1.779502e-11, 
    1.786963e-11, 1.791257e-11, 1.807871e-11, 1.811531e-11, 1.814924e-11, 
    1.821636e-11, 1.830262e-11, 1.845431e-11, 1.858669e-11, 1.870787e-11, 
    1.869898e-11, 1.870211e-11, 1.87292e-11, 1.86621e-11, 1.874023e-11, 
    1.875334e-11, 1.871905e-11, 1.891847e-11, 1.886142e-11, 1.89198e-11, 
    1.888265e-11, 1.795756e-11, 1.800301e-11, 1.797845e-11, 1.802465e-11, 
    1.799209e-11, 1.813701e-11, 1.818055e-11, 1.838484e-11, 1.830092e-11, 
    1.843457e-11, 1.831449e-11, 1.833574e-11, 1.843889e-11, 1.832097e-11, 
    1.857937e-11, 1.8404e-11, 1.873026e-11, 1.855456e-11, 1.874128e-11, 
    1.870734e-11, 1.876356e-11, 1.881396e-11, 1.887745e-11, 1.899477e-11, 
    1.896758e-11, 1.906587e-11, 1.807086e-11, 1.812995e-11, 1.812476e-11, 
    1.818669e-11, 1.823253e-11, 1.833207e-11, 1.849212e-11, 1.843188e-11, 
    1.854255e-11, 1.85648e-11, 1.839669e-11, 1.849982e-11, 1.816955e-11, 
    1.822274e-11, 1.819108e-11, 1.807551e-11, 1.844573e-11, 1.825536e-11, 
    1.860749e-11, 1.850393e-11, 1.880677e-11, 1.865591e-11, 1.895262e-11, 
    1.907994e-11, 1.920013e-11, 1.934084e-11, 1.816225e-11, 1.812206e-11, 
    1.819406e-11, 1.829382e-11, 1.838662e-11, 1.851024e-11, 1.852291e-11, 
    1.854611e-11, 1.860626e-11, 1.865688e-11, 1.855343e-11, 1.866958e-11, 
    1.823505e-11, 1.84623e-11, 1.810686e-11, 1.821359e-11, 1.828794e-11, 
    1.825533e-11, 1.8425e-11, 1.846507e-11, 1.862823e-11, 1.854383e-11, 
    1.904847e-11, 1.882458e-11, 1.944829e-11, 1.927324e-11, 1.810802e-11, 
    1.816212e-11, 1.835085e-11, 1.826096e-11, 1.851851e-11, 1.858211e-11, 
    1.863388e-11, 1.870011e-11, 1.870728e-11, 1.874657e-11, 1.86822e-11, 
    1.874404e-11, 1.85105e-11, 1.861473e-11, 1.832926e-11, 1.839858e-11, 
    1.836668e-11, 1.833171e-11, 1.843973e-11, 1.855505e-11, 1.855754e-11, 
    1.859458e-11, 1.869902e-11, 1.851956e-11, 1.907738e-11, 1.873211e-11, 
    1.822118e-11, 1.832564e-11, 1.834062e-11, 1.83001e-11, 1.857573e-11, 
    1.847568e-11, 1.874562e-11, 1.867253e-11, 1.879235e-11, 1.873277e-11, 
    1.872401e-11, 1.864761e-11, 1.860009e-11, 1.848025e-11, 1.838297e-11, 
    1.830598e-11, 1.832387e-11, 1.840848e-11, 1.856212e-11, 1.870792e-11, 
    1.867594e-11, 1.878324e-11, 1.849979e-11, 1.861843e-11, 1.857253e-11, 
    1.869231e-11, 1.843027e-11, 1.865323e-11, 1.837344e-11, 1.839791e-11, 
    1.847369e-11, 1.862647e-11, 1.866038e-11, 1.869656e-11, 1.867424e-11, 
    1.856603e-11, 1.854834e-11, 1.847186e-11, 1.845075e-11, 1.839258e-11, 
    1.834447e-11, 1.838842e-11, 1.843461e-11, 1.856609e-11, 1.868485e-11, 
    1.881467e-11, 1.88465e-11, 1.899862e-11, 1.887471e-11, 1.90793e-11, 
    1.890525e-11, 1.920694e-11, 1.866623e-11, 1.89002e-11, 1.847715e-11, 
    1.852256e-11, 1.860478e-11, 1.879391e-11, 1.869174e-11, 1.881126e-11, 
    1.854765e-11, 1.841139e-11, 1.837624e-11, 1.831065e-11, 1.837774e-11, 
    1.837228e-11, 1.843655e-11, 1.841589e-11, 1.857046e-11, 1.848737e-11, 
    1.872378e-11, 1.881032e-11, 1.905555e-11, 1.920644e-11, 1.936053e-11, 
    1.942868e-11, 1.944944e-11, 1.945812e-11,
  1.677788e-11, 1.692675e-11, 1.689777e-11, 1.701816e-11, 1.695133e-11, 
    1.703023e-11, 1.680802e-11, 1.693266e-11, 1.685305e-11, 1.679126e-11, 
    1.725282e-11, 1.702354e-11, 1.749245e-11, 1.734519e-11, 1.771615e-11, 
    1.746949e-11, 1.776607e-11, 1.770903e-11, 1.788097e-11, 1.783165e-11, 
    1.80523e-11, 1.790376e-11, 1.816716e-11, 1.801679e-11, 1.804027e-11, 
    1.789887e-11, 1.706959e-11, 1.72242e-11, 1.706045e-11, 1.708245e-11, 
    1.707258e-11, 1.695271e-11, 1.689243e-11, 1.676653e-11, 1.678936e-11, 
    1.688185e-11, 1.709235e-11, 1.702078e-11, 1.720144e-11, 1.719735e-11, 
    1.739941e-11, 1.730818e-11, 1.764931e-11, 1.755207e-11, 1.78337e-11, 
    1.776269e-11, 1.783036e-11, 1.780984e-11, 1.783063e-11, 1.772654e-11, 
    1.77711e-11, 1.767963e-11, 1.732524e-11, 1.742907e-11, 1.712019e-11, 
    1.693558e-11, 1.681347e-11, 1.672705e-11, 1.673926e-11, 1.676253e-11, 
    1.688239e-11, 1.699543e-11, 1.708179e-11, 1.713966e-11, 1.719676e-11, 
    1.737006e-11, 1.746213e-11, 1.766899e-11, 1.76316e-11, 1.769498e-11, 
    1.775564e-11, 1.785766e-11, 1.784085e-11, 1.788585e-11, 1.769332e-11, 
    1.782117e-11, 1.761031e-11, 1.766787e-11, 1.721224e-11, 1.704008e-11, 
    1.696708e-11, 1.690333e-11, 1.674864e-11, 1.68554e-11, 1.681328e-11, 
    1.691357e-11, 1.697743e-11, 1.694584e-11, 1.714124e-11, 1.706516e-11, 
    1.746759e-11, 1.729376e-11, 1.774856e-11, 1.763927e-11, 1.77748e-11, 
    1.770559e-11, 1.782424e-11, 1.771744e-11, 1.790262e-11, 1.794305e-11, 
    1.791542e-11, 1.802167e-11, 1.771153e-11, 1.783036e-11, 1.694495e-11, 
    1.69501e-11, 1.697411e-11, 1.686868e-11, 1.686224e-11, 1.67659e-11, 
    1.685162e-11, 1.688817e-11, 1.698114e-11, 1.703622e-11, 1.708866e-11, 
    1.72042e-11, 1.733362e-11, 1.751531e-11, 1.764635e-11, 1.773441e-11, 
    1.768039e-11, 1.772808e-11, 1.767477e-11, 1.764981e-11, 1.792789e-11, 
    1.777152e-11, 1.800637e-11, 1.799334e-11, 1.788692e-11, 1.799481e-11, 
    1.695372e-11, 1.692409e-11, 1.682136e-11, 1.690173e-11, 1.675543e-11, 
    1.683724e-11, 1.688436e-11, 1.706673e-11, 1.710693e-11, 1.714422e-11, 
    1.721798e-11, 1.731284e-11, 1.747978e-11, 1.76256e-11, 1.775917e-11, 
    1.774937e-11, 1.775282e-11, 1.778271e-11, 1.770871e-11, 1.779487e-11, 
    1.780934e-11, 1.77715e-11, 1.79916e-11, 1.79286e-11, 1.799307e-11, 
    1.795204e-11, 1.693372e-11, 1.698361e-11, 1.695664e-11, 1.700736e-11, 
    1.697162e-11, 1.713079e-11, 1.717864e-11, 1.740331e-11, 1.731097e-11, 
    1.745805e-11, 1.732589e-11, 1.734927e-11, 1.746283e-11, 1.733302e-11, 
    1.761753e-11, 1.742441e-11, 1.778387e-11, 1.759021e-11, 1.779603e-11, 
    1.775859e-11, 1.782061e-11, 1.787622e-11, 1.79463e-11, 1.807589e-11, 
    1.804585e-11, 1.815446e-11, 1.70581e-11, 1.712302e-11, 1.711731e-11, 
    1.718536e-11, 1.723576e-11, 1.734523e-11, 1.752141e-11, 1.745508e-11, 
    1.757696e-11, 1.760146e-11, 1.741634e-11, 1.752989e-11, 1.716654e-11, 
    1.722501e-11, 1.719019e-11, 1.706321e-11, 1.747034e-11, 1.726088e-11, 
    1.764851e-11, 1.753442e-11, 1.786828e-11, 1.77019e-11, 1.802932e-11, 
    1.817002e-11, 1.830293e-11, 1.845869e-11, 1.715851e-11, 1.711435e-11, 
    1.719347e-11, 1.730317e-11, 1.740526e-11, 1.754136e-11, 1.755532e-11, 
    1.758088e-11, 1.764715e-11, 1.770295e-11, 1.758895e-11, 1.771695e-11, 
    1.723856e-11, 1.748857e-11, 1.709765e-11, 1.721495e-11, 1.72967e-11, 
    1.726083e-11, 1.744751e-11, 1.749162e-11, 1.767138e-11, 1.757837e-11, 
    1.813524e-11, 1.788796e-11, 1.85777e-11, 1.838384e-11, 1.709892e-11, 
    1.715836e-11, 1.73659e-11, 1.726702e-11, 1.755047e-11, 1.762054e-11, 
    1.76776e-11, 1.775063e-11, 1.775853e-11, 1.780187e-11, 1.773087e-11, 
    1.779907e-11, 1.754166e-11, 1.765649e-11, 1.734214e-11, 1.741842e-11, 
    1.738332e-11, 1.734483e-11, 1.746372e-11, 1.759074e-11, 1.759347e-11, 
    1.763428e-11, 1.774947e-11, 1.755163e-11, 1.816723e-11, 1.778596e-11, 
    1.722328e-11, 1.733818e-11, 1.735464e-11, 1.731007e-11, 1.761351e-11, 
    1.75033e-11, 1.780082e-11, 1.77202e-11, 1.785237e-11, 1.778664e-11, 
    1.777698e-11, 1.769273e-11, 1.764036e-11, 1.750834e-11, 1.740125e-11, 
    1.731653e-11, 1.733622e-11, 1.742933e-11, 1.759852e-11, 1.775924e-11, 
    1.772398e-11, 1.784231e-11, 1.752985e-11, 1.766058e-11, 1.761e-11, 
    1.774202e-11, 1.745331e-11, 1.769898e-11, 1.739075e-11, 1.741768e-11, 
    1.750112e-11, 1.766945e-11, 1.770681e-11, 1.774671e-11, 1.772209e-11, 
    1.760283e-11, 1.758333e-11, 1.749909e-11, 1.747585e-11, 1.741182e-11, 
    1.735887e-11, 1.740724e-11, 1.745809e-11, 1.760289e-11, 1.77338e-11, 
    1.787701e-11, 1.791214e-11, 1.808017e-11, 1.794331e-11, 1.816936e-11, 
    1.797706e-11, 1.83105e-11, 1.771329e-11, 1.797145e-11, 1.750492e-11, 
    1.755493e-11, 1.764553e-11, 1.785411e-11, 1.77414e-11, 1.787325e-11, 
    1.758257e-11, 1.743254e-11, 1.739383e-11, 1.732167e-11, 1.739548e-11, 
    1.738947e-11, 1.746021e-11, 1.743747e-11, 1.760771e-11, 1.751617e-11, 
    1.777673e-11, 1.787221e-11, 1.814305e-11, 1.830992e-11, 1.848047e-11, 
    1.855596e-11, 1.857897e-11, 1.858859e-11,
  1.721998e-11, 1.738378e-11, 1.735188e-11, 1.748443e-11, 1.741085e-11, 
    1.749772e-11, 1.725313e-11, 1.73903e-11, 1.730267e-11, 1.72347e-11, 
    1.774304e-11, 1.749035e-11, 1.80074e-11, 1.784488e-11, 1.825451e-11, 
    1.798206e-11, 1.830969e-11, 1.824663e-11, 1.843675e-11, 1.838219e-11, 
    1.862639e-11, 1.846196e-11, 1.87536e-11, 1.858707e-11, 1.861307e-11, 
    1.845655e-11, 1.754107e-11, 1.771148e-11, 1.7531e-11, 1.755524e-11, 
    1.754436e-11, 1.741236e-11, 1.734602e-11, 1.72075e-11, 1.723261e-11, 
    1.733437e-11, 1.756615e-11, 1.748731e-11, 1.768635e-11, 1.768185e-11, 
    1.79047e-11, 1.780405e-11, 1.818063e-11, 1.807321e-11, 1.838447e-11, 
    1.830595e-11, 1.838077e-11, 1.835807e-11, 1.838107e-11, 1.826598e-11, 
    1.831525e-11, 1.821413e-11, 1.782288e-11, 1.793743e-11, 1.759681e-11, 
    1.739352e-11, 1.725914e-11, 1.716408e-11, 1.71775e-11, 1.72031e-11, 
    1.733497e-11, 1.745939e-11, 1.75545e-11, 1.761826e-11, 1.76812e-11, 
    1.787234e-11, 1.797393e-11, 1.820239e-11, 1.816106e-11, 1.82311e-11, 
    1.829815e-11, 1.841096e-11, 1.839237e-11, 1.844216e-11, 1.822926e-11, 
    1.837062e-11, 1.813754e-11, 1.820115e-11, 1.76983e-11, 1.750856e-11, 
    1.742819e-11, 1.735801e-11, 1.718783e-11, 1.730526e-11, 1.725892e-11, 
    1.736928e-11, 1.743957e-11, 1.740479e-11, 1.762001e-11, 1.753618e-11, 
    1.797996e-11, 1.778815e-11, 1.829032e-11, 1.816954e-11, 1.831933e-11, 
    1.824282e-11, 1.8374e-11, 1.825592e-11, 1.846071e-11, 1.850544e-11, 
    1.847487e-11, 1.859246e-11, 1.824938e-11, 1.838077e-11, 1.740381e-11, 
    1.740948e-11, 1.743592e-11, 1.731987e-11, 1.731279e-11, 1.720681e-11, 
    1.73011e-11, 1.734132e-11, 1.744365e-11, 1.750432e-11, 1.756208e-11, 
    1.76894e-11, 1.783212e-11, 1.803263e-11, 1.817736e-11, 1.827468e-11, 
    1.821497e-11, 1.826768e-11, 1.820877e-11, 1.818118e-11, 1.848867e-11, 
    1.831571e-11, 1.857553e-11, 1.85611e-11, 1.844334e-11, 1.856273e-11, 
    1.741347e-11, 1.738085e-11, 1.726781e-11, 1.735624e-11, 1.719528e-11, 
    1.728529e-11, 1.733714e-11, 1.753793e-11, 1.75822e-11, 1.762329e-11, 
    1.770459e-11, 1.780919e-11, 1.799341e-11, 1.815444e-11, 1.830205e-11, 
    1.829122e-11, 1.829503e-11, 1.832808e-11, 1.824627e-11, 1.834152e-11, 
    1.835753e-11, 1.831569e-11, 1.855917e-11, 1.848945e-11, 1.85608e-11, 
    1.851539e-11, 1.739145e-11, 1.744637e-11, 1.741668e-11, 1.747253e-11, 
    1.743317e-11, 1.760851e-11, 1.766124e-11, 1.790901e-11, 1.780713e-11, 
    1.796942e-11, 1.782359e-11, 1.784938e-11, 1.797472e-11, 1.783145e-11, 
    1.814554e-11, 1.79323e-11, 1.832936e-11, 1.811537e-11, 1.834281e-11, 
    1.830141e-11, 1.836998e-11, 1.84315e-11, 1.850903e-11, 1.86525e-11, 
    1.861923e-11, 1.873953e-11, 1.752841e-11, 1.759994e-11, 1.759364e-11, 
    1.766864e-11, 1.77242e-11, 1.784492e-11, 1.803937e-11, 1.796613e-11, 
    1.81007e-11, 1.812777e-11, 1.792337e-11, 1.804873e-11, 1.764789e-11, 
    1.771236e-11, 1.767396e-11, 1.753405e-11, 1.798299e-11, 1.77519e-11, 
    1.817975e-11, 1.805373e-11, 1.842272e-11, 1.823876e-11, 1.860093e-11, 
    1.875679e-11, 1.890408e-11, 1.907688e-11, 1.763904e-11, 1.759037e-11, 
    1.767757e-11, 1.779854e-11, 1.791116e-11, 1.80614e-11, 1.807681e-11, 
    1.810503e-11, 1.817824e-11, 1.823991e-11, 1.811396e-11, 1.825538e-11, 
    1.772731e-11, 1.800312e-11, 1.757199e-11, 1.770127e-11, 1.77914e-11, 
    1.775184e-11, 1.795777e-11, 1.800647e-11, 1.820503e-11, 1.810226e-11, 
    1.871826e-11, 1.84445e-11, 1.920897e-11, 1.899382e-11, 1.757338e-11, 
    1.763888e-11, 1.786773e-11, 1.775867e-11, 1.807145e-11, 1.814885e-11, 
    1.821189e-11, 1.829261e-11, 1.830134e-11, 1.834927e-11, 1.827077e-11, 
    1.834616e-11, 1.806172e-11, 1.818857e-11, 1.784151e-11, 1.792568e-11, 
    1.788693e-11, 1.784448e-11, 1.797567e-11, 1.811593e-11, 1.811894e-11, 
    1.816404e-11, 1.829138e-11, 1.807273e-11, 1.875373e-11, 1.833171e-11, 
    1.771043e-11, 1.783715e-11, 1.78553e-11, 1.780613e-11, 1.814108e-11, 
    1.801937e-11, 1.83481e-11, 1.825897e-11, 1.840512e-11, 1.833242e-11, 
    1.832174e-11, 1.822861e-11, 1.817074e-11, 1.802494e-11, 1.790673e-11, 
    1.781326e-11, 1.783497e-11, 1.793772e-11, 1.812453e-11, 1.830213e-11, 
    1.826315e-11, 1.839399e-11, 1.804868e-11, 1.819309e-11, 1.813721e-11, 
    1.828309e-11, 1.796419e-11, 1.823556e-11, 1.789513e-11, 1.792486e-11, 
    1.801695e-11, 1.82029e-11, 1.824417e-11, 1.828828e-11, 1.826106e-11, 
    1.812929e-11, 1.810775e-11, 1.801471e-11, 1.798907e-11, 1.791838e-11, 
    1.785997e-11, 1.791333e-11, 1.796946e-11, 1.812935e-11, 1.827401e-11, 
    1.843237e-11, 1.847123e-11, 1.865726e-11, 1.850575e-11, 1.875609e-11, 
    1.854314e-11, 1.891252e-11, 1.825136e-11, 1.85369e-11, 1.802115e-11, 
    1.807638e-11, 1.817647e-11, 1.840706e-11, 1.82824e-11, 1.842823e-11, 
    1.81069e-11, 1.794126e-11, 1.789854e-11, 1.781893e-11, 1.790036e-11, 
    1.789373e-11, 1.79718e-11, 1.794669e-11, 1.813467e-11, 1.803358e-11, 
    1.832147e-11, 1.842708e-11, 1.87269e-11, 1.891185e-11, 1.910102e-11, 
    1.918483e-11, 1.921037e-11, 1.922105e-11,
  1.87948e-11, 1.897033e-11, 1.893613e-11, 1.907825e-11, 1.899934e-11, 
    1.90925e-11, 1.883031e-11, 1.897732e-11, 1.888339e-11, 1.881056e-11, 
    1.93558e-11, 1.90846e-11, 1.963983e-11, 1.946515e-11, 1.990568e-11, 
    1.961259e-11, 1.996508e-11, 1.989718e-11, 2.010193e-11, 2.004315e-11, 
    2.030639e-11, 2.01291e-11, 2.044363e-11, 2.026396e-11, 2.029201e-11, 
    2.012327e-11, 1.9139e-11, 1.932192e-11, 1.912819e-11, 1.91542e-11, 
    1.914253e-11, 1.900096e-11, 1.892986e-11, 1.878142e-11, 1.880832e-11, 
    1.891736e-11, 1.916591e-11, 1.908133e-11, 1.92949e-11, 1.929006e-11, 
    1.952942e-11, 1.942129e-11, 1.982615e-11, 1.971059e-11, 2.00456e-11, 
    1.996104e-11, 2.004163e-11, 2.001717e-11, 2.004195e-11, 1.991801e-11, 
    1.997106e-11, 1.98622e-11, 1.944151e-11, 1.956461e-11, 1.919881e-11, 
    1.898078e-11, 1.883674e-11, 1.873492e-11, 1.87493e-11, 1.877672e-11, 
    1.8918e-11, 1.905139e-11, 1.91534e-11, 1.922182e-11, 1.928937e-11, 
    1.949468e-11, 1.960384e-11, 1.984957e-11, 1.980509e-11, 1.988047e-11, 
    1.995264e-11, 2.007415e-11, 2.005412e-11, 2.010776e-11, 1.987848e-11, 
    2.003069e-11, 1.977978e-11, 1.984822e-11, 1.930777e-11, 1.910412e-11, 
    1.901796e-11, 1.89427e-11, 1.876035e-11, 1.888617e-11, 1.883652e-11, 
    1.895477e-11, 1.903014e-11, 1.899284e-11, 1.922369e-11, 1.913375e-11, 
    1.961033e-11, 1.940422e-11, 1.994421e-11, 1.981421e-11, 1.997545e-11, 
    1.989308e-11, 2.003434e-11, 1.990718e-11, 2.012775e-11, 2.017597e-11, 
    2.014301e-11, 2.026978e-11, 1.990014e-11, 2.004163e-11, 1.89918e-11, 
    1.899787e-11, 1.902621e-11, 1.890183e-11, 1.889424e-11, 1.878068e-11, 
    1.88817e-11, 1.892481e-11, 1.903451e-11, 1.909957e-11, 1.916153e-11, 
    1.929817e-11, 1.945145e-11, 1.966695e-11, 1.982262e-11, 1.992737e-11, 
    1.98631e-11, 1.991984e-11, 1.985642e-11, 1.982674e-11, 2.015789e-11, 
    1.997155e-11, 2.025151e-11, 2.023596e-11, 2.010904e-11, 2.023771e-11, 
    1.900215e-11, 1.896717e-11, 1.884603e-11, 1.894079e-11, 1.876834e-11, 
    1.886476e-11, 1.892034e-11, 1.913563e-11, 1.918312e-11, 1.922722e-11, 
    1.931448e-11, 1.942681e-11, 1.962478e-11, 1.979797e-11, 1.995684e-11, 
    1.994518e-11, 1.994928e-11, 1.998487e-11, 1.989679e-11, 1.999935e-11, 
    2.00166e-11, 1.997153e-11, 2.023388e-11, 2.015873e-11, 2.023563e-11, 
    2.018668e-11, 1.897853e-11, 1.903743e-11, 1.900559e-11, 1.906548e-11, 
    1.902328e-11, 1.921136e-11, 1.926796e-11, 1.953407e-11, 1.94246e-11, 
    1.959899e-11, 1.944227e-11, 1.946999e-11, 1.96047e-11, 1.945072e-11, 
    1.97884e-11, 1.95591e-11, 1.998625e-11, 1.975595e-11, 2.000074e-11, 
    1.995615e-11, 2.003e-11, 2.009628e-11, 2.017983e-11, 2.033454e-11, 
    2.029865e-11, 2.042843e-11, 1.912541e-11, 1.920216e-11, 1.91954e-11, 
    1.927588e-11, 1.933554e-11, 1.946519e-11, 1.967419e-11, 1.959545e-11, 
    1.974015e-11, 1.976927e-11, 1.954949e-11, 1.968427e-11, 1.925362e-11, 
    1.932283e-11, 1.928161e-11, 1.913147e-11, 1.961358e-11, 1.936529e-11, 
    1.98252e-11, 1.968963e-11, 2.008682e-11, 1.988872e-11, 2.027891e-11, 
    2.044708e-11, 2.060608e-11, 2.079283e-11, 1.924412e-11, 1.919189e-11, 
    1.928547e-11, 1.941538e-11, 1.953636e-11, 1.969788e-11, 1.971445e-11, 
    1.974481e-11, 1.982358e-11, 1.988994e-11, 1.975442e-11, 1.99066e-11, 
    1.933891e-11, 1.963522e-11, 1.917217e-11, 1.931093e-11, 1.940771e-11, 
    1.936522e-11, 1.958646e-11, 1.963881e-11, 1.985241e-11, 1.974182e-11, 
    2.04055e-11, 2.01103e-11, 2.093567e-11, 2.070306e-11, 1.917366e-11, 
    1.924394e-11, 1.948971e-11, 1.937255e-11, 1.970869e-11, 1.979195e-11, 
    1.985978e-11, 1.994669e-11, 1.995608e-11, 2.000769e-11, 1.992316e-11, 
    2.000435e-11, 1.969823e-11, 1.983469e-11, 1.946152e-11, 1.955197e-11, 
    1.951033e-11, 1.946471e-11, 1.96057e-11, 1.975655e-11, 1.975978e-11, 
    1.980829e-11, 1.99454e-11, 1.971006e-11, 2.04438e-11, 1.998883e-11, 
    1.932075e-11, 1.945686e-11, 1.947634e-11, 1.942352e-11, 1.978359e-11, 
    1.965268e-11, 2.000643e-11, 1.991046e-11, 2.006785e-11, 1.998955e-11, 
    1.997805e-11, 1.987778e-11, 1.981551e-11, 1.965868e-11, 1.95316e-11, 
    1.943117e-11, 1.94545e-11, 1.956491e-11, 1.97658e-11, 1.995694e-11, 
    1.991498e-11, 2.005586e-11, 1.968421e-11, 1.983956e-11, 1.977943e-11, 
    1.993643e-11, 1.959336e-11, 1.98853e-11, 1.951914e-11, 1.955108e-11, 
    1.965009e-11, 1.985013e-11, 1.989453e-11, 1.994202e-11, 1.991271e-11, 
    1.977091e-11, 1.974773e-11, 1.964768e-11, 1.962011e-11, 1.954412e-11, 
    1.948135e-11, 1.95387e-11, 1.959904e-11, 1.977097e-11, 1.992666e-11, 
    2.009722e-11, 2.013909e-11, 2.03397e-11, 2.017631e-11, 2.044635e-11, 
    2.021665e-11, 2.061524e-11, 1.990229e-11, 2.02099e-11, 1.96546e-11, 
    1.971399e-11, 1.982168e-11, 2.006995e-11, 1.993569e-11, 2.009276e-11, 
    1.974683e-11, 1.956873e-11, 1.952279e-11, 1.943727e-11, 1.952475e-11, 
    1.951763e-11, 1.960153e-11, 1.957455e-11, 1.977669e-11, 1.966796e-11, 
    1.997776e-11, 2.009152e-11, 2.041481e-11, 2.061449e-11, 2.081892e-11, 
    2.090955e-11, 2.093718e-11, 2.094874e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
