netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to patch-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to patch-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "patch-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total patch-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float RSCANOPY(time, lndgrid) ;
		RSCANOPY:long_name = "canopy resistance" ;
		RSCANOPY:units = " s m-1" ;
		RSCANOPY:cell_methods = "time: mean" ;
		RSCANOPY:_FillValue = 1.e+36f ;
		RSCANOPY:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new Patches" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total patch-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C eallocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 11/05/14 11:51:47" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "11/05/14" ;

 time_written =
  "11:51:47" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.059954e-14, 5.073669e-14, 5.071005e-14, 5.082057e-14, 5.075929e-14, 
    5.083163e-14, 5.062738e-14, 5.074212e-14, 5.066889e-14, 5.061192e-14, 
    5.103474e-14, 5.082551e-14, 5.125189e-14, 5.111869e-14, 5.145308e-14, 
    5.123114e-14, 5.149779e-14, 5.144673e-14, 5.160045e-14, 5.155644e-14, 
    5.175276e-14, 5.162077e-14, 5.185447e-14, 5.172128e-14, 5.174211e-14, 
    5.16164e-14, 5.086768e-14, 5.10087e-14, 5.085931e-14, 5.087943e-14, 
    5.087041e-14, 5.076055e-14, 5.070512e-14, 5.058908e-14, 5.061016e-14, 
    5.06954e-14, 5.088848e-14, 5.0823e-14, 5.098805e-14, 5.098433e-14, 
    5.116781e-14, 5.108512e-14, 5.139314e-14, 5.130568e-14, 5.155828e-14, 
    5.149479e-14, 5.155529e-14, 5.153695e-14, 5.155552e-14, 5.146241e-14, 
    5.150231e-14, 5.142036e-14, 5.11006e-14, 5.119464e-14, 5.091392e-14, 
    5.074477e-14, 5.06324e-14, 5.055258e-14, 5.056387e-14, 5.058537e-14, 
    5.06959e-14, 5.079976e-14, 5.087884e-14, 5.093172e-14, 5.098379e-14, 
    5.114119e-14, 5.122451e-14, 5.14108e-14, 5.137723e-14, 5.143411e-14, 
    5.148848e-14, 5.157965e-14, 5.156465e-14, 5.160479e-14, 5.143264e-14, 
    5.154707e-14, 5.13581e-14, 5.140981e-14, 5.099781e-14, 5.084067e-14, 
    5.077371e-14, 5.071517e-14, 5.057254e-14, 5.067105e-14, 5.063222e-14, 
    5.07246e-14, 5.078325e-14, 5.075425e-14, 5.093316e-14, 5.086363e-14, 
    5.122944e-14, 5.1072e-14, 5.148214e-14, 5.138413e-14, 5.150562e-14, 
    5.144365e-14, 5.154981e-14, 5.145427e-14, 5.161974e-14, 5.165573e-14, 
    5.163114e-14, 5.172563e-14, 5.144897e-14, 5.155527e-14, 5.075343e-14, 
    5.075816e-14, 5.07802e-14, 5.068327e-14, 5.067735e-14, 5.058849e-14, 
    5.066757e-14, 5.070122e-14, 5.078666e-14, 5.083714e-14, 5.088512e-14, 
    5.099056e-14, 5.110819e-14, 5.127253e-14, 5.139048e-14, 5.146948e-14, 
    5.142105e-14, 5.14638e-14, 5.141601e-14, 5.13936e-14, 5.164224e-14, 
    5.150268e-14, 5.171204e-14, 5.170047e-14, 5.160574e-14, 5.170177e-14, 
    5.076148e-14, 5.073426e-14, 5.063968e-14, 5.071371e-14, 5.057882e-14, 
    5.065432e-14, 5.069771e-14, 5.086505e-14, 5.090182e-14, 5.093587e-14, 
    5.100312e-14, 5.108935e-14, 5.124047e-14, 5.137183e-14, 5.149164e-14, 
    5.148287e-14, 5.148596e-14, 5.15127e-14, 5.144644e-14, 5.152357e-14, 
    5.15365e-14, 5.150268e-14, 5.169892e-14, 5.164289e-14, 5.170022e-14, 
    5.166375e-14, 5.074312e-14, 5.078892e-14, 5.076417e-14, 5.081069e-14, 
    5.077791e-14, 5.09236e-14, 5.096725e-14, 5.117132e-14, 5.108764e-14, 
    5.122083e-14, 5.110119e-14, 5.112239e-14, 5.122512e-14, 5.110767e-14, 
    5.136457e-14, 5.11904e-14, 5.151374e-14, 5.133997e-14, 5.152461e-14, 
    5.149113e-14, 5.154658e-14, 5.159621e-14, 5.165864e-14, 5.17737e-14, 
    5.174707e-14, 5.184326e-14, 5.085717e-14, 5.091651e-14, 5.091131e-14, 
    5.09734e-14, 5.101929e-14, 5.111874e-14, 5.127804e-14, 5.121817e-14, 
    5.132809e-14, 5.135014e-14, 5.118314e-14, 5.128568e-14, 5.095623e-14, 
    5.100949e-14, 5.09778e-14, 5.086184e-14, 5.123193e-14, 5.104212e-14, 
    5.139242e-14, 5.128977e-14, 5.158913e-14, 5.144032e-14, 5.173241e-14, 
    5.185698e-14, 5.197423e-14, 5.211096e-14, 5.094891e-14, 5.09086e-14, 
    5.098079e-14, 5.108055e-14, 5.117311e-14, 5.129603e-14, 5.130861e-14, 
    5.133162e-14, 5.139121e-14, 5.144128e-14, 5.133886e-14, 5.145384e-14, 
    5.102179e-14, 5.124841e-14, 5.089334e-14, 5.100033e-14, 5.107468e-14, 
    5.10421e-14, 5.121133e-14, 5.125118e-14, 5.141295e-14, 5.132936e-14, 
    5.182623e-14, 5.160665e-14, 5.221505e-14, 5.204533e-14, 5.089451e-14, 
    5.094879e-14, 5.113746e-14, 5.104773e-14, 5.130424e-14, 5.136729e-14, 
    5.141855e-14, 5.148399e-14, 5.149107e-14, 5.152983e-14, 5.14663e-14, 
    5.152733e-14, 5.129629e-14, 5.13996e-14, 5.111594e-14, 5.118502e-14, 
    5.115325e-14, 5.111838e-14, 5.122598e-14, 5.134047e-14, 5.134296e-14, 
    5.137964e-14, 5.148286e-14, 5.130528e-14, 5.185446e-14, 5.151552e-14, 
    5.100794e-14, 5.111231e-14, 5.112726e-14, 5.108684e-14, 5.136097e-14, 
    5.126171e-14, 5.152889e-14, 5.145675e-14, 5.157494e-14, 5.151622e-14, 
    5.150757e-14, 5.143211e-14, 5.13851e-14, 5.126625e-14, 5.116947e-14, 
    5.109271e-14, 5.111056e-14, 5.119488e-14, 5.134748e-14, 5.149169e-14, 
    5.146011e-14, 5.156596e-14, 5.128566e-14, 5.140325e-14, 5.13578e-14, 
    5.147628e-14, 5.121657e-14, 5.143764e-14, 5.115998e-14, 5.118436e-14, 
    5.125974e-14, 5.14112e-14, 5.144474e-14, 5.148047e-14, 5.145843e-14, 
    5.135136e-14, 5.133383e-14, 5.125791e-14, 5.123692e-14, 5.117906e-14, 
    5.113111e-14, 5.11749e-14, 5.122088e-14, 5.135142e-14, 5.146892e-14, 
    5.15969e-14, 5.162822e-14, 5.177745e-14, 5.165593e-14, 5.185633e-14, 
    5.168589e-14, 5.198083e-14, 5.14505e-14, 5.168095e-14, 5.126318e-14, 
    5.130827e-14, 5.138973e-14, 5.157645e-14, 5.147573e-14, 5.159354e-14, 
    5.133314e-14, 5.119777e-14, 5.116277e-14, 5.109737e-14, 5.116427e-14, 
    5.115883e-14, 5.122281e-14, 5.120226e-14, 5.135575e-14, 5.127333e-14, 
    5.150735e-14, 5.159262e-14, 5.183317e-14, 5.198036e-14, 5.213007e-14, 
    5.219608e-14, 5.221617e-14, 5.222456e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.443775e-15, -7.436983e-15, -7.438304e-15, -7.432832e-15, -7.435868e-15, 
    -7.432286e-15, -7.442398e-15, -7.436712e-15, -7.440342e-15, 
    -7.443165e-15, -7.422236e-15, -7.432589e-15, -7.411532e-15, 
    -7.418107e-15, -7.401614e-15, -7.41255e-15, -7.399413e-15, -7.401933e-15, 
    -7.394364e-15, -7.396531e-15, -7.386857e-15, -7.393364e-15, 
    -7.381857e-15, -7.388412e-15, -7.387384e-15, -7.393578e-15, 
    -7.430507e-15, -7.423522e-15, -7.43092e-15, -7.429923e-15, -7.430371e-15, 
    -7.435803e-15, -7.438542e-15, -7.444297e-15, -7.443252e-15, 
    -7.439027e-15, -7.429475e-15, -7.432717e-15, -7.424561e-15, 
    -7.424745e-15, -7.415684e-15, -7.419766e-15, -7.404574e-15, 
    -7.408887e-15, -7.396441e-15, -7.399566e-15, -7.396586e-15, -7.39749e-15, 
    -7.396575e-15, -7.40116e-15, -7.399194e-15, -7.403233e-15, -7.419001e-15, 
    -7.414358e-15, -7.428219e-15, -7.436576e-15, -7.442148e-15, 
    -7.446106e-15, -7.445546e-15, -7.444478e-15, -7.439002e-15, 
    -7.433866e-15, -7.429956e-15, -7.427345e-15, -7.424772e-15, 
    -7.416986e-15, -7.412881e-15, -7.4037e-15, -7.405359e-15, -7.402552e-15, 
    -7.399877e-15, -7.395386e-15, -7.396126e-15, -7.394148e-15, 
    -7.402628e-15, -7.396989e-15, -7.406304e-15, -7.403753e-15, 
    -7.424059e-15, -7.431843e-15, -7.435145e-15, -7.438049e-15, 
    -7.445116e-15, -7.440233e-15, -7.442156e-15, -7.437585e-15, 
    -7.434683e-15, -7.436118e-15, -7.427273e-15, -7.430707e-15, 
    -7.412638e-15, -7.42041e-15, -7.400189e-15, -7.405019e-15, -7.399034e-15, 
    -7.402087e-15, -7.396855e-15, -7.401564e-15, -7.393413e-15, 
    -7.391638e-15, -7.39285e-15, -7.388202e-15, -7.401825e-15, -7.396586e-15, 
    -7.436158e-15, -7.435924e-15, -7.434834e-15, -7.439628e-15, 
    -7.439922e-15, -7.444325e-15, -7.440408e-15, -7.43874e-15, -7.434516e-15, 
    -7.432017e-15, -7.429644e-15, -7.424435e-15, -7.418624e-15, 
    -7.410517e-15, -7.404705e-15, -7.400814e-15, -7.403201e-15, 
    -7.401094e-15, -7.403449e-15, -7.404554e-15, -7.392302e-15, 
    -7.399175e-15, -7.38887e-15, -7.38944e-15, -7.3941e-15, -7.389376e-15, 
    -7.435759e-15, -7.437108e-15, -7.441788e-15, -7.438125e-15, 
    -7.444806e-15, -7.441062e-15, -7.438911e-15, -7.430633e-15, -7.42882e-15, 
    -7.427137e-15, -7.423816e-15, -7.419557e-15, -7.412098e-15, 
    -7.405623e-15, -7.399722e-15, -7.400155e-15, -7.400003e-15, 
    -7.398684e-15, -7.401948e-15, -7.398148e-15, -7.39751e-15, -7.399178e-15, 
    -7.389516e-15, -7.392274e-15, -7.389452e-15, -7.391248e-15, -7.43667e-15, 
    -7.434402e-15, -7.435627e-15, -7.433324e-15, -7.434945e-15, 
    -7.427739e-15, -7.425581e-15, -7.415505e-15, -7.41964e-15, -7.413065e-15, 
    -7.418973e-15, -7.417925e-15, -7.412844e-15, -7.418654e-15, 
    -7.405977e-15, -7.414561e-15, -7.398633e-15, -7.407184e-15, 
    -7.398098e-15, -7.399748e-15, -7.397017e-15, -7.394571e-15, 
    -7.391498e-15, -7.385833e-15, -7.387145e-15, -7.382413e-15, 
    -7.431027e-15, -7.42809e-15, -7.428352e-15, -7.425284e-15, -7.423016e-15, 
    -7.418108e-15, -7.410247e-15, -7.413201e-15, -7.407783e-15, 
    -7.406694e-15, -7.41493e-15, -7.409869e-15, -7.42613e-15, -7.423495e-15, 
    -7.425065e-15, -7.430794e-15, -7.412517e-15, -7.421884e-15, 
    -7.404609e-15, -7.40967e-15, -7.39492e-15, -7.402245e-15, -7.387866e-15, 
    -7.381729e-15, -7.375974e-15, -7.369244e-15, -7.426494e-15, 
    -7.428486e-15, -7.424921e-15, -7.419987e-15, -7.415423e-15, 
    -7.409361e-15, -7.408742e-15, -7.407607e-15, -7.404671e-15, 
    -7.402203e-15, -7.407246e-15, -7.401585e-15, -7.422878e-15, 
    -7.411707e-15, -7.429237e-15, -7.423946e-15, -7.420278e-15, -7.42189e-15, 
    -7.41354e-15, -7.411575e-15, -7.403596e-15, -7.40772e-15, -7.38324e-15, 
    -7.39405e-15, -7.364138e-15, -7.372472e-15, -7.429182e-15, -7.426501e-15, 
    -7.41718e-15, -7.421612e-15, -7.408957e-15, -7.405848e-15, -7.403325e-15, 
    -7.400097e-15, -7.39975e-15, -7.397839e-15, -7.400971e-15, -7.397965e-15, 
    -7.409348e-15, -7.404257e-15, -7.418247e-15, -7.414835e-15, 
    -7.416405e-15, -7.418127e-15, -7.412816e-15, -7.407165e-15, 
    -7.407049e-15, -7.405238e-15, -7.40013e-15, -7.408907e-15, -7.381838e-15, 
    -7.398524e-15, -7.423579e-15, -7.418417e-15, -7.417686e-15, 
    -7.419683e-15, -7.40616e-15, -7.411054e-15, -7.397887e-15, -7.401442e-15, 
    -7.39562e-15, -7.398511e-15, -7.398937e-15, -7.402655e-15, -7.40497e-15, 
    -7.410828e-15, -7.415602e-15, -7.419394e-15, -7.418512e-15, 
    -7.414347e-15, -7.406821e-15, -7.399717e-15, -7.401271e-15, 
    -7.396062e-15, -7.409874e-15, -7.404073e-15, -7.406313e-15, 
    -7.400478e-15, -7.413279e-15, -7.402362e-15, -7.416073e-15, -7.41487e-15, 
    -7.411151e-15, -7.403678e-15, -7.402033e-15, -7.400269e-15, 
    -7.401359e-15, -7.406631e-15, -7.407497e-15, -7.411243e-15, 
    -7.412274e-15, -7.415132e-15, -7.417498e-15, -7.415336e-15, 
    -7.413065e-15, -7.406631e-15, -7.400839e-15, -7.394536e-15, 
    -7.392996e-15, -7.385637e-15, -7.39162e-15, -7.381745e-15, -7.39013e-15, 
    -7.375631e-15, -7.401736e-15, -7.390386e-15, -7.410983e-15, -7.40876e-15, 
    -7.404737e-15, -7.395536e-15, -7.400506e-15, -7.394697e-15, 
    -7.407532e-15, -7.414201e-15, -7.415935e-15, -7.419162e-15, 
    -7.415862e-15, -7.41613e-15, -7.412973e-15, -7.413988e-15, -7.406417e-15, 
    -7.410483e-15, -7.398946e-15, -7.394744e-15, -7.382907e-15, 
    -7.375666e-15, -7.368315e-15, -7.365073e-15, -7.364087e-15, -7.363674e-15 ;

 CH4_SURF_DIFF_UNSAT =
  4.819795e-14, 4.768278e-14, 4.778307e-14, 4.736664e-14, 4.75978e-14, 
    4.732492e-14, 4.809367e-14, 4.766227e-14, 4.793781e-14, 4.815169e-14, 
    4.655558e-14, 4.734805e-14, 4.572907e-14, 4.623714e-14, 4.495829e-14, 
    4.580818e-14, 4.478647e-14, 4.498296e-14, 4.43912e-14, 4.456092e-14, 
    4.380184e-14, 4.431282e-14, 4.340732e-14, 4.392404e-14, 4.384326e-14, 
    4.432964e-14, 4.718894e-14, 4.665441e-14, 4.722054e-14, 4.714443e-14, 
    4.71786e-14, 4.7593e-14, 4.78014e-14, 4.823732e-14, 4.815828e-14, 
    4.78381e-14, 4.71102e-14, 4.735768e-14, 4.673347e-14, 4.674759e-14, 
    4.60501e-14, 4.636491e-14, 4.518864e-14, 4.552374e-14, 4.455384e-14, 
    4.479822e-14, 4.456531e-14, 4.463598e-14, 4.456439e-14, 4.492267e-14, 
    4.476925e-14, 4.508424e-14, 4.630598e-14, 4.594773e-14, 4.701406e-14, 
    4.765205e-14, 4.807475e-14, 4.837402e-14, 4.833174e-14, 4.82511e-14, 
    4.783622e-14, 4.744533e-14, 4.714683e-14, 4.694685e-14, 4.674962e-14, 
    4.615105e-14, 4.583364e-14, 4.512077e-14, 4.524969e-14, 4.503129e-14, 
    4.482251e-14, 4.447138e-14, 4.452923e-14, 4.437435e-14, 4.503711e-14, 
    4.459687e-14, 4.532307e-14, 4.512472e-14, 4.669567e-14, 4.729096e-14, 
    4.754314e-14, 4.776378e-14, 4.829922e-14, 4.792962e-14, 4.807541e-14, 
    4.772843e-14, 4.750756e-14, 4.761685e-14, 4.694138e-14, 4.720429e-14, 
    4.581481e-14, 4.641461e-14, 4.484688e-14, 4.522324e-14, 4.475657e-14, 
    4.499486e-14, 4.458635e-14, 4.495405e-14, 4.43167e-14, 4.41776e-14, 
    4.427266e-14, 4.390735e-14, 4.49744e-14, 4.456528e-14, 4.76199e-14, 
    4.760208e-14, 4.751906e-14, 4.788367e-14, 4.790596e-14, 4.823947e-14, 
    4.794277e-14, 4.781625e-14, 4.749477e-14, 4.730429e-14, 4.712304e-14, 
    4.672389e-14, 4.6277e-14, 4.565034e-14, 4.519887e-14, 4.489561e-14, 
    4.508164e-14, 4.491741e-14, 4.510098e-14, 4.518697e-14, 4.422971e-14, 
    4.47678e-14, 4.395994e-14, 4.400474e-14, 4.437065e-14, 4.399969e-14, 
    4.758957e-14, 4.769209e-14, 4.804749e-14, 4.776942e-14, 4.827576e-14, 
    4.799248e-14, 4.782937e-14, 4.719873e-14, 4.705995e-14, 4.693105e-14, 
    4.667631e-14, 4.634881e-14, 4.577284e-14, 4.527029e-14, 4.481037e-14, 
    4.484412e-14, 4.483223e-14, 4.472932e-14, 4.49841e-14, 4.468746e-14, 
    4.46376e-14, 4.47679e-14, 4.401073e-14, 4.422736e-14, 4.400569e-14, 
    4.414677e-14, 4.765878e-14, 4.748622e-14, 4.757948e-14, 4.740404e-14, 
    4.752763e-14, 4.697733e-14, 4.681201e-14, 4.60365e-14, 4.635525e-14, 
    4.584778e-14, 4.630379e-14, 4.622305e-14, 4.583107e-14, 4.627919e-14, 
    4.529798e-14, 4.596367e-14, 4.472532e-14, 4.5392e-14, 4.468346e-14, 
    4.481237e-14, 4.459892e-14, 4.440751e-14, 4.41665e-14, 4.372092e-14, 
    4.38242e-14, 4.345103e-14, 4.722867e-14, 4.700425e-14, 4.702407e-14, 
    4.678896e-14, 4.661488e-14, 4.623705e-14, 4.562936e-14, 4.585814e-14, 
    4.543798e-14, 4.535351e-14, 4.599176e-14, 4.560008e-14, 4.685392e-14, 
    4.665187e-14, 4.677224e-14, 4.721095e-14, 4.580537e-14, 4.652804e-14, 
    4.519139e-14, 4.558456e-14, 4.443481e-14, 4.500742e-14, 4.388102e-14, 
    4.339734e-14, 4.29413e-14, 4.240674e-14, 4.688169e-14, 4.703433e-14, 
    4.6761e-14, 4.638205e-14, 4.60299e-14, 4.556059e-14, 4.551253e-14, 
    4.542444e-14, 4.519613e-14, 4.500393e-14, 4.539652e-14, 4.495572e-14, 
    4.660487e-14, 4.574252e-14, 4.709194e-14, 4.668658e-14, 4.640444e-14, 
    4.652832e-14, 4.588428e-14, 4.573213e-14, 4.511256e-14, 4.543313e-14, 
    4.351678e-14, 4.436698e-14, 4.199897e-14, 4.266351e-14, 4.708761e-14, 
    4.688224e-14, 4.616563e-14, 4.650696e-14, 4.552924e-14, 4.528776e-14, 
    4.509127e-14, 4.483971e-14, 4.481257e-14, 4.466334e-14, 4.490781e-14, 
    4.467303e-14, 4.555959e-14, 4.516393e-14, 4.624775e-14, 4.598451e-14, 
    4.610568e-14, 4.623845e-14, 4.582836e-14, 4.539033e-14, 4.538106e-14, 
    4.524037e-14, 4.484318e-14, 4.552528e-14, 4.34066e-14, 4.471766e-14, 
    4.665804e-14, 4.626122e-14, 4.620458e-14, 4.635843e-14, 4.531198e-14, 
    4.569182e-14, 4.466699e-14, 4.494454e-14, 4.44896e-14, 4.471579e-14, 
    4.474905e-14, 4.503914e-14, 4.52195e-14, 4.567441e-14, 4.604375e-14, 
    4.633613e-14, 4.62682e-14, 4.594687e-14, 4.536353e-14, 4.481007e-14, 
    4.493143e-14, 4.452421e-14, 4.560031e-14, 4.514978e-14, 4.532401e-14, 
    4.48694e-14, 4.586419e-14, 4.501712e-14, 4.608005e-14, 4.598712e-14, 
    4.569936e-14, 4.511912e-14, 4.499065e-14, 4.485321e-14, 4.493805e-14, 
    4.534871e-14, 4.541595e-14, 4.570638e-14, 4.578644e-14, 4.600736e-14, 
    4.619002e-14, 4.602312e-14, 4.584766e-14, 4.534858e-14, 4.489763e-14, 
    4.440477e-14, 4.4284e-14, 4.370595e-14, 4.417651e-14, 4.339925e-14, 
    4.406008e-14, 4.291485e-14, 4.496805e-14, 4.407966e-14, 4.568628e-14, 
    4.551388e-14, 4.520154e-14, 4.448341e-14, 4.487154e-14, 4.441759e-14, 
    4.541859e-14, 4.593573e-14, 4.60694e-14, 4.631836e-14, 4.606371e-14, 
    4.608444e-14, 4.584045e-14, 4.59189e-14, 4.533199e-14, 4.564748e-14, 
    4.474986e-14, 4.44212e-14, 4.349014e-14, 4.291712e-14, 4.23323e-14, 
    4.207353e-14, 4.199471e-14, 4.196174e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.93195e-23, 1.931952e-23, 1.931949e-23, 1.93195e-23, 1.931947e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931945e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931945e-23, 
    1.931946e-23, 1.931951e-23, 1.93195e-23, 1.931952e-23, 1.931951e-23, 
    1.931951e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931951e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.93195e-23, 1.931949e-23, 1.931951e-23, 
    1.931952e-23, 1.931953e-23, 1.931954e-23, 1.931954e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931951e-23, 1.931952e-23, 
    1.931952e-23, 1.931953e-23, 1.931954e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931952e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931947e-23, 1.931947e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931945e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 
    1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 1.931954e-23, 
    1.931953e-23, 1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.93195e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931948e-23, 1.931951e-23, 
    1.93195e-23, 1.931951e-23, 1.931952e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 
    1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.93195e-23, 1.931949e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931945e-23, 1.931946e-23, 1.931942e-23, 1.931943e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931948e-23, 1.93195e-23, 1.931949e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931944e-23, 1.931947e-23, 
    1.93195e-23, 1.93195e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931949e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931944e-23, 
    1.931946e-23, 1.931944e-23, 1.931947e-23, 1.931946e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 
    1.931948e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931949e-23, 
    1.931947e-23, 1.931946e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975387e-24, 
    1.975386e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975384e-24, 1.975386e-24, 1.975382e-24, 1.975383e-24, 1.97538e-24, 
    1.975382e-24, 1.975379e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 
    1.975377e-24, 1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975377e-24, 
    1.975378e-24, 1.975386e-24, 1.975384e-24, 1.975386e-24, 1.975385e-24, 
    1.975385e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975385e-24, 1.975386e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975383e-24, 1.97538e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 1.975385e-24, 
    1.975387e-24, 1.975388e-24, 1.975389e-24, 1.975389e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 
    1.975383e-24, 1.975382e-24, 1.97538e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 1.97538e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975384e-24, 1.975386e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975387e-24, 1.975385e-24, 1.975386e-24, 
    1.975382e-24, 1.975383e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.975378e-24, 1.975378e-24, 
    1.975378e-24, 1.975377e-24, 1.97538e-24, 1.975379e-24, 1.975387e-24, 
    1.975387e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975388e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975387e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975388e-24, 1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975378e-24, 1.975387e-24, 1.975386e-24, 1.975387e-24, 1.975386e-24, 
    1.975386e-24, 1.975385e-24, 1.975384e-24, 1.975382e-24, 1.975383e-24, 
    1.975382e-24, 1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975383e-24, 
    1.97538e-24, 1.975382e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975376e-24, 
    1.975377e-24, 1.975376e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975384e-24, 1.975383e-24, 1.975381e-24, 1.975382e-24, 
    1.975381e-24, 1.975381e-24, 1.975382e-24, 1.975381e-24, 1.975385e-24, 
    1.975384e-24, 1.975384e-24, 1.975386e-24, 1.975382e-24, 1.975384e-24, 
    1.97538e-24, 1.975381e-24, 1.975378e-24, 1.97538e-24, 1.975377e-24, 
    1.975376e-24, 1.975374e-24, 1.975373e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 
    1.975384e-24, 1.975382e-24, 1.975385e-24, 1.975384e-24, 1.975383e-24, 
    1.975384e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975381e-24, 
    1.975376e-24, 1.975378e-24, 1.975372e-24, 1.975374e-24, 1.975385e-24, 
    1.975385e-24, 1.975383e-24, 1.975384e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 
    1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975376e-24, 1.975379e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975383e-24, 1.97538e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 1.975382e-24, 
    1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.975379e-24, 1.975382e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 
    1.975381e-24, 1.975381e-24, 1.975382e-24, 1.975382e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.975381e-24, 1.975379e-24, 
    1.975378e-24, 1.975378e-24, 1.975376e-24, 1.975378e-24, 1.975376e-24, 
    1.975377e-24, 1.975374e-24, 1.97538e-24, 1.975377e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 
    1.975381e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.975379e-24, 1.975378e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24 ;

 CONC_CH4_SAT =
  3.512651e-08, 3.512537e-08, 3.512561e-08, 3.512466e-08, 3.51252e-08, 
    3.512457e-08, 3.512629e-08, 3.512531e-08, 3.512595e-08, 3.512643e-08, 
    3.512276e-08, 3.512462e-08, 3.512091e-08, 3.512212e-08, 3.511906e-08, 
    3.512107e-08, 3.511866e-08, 3.511916e-08, 3.511772e-08, 3.511814e-08, 
    3.511618e-08, 3.511753e-08, 3.511521e-08, 3.511653e-08, 3.511631e-08, 
    3.511757e-08, 3.512429e-08, 3.512298e-08, 3.512435e-08, 3.512417e-08, 
    3.512426e-08, 3.512518e-08, 3.512561e-08, 3.512662e-08, 3.512644e-08, 
    3.512572e-08, 3.512409e-08, 3.512467e-08, 3.512327e-08, 3.512331e-08, 
    3.512169e-08, 3.512243e-08, 3.511965e-08, 3.512046e-08, 3.511812e-08, 
    3.511872e-08, 3.511814e-08, 3.511832e-08, 3.511814e-08, 3.511901e-08, 
    3.511864e-08, 3.511941e-08, 3.512228e-08, 3.512144e-08, 3.512389e-08, 
    3.512526e-08, 3.512625e-08, 3.512691e-08, 3.512682e-08, 3.512663e-08, 
    3.512571e-08, 3.512486e-08, 3.512421e-08, 3.512375e-08, 3.512331e-08, 
    3.512186e-08, 3.512115e-08, 3.511947e-08, 3.511981e-08, 3.511926e-08, 
    3.511878e-08, 3.511791e-08, 3.511806e-08, 3.511767e-08, 3.51193e-08, 
    3.511821e-08, 3.511999e-08, 3.511951e-08, 3.512307e-08, 3.512452e-08, 
    3.512502e-08, 3.512556e-08, 3.512674e-08, 3.512592e-08, 3.512624e-08, 
    3.51255e-08, 3.5125e-08, 3.512525e-08, 3.512374e-08, 3.512433e-08, 
    3.512111e-08, 3.512252e-08, 3.511883e-08, 3.511974e-08, 3.511862e-08, 
    3.51192e-08, 3.511819e-08, 3.51191e-08, 3.511753e-08, 3.511717e-08, 
    3.511741e-08, 3.511651e-08, 3.511915e-08, 3.511813e-08, 3.512525e-08, 
    3.512521e-08, 3.512503e-08, 3.512582e-08, 3.512587e-08, 3.512661e-08, 
    3.512596e-08, 3.512567e-08, 3.512498e-08, 3.512455e-08, 3.512414e-08, 
    3.512324e-08, 3.51222e-08, 3.512074e-08, 3.511968e-08, 3.511896e-08, 
    3.511941e-08, 3.511901e-08, 3.511946e-08, 3.511967e-08, 3.51173e-08, 
    3.511863e-08, 3.511664e-08, 3.511676e-08, 3.511765e-08, 3.511675e-08, 
    3.512518e-08, 3.512542e-08, 3.512619e-08, 3.512559e-08, 3.51267e-08, 
    3.512606e-08, 3.512569e-08, 3.512429e-08, 3.512401e-08, 3.512371e-08, 
    3.512314e-08, 3.512239e-08, 3.512103e-08, 3.511984e-08, 3.511875e-08, 
    3.511883e-08, 3.511881e-08, 3.511855e-08, 3.511917e-08, 3.511844e-08, 
    3.511831e-08, 3.511864e-08, 3.511677e-08, 3.511731e-08, 3.511676e-08, 
    3.511711e-08, 3.512535e-08, 3.512496e-08, 3.512516e-08, 3.512476e-08, 
    3.512504e-08, 3.512379e-08, 3.51234e-08, 3.512163e-08, 3.51224e-08, 
    3.51212e-08, 3.512229e-08, 3.512209e-08, 3.512111e-08, 3.512224e-08, 
    3.511988e-08, 3.512144e-08, 3.511854e-08, 3.512008e-08, 3.511844e-08, 
    3.511876e-08, 3.511824e-08, 3.511775e-08, 3.511716e-08, 3.511601e-08, 
    3.511629e-08, 3.511534e-08, 3.512438e-08, 3.512386e-08, 3.512393e-08, 
    3.51234e-08, 3.512299e-08, 3.512214e-08, 3.51207e-08, 3.512125e-08, 
    3.512026e-08, 3.512006e-08, 3.512157e-08, 3.512062e-08, 3.512353e-08, 
    3.512304e-08, 3.512335e-08, 3.512433e-08, 3.512109e-08, 3.512276e-08, 
    3.511966e-08, 3.51206e-08, 3.511782e-08, 3.511919e-08, 3.511643e-08, 
    3.511515e-08, 3.511403e-08, 3.511256e-08, 3.51236e-08, 3.512395e-08, 
    3.512334e-08, 3.512243e-08, 3.512165e-08, 3.512054e-08, 3.512044e-08, 
    3.512022e-08, 3.511969e-08, 3.511922e-08, 3.512013e-08, 3.51191e-08, 
    3.512288e-08, 3.512096e-08, 3.512406e-08, 3.512312e-08, 3.51225e-08, 
    3.51228e-08, 3.512132e-08, 3.512096e-08, 3.511946e-08, 3.512025e-08, 
    3.511544e-08, 3.511762e-08, 3.51115e-08, 3.511326e-08, 3.512407e-08, 
    3.512361e-08, 3.512195e-08, 3.512275e-08, 3.512048e-08, 3.511989e-08, 
    3.511943e-08, 3.511881e-08, 3.511875e-08, 3.511838e-08, 3.511899e-08, 
    3.511841e-08, 3.512054e-08, 3.51196e-08, 3.512217e-08, 3.512154e-08, 
    3.512184e-08, 3.512215e-08, 3.512119e-08, 3.512011e-08, 3.512013e-08, 
    3.511977e-08, 3.511868e-08, 3.512047e-08, 3.511509e-08, 3.51184e-08, 
    3.51231e-08, 3.512215e-08, 3.512206e-08, 3.512242e-08, 3.511995e-08, 
    3.512086e-08, 3.511839e-08, 3.511908e-08, 3.511796e-08, 3.511852e-08, 
    3.51186e-08, 3.511931e-08, 3.511973e-08, 3.512081e-08, 3.512168e-08, 
    3.512237e-08, 3.512222e-08, 3.512145e-08, 3.512005e-08, 3.511873e-08, 
    3.511902e-08, 3.511805e-08, 3.512065e-08, 3.511955e-08, 3.511996e-08, 
    3.511889e-08, 3.512126e-08, 3.511913e-08, 3.512178e-08, 3.512156e-08, 
    3.512087e-08, 3.511945e-08, 3.511919e-08, 3.511884e-08, 3.511906e-08, 
    3.512002e-08, 3.51202e-08, 3.51209e-08, 3.512107e-08, 3.512161e-08, 
    3.512204e-08, 3.512164e-08, 3.512121e-08, 3.512004e-08, 3.511894e-08, 
    3.511774e-08, 3.511746e-08, 3.511591e-08, 3.511712e-08, 3.511506e-08, 
    3.511673e-08, 3.511385e-08, 3.511906e-08, 3.511686e-08, 3.512086e-08, 
    3.512045e-08, 3.511966e-08, 3.51179e-08, 3.511889e-08, 3.511774e-08, 
    3.512021e-08, 3.51214e-08, 3.512175e-08, 3.512232e-08, 3.512174e-08, 
    3.512179e-08, 3.512122e-08, 3.512141e-08, 3.512e-08, 3.512076e-08, 
    3.511859e-08, 3.511776e-08, 3.511542e-08, 3.511392e-08, 3.511242e-08, 
    3.511172e-08, 3.511152e-08, 3.511142e-08,
  6.069577e-11, 6.077409e-11, 6.07589e-11, 6.082198e-11, 6.078706e-11, 
    6.082831e-11, 6.071172e-11, 6.077714e-11, 6.073542e-11, 6.070291e-11, 
    6.094412e-11, 6.082481e-11, 6.107431e-11, 6.09925e-11, 6.119989e-11, 
    6.10613e-11, 6.122784e-11, 6.119606e-11, 6.129207e-11, 6.126459e-11, 
    6.138691e-11, 6.130475e-11, 6.145052e-11, 6.136739e-11, 6.138034e-11, 
    6.130201e-11, 6.084899e-11, 6.092923e-11, 6.084419e-11, 6.085565e-11, 
    6.085054e-11, 6.078772e-11, 6.075596e-11, 6.068989e-11, 6.070192e-11, 
    6.075049e-11, 6.08608e-11, 6.082346e-11, 6.091785e-11, 6.091572e-11, 
    6.102197e-11, 6.097333e-11, 6.116261e-11, 6.110806e-11, 6.126574e-11, 
    6.122609e-11, 6.126385e-11, 6.125242e-11, 6.126399e-11, 6.120585e-11, 
    6.123076e-11, 6.117962e-11, 6.098216e-11, 6.103868e-11, 6.087538e-11, 
    6.077853e-11, 6.071457e-11, 6.066905e-11, 6.067549e-11, 6.068772e-11, 
    6.075077e-11, 6.081018e-11, 6.08554e-11, 6.088562e-11, 6.091541e-11, 
    6.100513e-11, 6.105723e-11, 6.117355e-11, 6.115271e-11, 6.118812e-11, 
    6.122215e-11, 6.127904e-11, 6.12697e-11, 6.129473e-11, 6.11873e-11, 
    6.125866e-11, 6.114081e-11, 6.117304e-11, 6.092297e-11, 6.083356e-11, 
    6.079508e-11, 6.076181e-11, 6.068042e-11, 6.07366e-11, 6.071444e-11, 
    6.076726e-11, 6.080075e-11, 6.078421e-11, 6.088645e-11, 6.084669e-11, 
    6.106032e-11, 6.096576e-11, 6.121818e-11, 6.1157e-11, 6.123286e-11, 
    6.119419e-11, 6.126039e-11, 6.120081e-11, 6.130408e-11, 6.132649e-11, 
    6.131116e-11, 6.137019e-11, 6.119749e-11, 6.126379e-11, 6.078372e-11, 
    6.078641e-11, 6.079903e-11, 6.074357e-11, 6.07402e-11, 6.068954e-11, 
    6.073467e-11, 6.075385e-11, 6.080273e-11, 6.083154e-11, 6.085896e-11, 
    6.091923e-11, 6.098643e-11, 6.108726e-11, 6.116097e-11, 6.121031e-11, 
    6.118009e-11, 6.120676e-11, 6.117692e-11, 6.116296e-11, 6.131805e-11, 
    6.123095e-11, 6.136171e-11, 6.13545e-11, 6.12953e-11, 6.135531e-11, 
    6.078831e-11, 6.07728e-11, 6.071873e-11, 6.076104e-11, 6.068403e-11, 
    6.072707e-11, 6.075178e-11, 6.08474e-11, 6.086853e-11, 6.088796e-11, 
    6.092644e-11, 6.097575e-11, 6.106728e-11, 6.114927e-11, 6.122415e-11, 
    6.121868e-11, 6.12206e-11, 6.123726e-11, 6.119591e-11, 6.124405e-11, 
    6.125207e-11, 6.123101e-11, 6.135353e-11, 6.131855e-11, 6.135435e-11, 
    6.133159e-11, 6.077785e-11, 6.080399e-11, 6.078986e-11, 6.08164e-11, 
    6.079766e-11, 6.088084e-11, 6.090577e-11, 6.102405e-11, 6.097475e-11, 
    6.1055e-11, 6.098253e-11, 6.099462e-11, 6.105747e-11, 6.098626e-11, 
    6.114464e-11, 6.103589e-11, 6.12379e-11, 6.112919e-11, 6.12447e-11, 
    6.122382e-11, 6.125844e-11, 6.128938e-11, 6.132837e-11, 6.140012e-11, 
    6.138354e-11, 6.144359e-11, 6.0843e-11, 6.087685e-11, 6.087397e-11, 
    6.090945e-11, 6.093566e-11, 6.099259e-11, 6.109076e-11, 6.105345e-11, 
    6.112206e-11, 6.113579e-11, 6.10316e-11, 6.109548e-11, 6.089957e-11, 
    6.092993e-11, 6.091193e-11, 6.084561e-11, 6.10619e-11, 6.094861e-11, 
    6.116216e-11, 6.10981e-11, 6.128495e-11, 6.119197e-11, 6.137438e-11, 
    6.145195e-11, 6.152539e-11, 6.161053e-11, 6.089543e-11, 6.087242e-11, 
    6.09137e-11, 6.09706e-11, 6.102529e-11, 6.110199e-11, 6.110989e-11, 
    6.112422e-11, 6.116146e-11, 6.11927e-11, 6.112865e-11, 6.120054e-11, 
    6.093677e-11, 6.107222e-11, 6.086363e-11, 6.092468e-11, 6.096729e-11, 
    6.09487e-11, 6.104921e-11, 6.107406e-11, 6.117492e-11, 6.112286e-11, 
    6.143272e-11, 6.129575e-11, 6.167565e-11, 6.156961e-11, 6.086436e-11, 
    6.089539e-11, 6.10032e-11, 6.095194e-11, 6.110717e-11, 6.114648e-11, 
    6.117853e-11, 6.121929e-11, 6.122378e-11, 6.124793e-11, 6.120833e-11, 
    6.124641e-11, 6.110215e-11, 6.116666e-11, 6.099101e-11, 6.103273e-11, 
    6.101296e-11, 6.099241e-11, 6.105833e-11, 6.112963e-11, 6.113132e-11, 
    6.115414e-11, 6.121811e-11, 6.110781e-11, 6.145006e-11, 6.123857e-11, 
    6.092922e-11, 6.098874e-11, 6.099744e-11, 6.097435e-11, 6.114254e-11, 
    6.108059e-11, 6.124737e-11, 6.120236e-11, 6.127614e-11, 6.123946e-11, 
    6.123407e-11, 6.118698e-11, 6.115761e-11, 6.108339e-11, 6.102301e-11, 
    6.097772e-11, 6.098793e-11, 6.103885e-11, 6.113403e-11, 6.12241e-11, 
    6.120435e-11, 6.127054e-11, 6.109556e-11, 6.116888e-11, 6.11405e-11, 
    6.121453e-11, 6.105241e-11, 6.118997e-11, 6.101716e-11, 6.103236e-11, 
    6.107936e-11, 6.117374e-11, 6.119486e-11, 6.12171e-11, 6.120342e-11, 
    6.113648e-11, 6.112558e-11, 6.107825e-11, 6.10651e-11, 6.102906e-11, 
    6.099968e-11, 6.102644e-11, 6.105506e-11, 6.113657e-11, 6.120988e-11, 
    6.128979e-11, 6.13094e-11, 6.140222e-11, 6.132643e-11, 6.145121e-11, 
    6.134478e-11, 6.152909e-11, 6.119818e-11, 6.134199e-11, 6.108155e-11, 
    6.110969e-11, 6.116038e-11, 6.127689e-11, 6.121419e-11, 6.128759e-11, 
    6.112517e-11, 6.104058e-11, 6.101889e-11, 6.098035e-11, 6.101982e-11, 
    6.101643e-11, 6.105637e-11, 6.104355e-11, 6.113928e-11, 6.108788e-11, 
    6.123388e-11, 6.128705e-11, 6.143724e-11, 6.152905e-11, 6.162267e-11, 
    6.166387e-11, 6.167642e-11, 6.168165e-11,
  2.81559e-14, 2.822542e-14, 2.821193e-14, 2.826799e-14, 2.823693e-14, 
    2.827361e-14, 2.817004e-14, 2.822814e-14, 2.819107e-14, 2.816223e-14, 
    2.837678e-14, 2.82705e-14, 2.84913e-14, 2.841987e-14, 2.860066e-14, 
    2.848e-14, 2.862503e-14, 2.859731e-14, 2.86811e-14, 2.86571e-14, 
    2.876408e-14, 2.869218e-14, 2.88198e-14, 2.874698e-14, 2.875832e-14, 
    2.868979e-14, 2.829199e-14, 2.83635e-14, 2.828773e-14, 2.829793e-14, 
    2.829338e-14, 2.823753e-14, 2.820932e-14, 2.815068e-14, 2.816134e-14, 
    2.820446e-14, 2.830252e-14, 2.826929e-14, 2.83533e-14, 2.83514e-14, 
    2.844579e-14, 2.840276e-14, 2.856815e-14, 2.852064e-14, 2.86581e-14, 
    2.862349e-14, 2.865645e-14, 2.864647e-14, 2.865658e-14, 2.860584e-14, 
    2.862757e-14, 2.858297e-14, 2.841065e-14, 2.846031e-14, 2.831549e-14, 
    2.822939e-14, 2.817257e-14, 2.81322e-14, 2.81379e-14, 2.814875e-14, 
    2.820471e-14, 2.825748e-14, 2.82977e-14, 2.83246e-14, 2.835113e-14, 
    2.843119e-14, 2.847644e-14, 2.85777e-14, 2.855952e-14, 2.859039e-14, 
    2.862005e-14, 2.866972e-14, 2.866156e-14, 2.868343e-14, 2.858966e-14, 
    2.865193e-14, 2.854914e-14, 2.857723e-14, 2.835793e-14, 2.827827e-14, 
    2.82441e-14, 2.821451e-14, 2.814228e-14, 2.819212e-14, 2.817246e-14, 
    2.821934e-14, 2.824909e-14, 2.823439e-14, 2.832533e-14, 2.828994e-14, 
    2.847912e-14, 2.839602e-14, 2.861659e-14, 2.856326e-14, 2.86294e-14, 
    2.859566e-14, 2.865344e-14, 2.860144e-14, 2.86916e-14, 2.871119e-14, 
    2.869779e-14, 2.874942e-14, 2.859855e-14, 2.865641e-14, 2.823396e-14, 
    2.823636e-14, 2.824756e-14, 2.819831e-14, 2.819533e-14, 2.815036e-14, 
    2.819041e-14, 2.820744e-14, 2.825085e-14, 2.827647e-14, 2.830086e-14, 
    2.835454e-14, 2.841447e-14, 2.850255e-14, 2.856671e-14, 2.860972e-14, 
    2.858337e-14, 2.860663e-14, 2.858062e-14, 2.856844e-14, 2.870382e-14, 
    2.862775e-14, 2.874199e-14, 2.873568e-14, 2.868393e-14, 2.87364e-14, 
    2.823805e-14, 2.822425e-14, 2.817626e-14, 2.821382e-14, 2.814547e-14, 
    2.818367e-14, 2.820561e-14, 2.829059e-14, 2.830938e-14, 2.832668e-14, 
    2.836096e-14, 2.840492e-14, 2.848517e-14, 2.855653e-14, 2.86218e-14, 
    2.861702e-14, 2.86187e-14, 2.863324e-14, 2.859717e-14, 2.863917e-14, 
    2.864618e-14, 2.862779e-14, 2.873484e-14, 2.870425e-14, 2.873555e-14, 
    2.871564e-14, 2.822875e-14, 2.825198e-14, 2.823942e-14, 2.826302e-14, 
    2.824636e-14, 2.832036e-14, 2.834256e-14, 2.84476e-14, 2.840403e-14, 
    2.84745e-14, 2.841097e-14, 2.842176e-14, 2.847668e-14, 2.84143e-14, 
    2.855252e-14, 2.845791e-14, 2.863381e-14, 2.853907e-14, 2.863974e-14, 
    2.862151e-14, 2.865173e-14, 2.867875e-14, 2.871283e-14, 2.877563e-14, 
    2.876111e-14, 2.881371e-14, 2.828667e-14, 2.831679e-14, 2.831422e-14, 
    2.834582e-14, 2.836918e-14, 2.841994e-14, 2.850559e-14, 2.847313e-14, 
    2.853282e-14, 2.854478e-14, 2.845415e-14, 2.850971e-14, 2.833702e-14, 
    2.836409e-14, 2.834803e-14, 2.8289e-14, 2.84805e-14, 2.838074e-14, 
    2.856775e-14, 2.851198e-14, 2.867489e-14, 2.859375e-14, 2.875309e-14, 
    2.882108e-14, 2.888548e-14, 2.896034e-14, 2.833333e-14, 2.831284e-14, 
    2.83496e-14, 2.840035e-14, 2.844867e-14, 2.851536e-14, 2.852223e-14, 
    2.853471e-14, 2.856714e-14, 2.859437e-14, 2.853858e-14, 2.860121e-14, 
    2.837021e-14, 2.848947e-14, 2.830503e-14, 2.835941e-14, 2.839739e-14, 
    2.83808e-14, 2.846944e-14, 2.849105e-14, 2.857888e-14, 2.853351e-14, 
    2.880422e-14, 2.868434e-14, 2.901765e-14, 2.892435e-14, 2.830567e-14, 
    2.833329e-14, 2.842943e-14, 2.838368e-14, 2.851986e-14, 2.85541e-14, 
    2.858201e-14, 2.861757e-14, 2.862147e-14, 2.864256e-14, 2.8608e-14, 
    2.864123e-14, 2.85155e-14, 2.857167e-14, 2.841853e-14, 2.845513e-14, 
    2.843795e-14, 2.841977e-14, 2.847738e-14, 2.853944e-14, 2.854089e-14, 
    2.856078e-14, 2.861661e-14, 2.852043e-14, 2.881946e-14, 2.863445e-14, 
    2.836343e-14, 2.841653e-14, 2.842428e-14, 2.840367e-14, 2.855066e-14, 
    2.849674e-14, 2.864206e-14, 2.860279e-14, 2.866718e-14, 2.863517e-14, 
    2.863045e-14, 2.858938e-14, 2.856379e-14, 2.849918e-14, 2.844669e-14, 
    2.840667e-14, 2.841578e-14, 2.846046e-14, 2.854327e-14, 2.862177e-14, 
    2.860455e-14, 2.866229e-14, 2.850976e-14, 2.857362e-14, 2.854889e-14, 
    2.861341e-14, 2.847224e-14, 2.859205e-14, 2.84416e-14, 2.84548e-14, 
    2.849567e-14, 2.857787e-14, 2.859626e-14, 2.861566e-14, 2.860371e-14, 
    2.854539e-14, 2.85359e-14, 2.84947e-14, 2.848327e-14, 2.845194e-14, 
    2.842628e-14, 2.844966e-14, 2.847455e-14, 2.854547e-14, 2.860936e-14, 
    2.867912e-14, 2.869624e-14, 2.87775e-14, 2.871117e-14, 2.882047e-14, 
    2.872727e-14, 2.888879e-14, 2.859919e-14, 2.872479e-14, 2.849757e-14, 
    2.852205e-14, 2.856621e-14, 2.866786e-14, 2.861311e-14, 2.867721e-14, 
    2.853554e-14, 2.846197e-14, 2.84431e-14, 2.840903e-14, 2.844391e-14, 
    2.844097e-14, 2.847567e-14, 2.846453e-14, 2.854783e-14, 2.850308e-14, 
    2.86303e-14, 2.867673e-14, 2.880815e-14, 2.888871e-14, 2.897099e-14, 
    2.900726e-14, 2.901832e-14, 2.902293e-14,
  3.876818e-18, 3.890717e-18, 3.888014e-18, 3.899247e-18, 3.893021e-18, 
    3.900374e-18, 3.87963e-18, 3.891262e-18, 3.883838e-18, 3.878066e-18, 
    3.921084e-18, 3.899751e-18, 3.943763e-18, 3.929737e-18, 3.965168e-18, 
    3.941554e-18, 3.969944e-18, 3.964508e-18, 3.980938e-18, 3.976228e-18, 
    3.997239e-18, 3.983113e-18, 4.008194e-18, 3.993875e-18, 3.996105e-18, 
    3.982643e-18, 3.904058e-18, 3.918417e-18, 3.903204e-18, 3.90525e-18, 
    3.904336e-18, 3.893142e-18, 3.887495e-18, 3.875821e-18, 3.877888e-18, 
    3.88652e-18, 3.906171e-18, 3.899506e-18, 3.916359e-18, 3.915978e-18, 
    3.934866e-18, 3.926298e-18, 3.958797e-18, 3.949498e-18, 3.976425e-18, 
    3.969639e-18, 3.976102e-18, 3.974145e-18, 3.976128e-18, 3.96618e-18, 
    3.970439e-18, 3.961699e-18, 3.927882e-18, 3.937704e-18, 3.908773e-18, 
    3.891515e-18, 3.880136e-18, 3.872305e-18, 3.87339e-18, 3.875457e-18, 
    3.886571e-18, 3.897139e-18, 3.905202e-18, 3.910598e-18, 3.915923e-18, 
    3.932017e-18, 3.940859e-18, 3.960668e-18, 3.957108e-18, 3.963155e-18, 
    3.968966e-18, 3.978706e-18, 3.977105e-18, 3.981395e-18, 3.963009e-18, 
    3.975216e-18, 3.955076e-18, 3.960576e-18, 3.917299e-18, 3.901307e-18, 
    3.894461e-18, 3.888531e-18, 3.874224e-18, 3.88405e-18, 3.880114e-18, 
    3.889498e-18, 3.895458e-18, 3.892513e-18, 3.910746e-18, 3.903647e-18, 
    3.941383e-18, 3.924944e-18, 3.968288e-18, 3.95784e-18, 3.970797e-18, 
    3.964186e-18, 3.975512e-18, 3.965318e-18, 3.982999e-18, 3.986846e-18, 
    3.984215e-18, 3.994354e-18, 3.964751e-18, 3.976095e-18, 3.892427e-18, 
    3.892906e-18, 3.895151e-18, 3.885289e-18, 3.884691e-18, 3.875762e-18, 
    3.883705e-18, 3.887115e-18, 3.89581e-18, 3.900946e-18, 3.905838e-18, 
    3.91661e-18, 3.928653e-18, 3.945963e-18, 3.958515e-18, 3.96694e-18, 
    3.961778e-18, 3.966335e-18, 3.961238e-18, 3.958854e-18, 3.9854e-18, 
    3.970474e-18, 3.992894e-18, 3.991655e-18, 3.981494e-18, 3.991795e-18, 
    3.893245e-18, 3.890481e-18, 3.880875e-18, 3.888391e-18, 3.874832e-18, 
    3.882356e-18, 3.88675e-18, 3.90378e-18, 3.907546e-18, 3.911017e-18, 
    3.917898e-18, 3.926731e-18, 3.942563e-18, 3.956524e-18, 3.969307e-18, 
    3.968371e-18, 3.9687e-18, 3.971551e-18, 3.964481e-18, 3.972713e-18, 
    3.974088e-18, 3.970481e-18, 3.991488e-18, 3.985481e-18, 3.991628e-18, 
    3.987718e-18, 3.891381e-18, 3.896036e-18, 3.893519e-18, 3.898249e-18, 
    3.894911e-18, 3.909751e-18, 3.914208e-18, 3.935223e-18, 3.926553e-18, 
    3.940478e-18, 3.927947e-18, 3.930117e-18, 3.940906e-18, 3.928615e-18, 
    3.955739e-18, 3.937237e-18, 3.971661e-18, 3.953109e-18, 3.972824e-18, 
    3.969251e-18, 3.975175e-18, 3.980477e-18, 3.987167e-18, 3.999507e-18, 
    3.996651e-18, 4.006995e-18, 3.90299e-18, 3.909035e-18, 3.908516e-18, 
    3.914858e-18, 3.91955e-18, 3.92975e-18, 3.946556e-18, 3.940209e-18, 
    3.951881e-18, 3.954222e-18, 3.936499e-18, 3.947362e-18, 3.913095e-18, 
    3.91853e-18, 3.915303e-18, 3.903459e-18, 3.941651e-18, 3.921874e-18, 
    3.958721e-18, 3.947804e-18, 3.979719e-18, 3.963813e-18, 3.995076e-18, 
    4.008447e-18, 4.021123e-18, 4.035887e-18, 3.912351e-18, 3.908239e-18, 
    3.915617e-18, 3.925814e-18, 3.935429e-18, 3.948467e-18, 3.94981e-18, 
    3.952252e-18, 3.958599e-18, 3.963933e-18, 3.953011e-18, 3.965272e-18, 
    3.919764e-18, 3.943404e-18, 3.906673e-18, 3.91759e-18, 3.925219e-18, 
    3.921885e-18, 3.939487e-18, 3.943711e-18, 3.960901e-18, 3.952017e-18, 
    4.005132e-18, 3.981578e-18, 4.047197e-18, 4.028788e-18, 3.9068e-18, 
    3.912344e-18, 3.931661e-18, 3.922464e-18, 3.949346e-18, 3.956046e-18, 
    3.961511e-18, 3.96848e-18, 3.969243e-18, 3.973378e-18, 3.966602e-18, 
    3.973116e-18, 3.948495e-18, 3.959488e-18, 3.929466e-18, 3.936691e-18, 
    3.933334e-18, 3.929716e-18, 3.941039e-18, 3.953178e-18, 3.953461e-18, 
    3.957355e-18, 3.968299e-18, 3.949457e-18, 4.008136e-18, 3.971795e-18, 
    3.918394e-18, 3.929068e-18, 3.930622e-18, 3.926479e-18, 3.955373e-18, 
    3.944824e-18, 3.973281e-18, 3.965582e-18, 3.978206e-18, 3.971928e-18, 
    3.971004e-18, 3.962955e-18, 3.957943e-18, 3.945302e-18, 3.935043e-18, 
    3.927082e-18, 3.928914e-18, 3.937732e-18, 3.953927e-18, 3.969302e-18, 
    3.965928e-18, 3.977247e-18, 3.94737e-18, 3.95987e-18, 3.955028e-18, 
    3.967663e-18, 3.940035e-18, 3.963486e-18, 3.934047e-18, 3.936627e-18, 
    3.944614e-18, 3.960702e-18, 3.964302e-18, 3.968105e-18, 3.965762e-18, 
    3.954343e-18, 3.952484e-18, 3.944426e-18, 3.942191e-18, 3.936067e-18, 
    3.931023e-18, 3.935623e-18, 3.940487e-18, 3.954357e-18, 3.966871e-18, 
    3.980549e-18, 3.98391e-18, 3.999879e-18, 3.986845e-18, 4.008334e-18, 
    3.990013e-18, 4.021783e-18, 3.964881e-18, 3.989521e-18, 3.944986e-18, 
    3.949774e-18, 3.95842e-18, 3.978344e-18, 3.967604e-18, 3.980177e-18, 
    3.952413e-18, 3.938029e-18, 3.934341e-18, 3.927557e-18, 3.934499e-18, 
    3.933924e-18, 3.940704e-18, 3.938526e-18, 3.954819e-18, 3.946063e-18, 
    3.970974e-18, 3.980083e-18, 4.005902e-18, 4.021764e-18, 4.037984e-18, 
    4.045145e-18, 4.047328e-18, 4.048239e-18,
  1.666524e-22, 1.674562e-22, 1.672997e-22, 1.679502e-22, 1.675895e-22, 
    1.680155e-22, 1.668147e-22, 1.674878e-22, 1.670581e-22, 1.667243e-22, 
    1.692169e-22, 1.679794e-22, 1.705393e-22, 1.697187e-22, 1.718049e-22, 
    1.704089e-22, 1.720876e-22, 1.717656e-22, 1.727387e-22, 1.724596e-22, 
    1.737063e-22, 1.728676e-22, 1.743568e-22, 1.735063e-22, 1.736387e-22, 
    1.728398e-22, 1.682288e-22, 1.690621e-22, 1.681793e-22, 1.68298e-22, 
    1.682449e-22, 1.675966e-22, 1.672699e-22, 1.665952e-22, 1.66714e-22, 
    1.672134e-22, 1.683514e-22, 1.679651e-22, 1.68942e-22, 1.689199e-22, 
    1.700143e-22, 1.695189e-22, 1.714277e-22, 1.708778e-22, 1.724712e-22, 
    1.720693e-22, 1.724522e-22, 1.723361e-22, 1.724537e-22, 1.718646e-22, 
    1.721167e-22, 1.715993e-22, 1.69611e-22, 1.701813e-22, 1.685022e-22, 
    1.675027e-22, 1.66844e-22, 1.663937e-22, 1.664559e-22, 1.665744e-22, 
    1.672163e-22, 1.67828e-22, 1.682951e-22, 1.686079e-22, 1.689168e-22, 
    1.698516e-22, 1.703677e-22, 1.715385e-22, 1.713277e-22, 1.716856e-22, 
    1.720294e-22, 1.726065e-22, 1.725115e-22, 1.727659e-22, 1.716769e-22, 
    1.723998e-22, 1.712075e-22, 1.715328e-22, 1.689973e-22, 1.680694e-22, 
    1.676732e-22, 1.673297e-22, 1.665037e-22, 1.670704e-22, 1.668428e-22, 
    1.673855e-22, 1.677306e-22, 1.6756e-22, 1.686165e-22, 1.68205e-22, 
    1.703987e-22, 1.694404e-22, 1.719893e-22, 1.71371e-22, 1.721379e-22, 
    1.717464e-22, 1.724172e-22, 1.718134e-22, 1.728609e-22, 1.730892e-22, 
    1.729331e-22, 1.735345e-22, 1.717799e-22, 1.724518e-22, 1.675551e-22, 
    1.675829e-22, 1.677128e-22, 1.671422e-22, 1.671075e-22, 1.665918e-22, 
    1.670504e-22, 1.672477e-22, 1.677509e-22, 1.680485e-22, 1.68332e-22, 
    1.689566e-22, 1.696558e-22, 1.706691e-22, 1.71411e-22, 1.719095e-22, 
    1.716039e-22, 1.718736e-22, 1.71572e-22, 1.714309e-22, 1.730034e-22, 
    1.721189e-22, 1.734479e-22, 1.733743e-22, 1.727718e-22, 1.733826e-22, 
    1.676024e-22, 1.674424e-22, 1.668867e-22, 1.673215e-22, 1.665385e-22, 
    1.669724e-22, 1.672267e-22, 1.682128e-22, 1.684309e-22, 1.686323e-22, 
    1.690313e-22, 1.695441e-22, 1.704682e-22, 1.712933e-22, 1.720496e-22, 
    1.719942e-22, 1.720136e-22, 1.721825e-22, 1.717639e-22, 1.722513e-22, 
    1.723329e-22, 1.721192e-22, 1.733645e-22, 1.730081e-22, 1.733728e-22, 
    1.731407e-22, 1.674945e-22, 1.677641e-22, 1.676183e-22, 1.678923e-22, 
    1.67699e-22, 1.68559e-22, 1.688175e-22, 1.70035e-22, 1.695338e-22, 
    1.703451e-22, 1.696147e-22, 1.697408e-22, 1.703708e-22, 1.696534e-22, 
    1.71247e-22, 1.70154e-22, 1.721891e-22, 1.710917e-22, 1.722579e-22, 
    1.720463e-22, 1.723972e-22, 1.727115e-22, 1.731081e-22, 1.738407e-22, 
    1.73671e-22, 1.742855e-22, 1.681669e-22, 1.685174e-22, 1.684871e-22, 
    1.68855e-22, 1.691272e-22, 1.697194e-22, 1.70704e-22, 1.70329e-22, 
    1.710186e-22, 1.711571e-22, 1.7011e-22, 1.707517e-22, 1.687528e-22, 
    1.690683e-22, 1.688809e-22, 1.681941e-22, 1.704144e-22, 1.692623e-22, 
    1.714231e-22, 1.707777e-22, 1.726665e-22, 1.717246e-22, 1.735775e-22, 
    1.743721e-22, 1.751256e-22, 1.760052e-22, 1.687096e-22, 1.684711e-22, 
    1.688989e-22, 1.69491e-22, 1.700469e-22, 1.708169e-22, 1.708962e-22, 
    1.710406e-22, 1.714158e-22, 1.717315e-22, 1.710856e-22, 1.718107e-22, 
    1.691402e-22, 1.705179e-22, 1.683804e-22, 1.690138e-22, 1.694564e-22, 
    1.692628e-22, 1.702864e-22, 1.705358e-22, 1.715522e-22, 1.710266e-22, 
    1.741751e-22, 1.72777e-22, 1.766794e-22, 1.755822e-22, 1.683877e-22, 
    1.687091e-22, 1.698305e-22, 1.692963e-22, 1.708688e-22, 1.712649e-22, 
    1.715881e-22, 1.720008e-22, 1.720458e-22, 1.722908e-22, 1.718894e-22, 
    1.722752e-22, 1.708186e-22, 1.714685e-22, 1.697028e-22, 1.701214e-22, 
    1.699265e-22, 1.697174e-22, 1.70378e-22, 1.710956e-22, 1.71112e-22, 
    1.713424e-22, 1.71991e-22, 1.708753e-22, 1.743542e-22, 1.721979e-22, 
    1.690601e-22, 1.696801e-22, 1.697701e-22, 1.695294e-22, 1.712252e-22, 
    1.706016e-22, 1.72285e-22, 1.718291e-22, 1.725768e-22, 1.722049e-22, 
    1.721501e-22, 1.716736e-22, 1.713771e-22, 1.7063e-22, 1.700244e-22, 
    1.695644e-22, 1.696708e-22, 1.701829e-22, 1.711398e-22, 1.720494e-22, 
    1.718497e-22, 1.725199e-22, 1.707521e-22, 1.714912e-22, 1.712049e-22, 
    1.719523e-22, 1.703188e-22, 1.717058e-22, 1.699673e-22, 1.701175e-22, 
    1.705893e-22, 1.715407e-22, 1.717533e-22, 1.719786e-22, 1.718398e-22, 
    1.711644e-22, 1.710544e-22, 1.705781e-22, 1.704462e-22, 1.700845e-22, 
    1.697933e-22, 1.700583e-22, 1.703456e-22, 1.711651e-22, 1.719055e-22, 
    1.727158e-22, 1.729149e-22, 1.738632e-22, 1.730895e-22, 1.74366e-22, 
    1.73278e-22, 1.751656e-22, 1.717881e-22, 1.732483e-22, 1.706111e-22, 
    1.708941e-22, 1.714056e-22, 1.725853e-22, 1.719488e-22, 1.726939e-22, 
    1.710501e-22, 1.702006e-22, 1.699841e-22, 1.69592e-22, 1.699932e-22, 
    1.699602e-22, 1.703582e-22, 1.702296e-22, 1.711924e-22, 1.706748e-22, 
    1.721485e-22, 1.726883e-22, 1.742206e-22, 1.75164e-22, 1.761298e-22, 
    1.765568e-22, 1.76687e-22, 1.767414e-22,
  2.315837e-27, 2.330074e-27, 2.327301e-27, 2.338831e-27, 2.332435e-27, 
    2.339989e-27, 2.318712e-27, 2.330636e-27, 2.323022e-27, 2.317111e-27, 
    2.361327e-27, 2.339349e-27, 2.384825e-27, 2.37024e-27, 2.407394e-27, 
    2.382506e-27, 2.412441e-27, 2.406688e-27, 2.424072e-27, 2.419083e-27, 
    2.441395e-27, 2.426378e-27, 2.453051e-27, 2.437811e-27, 2.440184e-27, 
    2.425881e-27, 2.343771e-27, 2.358576e-27, 2.342893e-27, 2.345e-27, 
    2.344058e-27, 2.332562e-27, 2.326777e-27, 2.314805e-27, 2.316929e-27, 
    2.325773e-27, 2.345948e-27, 2.339092e-27, 2.356431e-27, 2.356039e-27, 
    2.375477e-27, 2.366685e-27, 2.400658e-27, 2.390852e-27, 2.419291e-27, 
    2.412111e-27, 2.418951e-27, 2.416877e-27, 2.418978e-27, 2.408456e-27, 
    2.412958e-27, 2.403721e-27, 2.368323e-27, 2.378449e-27, 2.348623e-27, 
    2.330903e-27, 2.319232e-27, 2.31121e-27, 2.312303e-27, 2.314433e-27, 
    2.325824e-27, 2.336662e-27, 2.344945e-27, 2.350498e-27, 2.355982e-27, 
    2.37261e-27, 2.38177e-27, 2.402638e-27, 2.398874e-27, 2.405263e-27, 
    2.411398e-27, 2.42171e-27, 2.420012e-27, 2.424561e-27, 2.405104e-27, 
    2.418016e-27, 2.396729e-27, 2.402534e-27, 2.357426e-27, 2.340942e-27, 
    2.333924e-27, 2.327832e-27, 2.313162e-27, 2.323241e-27, 2.319211e-27, 
    2.32882e-27, 2.334936e-27, 2.331911e-27, 2.35065e-27, 2.343348e-27, 
    2.382321e-27, 2.365292e-27, 2.410682e-27, 2.399647e-27, 2.413335e-27, 
    2.406345e-27, 2.418328e-27, 2.407541e-27, 2.426259e-27, 2.430345e-27, 
    2.427551e-27, 2.438313e-27, 2.406943e-27, 2.418946e-27, 2.331824e-27, 
    2.332317e-27, 2.334619e-27, 2.324512e-27, 2.323897e-27, 2.314746e-27, 
    2.322885e-27, 2.326381e-27, 2.335295e-27, 2.340572e-27, 2.345601e-27, 
    2.356692e-27, 2.369122e-27, 2.387135e-27, 2.40036e-27, 2.409256e-27, 
    2.403802e-27, 2.408616e-27, 2.403233e-27, 2.400715e-27, 2.42881e-27, 
    2.412997e-27, 2.436763e-27, 2.435445e-27, 2.424667e-27, 2.435594e-27, 
    2.332664e-27, 2.329827e-27, 2.319987e-27, 2.327685e-27, 2.313786e-27, 
    2.321506e-27, 2.32601e-27, 2.34349e-27, 2.347357e-27, 2.350932e-27, 
    2.358018e-27, 2.367133e-27, 2.383557e-27, 2.398262e-27, 2.411758e-27, 
    2.410768e-27, 2.411116e-27, 2.414133e-27, 2.406658e-27, 2.415363e-27, 
    2.416821e-27, 2.413001e-27, 2.435268e-27, 2.428891e-27, 2.435417e-27, 
    2.431264e-27, 2.33075e-27, 2.335529e-27, 2.332945e-27, 2.337803e-27, 
    2.334376e-27, 2.349634e-27, 2.354225e-27, 2.375847e-27, 2.366951e-27, 
    2.381365e-27, 2.368388e-27, 2.370633e-27, 2.381828e-27, 2.369077e-27, 
    2.39744e-27, 2.377966e-27, 2.41425e-27, 2.394673e-27, 2.415481e-27, 
    2.411699e-27, 2.417967e-27, 2.423587e-27, 2.430681e-27, 2.443799e-27, 
    2.440758e-27, 2.451769e-27, 2.342672e-27, 2.348893e-27, 2.348354e-27, 
    2.354886e-27, 2.359724e-27, 2.37025e-27, 2.387756e-27, 2.381076e-27, 
    2.393362e-27, 2.395832e-27, 2.377176e-27, 2.388607e-27, 2.353072e-27, 
    2.358679e-27, 2.355346e-27, 2.343157e-27, 2.382601e-27, 2.362127e-27, 
    2.400578e-27, 2.389069e-27, 2.422784e-27, 2.40596e-27, 2.439084e-27, 
    2.453329e-27, 2.4669e-27, 2.483114e-27, 2.352305e-27, 2.34807e-27, 
    2.355666e-27, 2.366193e-27, 2.376056e-27, 2.389768e-27, 2.39118e-27, 
    2.393755e-27, 2.400445e-27, 2.406078e-27, 2.39456e-27, 2.407493e-27, 
    2.359963e-27, 2.384442e-27, 2.346462e-27, 2.357711e-27, 2.365575e-27, 
    2.362132e-27, 2.380316e-27, 2.384759e-27, 2.402882e-27, 2.393505e-27, 
    2.449799e-27, 2.424762e-27, 2.495549e-27, 2.475314e-27, 2.346589e-27, 
    2.352295e-27, 2.37223e-27, 2.362729e-27, 2.390691e-27, 2.397755e-27, 
    2.403519e-27, 2.410888e-27, 2.411691e-27, 2.416068e-27, 2.408898e-27, 
    2.415788e-27, 2.389797e-27, 2.401386e-27, 2.369955e-27, 2.377381e-27, 
    2.373925e-27, 2.370214e-27, 2.381948e-27, 2.394738e-27, 2.395028e-27, 
    2.399138e-27, 2.410726e-27, 2.390808e-27, 2.453016e-27, 2.41442e-27, 
    2.358529e-27, 2.369555e-27, 2.371152e-27, 2.36687e-27, 2.397046e-27, 
    2.385932e-27, 2.415964e-27, 2.407821e-27, 2.421179e-27, 2.414532e-27, 
    2.413554e-27, 2.405046e-27, 2.399756e-27, 2.386438e-27, 2.375656e-27, 
    2.367493e-27, 2.369385e-27, 2.378477e-27, 2.395526e-27, 2.411757e-27, 
    2.408192e-27, 2.420162e-27, 2.388612e-27, 2.401792e-27, 2.396686e-27, 
    2.410022e-27, 2.380895e-27, 2.405634e-27, 2.374645e-27, 2.377311e-27, 
    2.385712e-27, 2.402678e-27, 2.406468e-27, 2.410492e-27, 2.408011e-27, 
    2.395963e-27, 2.394001e-27, 2.385511e-27, 2.383164e-27, 2.376721e-27, 
    2.371564e-27, 2.376257e-27, 2.381373e-27, 2.395975e-27, 2.409187e-27, 
    2.423665e-27, 2.427224e-27, 2.444209e-27, 2.430354e-27, 2.45323e-27, 
    2.433739e-27, 2.46765e-27, 2.407096e-27, 2.433198e-27, 2.3861e-27, 
    2.391142e-27, 2.400267e-27, 2.421336e-27, 2.409959e-27, 2.423276e-27, 
    2.393925e-27, 2.378793e-27, 2.374943e-27, 2.367984e-27, 2.375103e-27, 
    2.374521e-27, 2.381596e-27, 2.379305e-27, 2.396461e-27, 2.387234e-27, 
    2.413526e-27, 2.423174e-27, 2.450608e-27, 2.467613e-27, 2.485405e-27, 
    2.493285e-27, 2.495688e-27, 2.496693e-27,
  1.031222e-32, 1.039212e-32, 1.037655e-32, 1.044133e-32, 1.040537e-32, 
    1.044784e-32, 1.032836e-32, 1.039529e-32, 1.035253e-32, 1.031938e-32, 
    1.056919e-32, 1.044424e-32, 1.070412e-32, 1.06206e-32, 1.083302e-32, 
    1.06909e-32, 1.086189e-32, 1.082896e-32, 1.092851e-32, 1.089991e-32, 
    1.102798e-32, 1.094173e-32, 1.109501e-32, 1.100737e-32, 1.102101e-32, 
    1.093888e-32, 1.04691e-32, 1.055333e-32, 1.046416e-32, 1.047602e-32, 
    1.047071e-32, 1.040609e-32, 1.037363e-32, 1.030634e-32, 1.031836e-32, 
    1.036798e-32, 1.048135e-32, 1.044278e-32, 1.054089e-32, 1.053863e-32, 
    1.065081e-32, 1.060006e-32, 1.079449e-32, 1.073848e-32, 1.09011e-32, 
    1.085999e-32, 1.089916e-32, 1.088728e-32, 1.089931e-32, 1.083907e-32, 
    1.086484e-32, 1.081199e-32, 1.060953e-32, 1.066776e-32, 1.04964e-32, 
    1.03968e-32, 1.033128e-32, 1.028594e-32, 1.029212e-32, 1.030424e-32, 
    1.036827e-32, 1.042912e-32, 1.04757e-32, 1.050695e-32, 1.05383e-32, 
    1.063433e-32, 1.06867e-32, 1.080581e-32, 1.078428e-32, 1.082082e-32, 
    1.085591e-32, 1.091497e-32, 1.090524e-32, 1.093132e-32, 1.08199e-32, 
    1.089381e-32, 1.077203e-32, 1.080521e-32, 1.054669e-32, 1.045319e-32, 
    1.041377e-32, 1.037954e-32, 1.0297e-32, 1.035377e-32, 1.033117e-32, 
    1.038507e-32, 1.041942e-32, 1.040243e-32, 1.050781e-32, 1.046671e-32, 
    1.068984e-32, 1.059203e-32, 1.085181e-32, 1.07887e-32, 1.086699e-32, 
    1.082699e-32, 1.089559e-32, 1.083384e-32, 1.094105e-32, 1.09645e-32, 
    1.094847e-32, 1.101024e-32, 1.083041e-32, 1.089914e-32, 1.040194e-32, 
    1.040471e-32, 1.041764e-32, 1.03609e-32, 1.035745e-32, 1.030601e-32, 
    1.035176e-32, 1.037139e-32, 1.042144e-32, 1.04511e-32, 1.047939e-32, 
    1.05424e-32, 1.061415e-32, 1.071729e-32, 1.079278e-32, 1.084365e-32, 
    1.081245e-32, 1.083998e-32, 1.08092e-32, 1.07948e-32, 1.095569e-32, 
    1.086507e-32, 1.100134e-32, 1.099377e-32, 1.093193e-32, 1.099462e-32, 
    1.040666e-32, 1.039073e-32, 1.033551e-32, 1.03787e-32, 1.030055e-32, 
    1.034403e-32, 1.036932e-32, 1.046752e-32, 1.048927e-32, 1.05094e-32, 
    1.055004e-32, 1.060265e-32, 1.069688e-32, 1.07808e-32, 1.085796e-32, 
    1.08523e-32, 1.085429e-32, 1.087156e-32, 1.082878e-32, 1.08786e-32, 
    1.088696e-32, 1.086508e-32, 1.099275e-32, 1.095614e-32, 1.099361e-32, 
    1.096976e-32, 1.039591e-32, 1.042275e-32, 1.040824e-32, 1.043554e-32, 
    1.041628e-32, 1.05021e-32, 1.052819e-32, 1.065295e-32, 1.06016e-32, 
    1.068438e-32, 1.06099e-32, 1.062287e-32, 1.068705e-32, 1.061387e-32, 
    1.077612e-32, 1.066503e-32, 1.087224e-32, 1.076033e-32, 1.087928e-32, 
    1.085763e-32, 1.089352e-32, 1.092573e-32, 1.096642e-32, 1.104178e-32, 
    1.10243e-32, 1.108762e-32, 1.046291e-32, 1.049793e-32, 1.049488e-32, 
    1.053198e-32, 1.055989e-32, 1.062065e-32, 1.072082e-32, 1.068272e-32, 
    1.075281e-32, 1.076691e-32, 1.066049e-32, 1.072568e-32, 1.052154e-32, 
    1.055388e-32, 1.053464e-32, 1.046565e-32, 1.069143e-32, 1.057377e-32, 
    1.079403e-32, 1.072831e-32, 1.092113e-32, 1.082481e-32, 1.101467e-32, 
    1.109664e-32, 1.117488e-32, 1.126912e-32, 1.051713e-32, 1.049328e-32, 
    1.053648e-32, 1.059724e-32, 1.065412e-32, 1.07323e-32, 1.074035e-32, 
    1.075505e-32, 1.079326e-32, 1.082547e-32, 1.075966e-32, 1.083356e-32, 
    1.056131e-32, 1.070193e-32, 1.048424e-32, 1.05483e-32, 1.059366e-32, 
    1.057378e-32, 1.067838e-32, 1.070372e-32, 1.08072e-32, 1.075362e-32, 
    1.107632e-32, 1.093249e-32, 1.134241e-32, 1.122377e-32, 1.048495e-32, 
    1.051706e-32, 1.06321e-32, 1.057722e-32, 1.073756e-32, 1.07779e-32, 
    1.081083e-32, 1.085299e-32, 1.085758e-32, 1.088265e-32, 1.08416e-32, 
    1.088104e-32, 1.073246e-32, 1.079864e-32, 1.061894e-32, 1.066167e-32, 
    1.064186e-32, 1.062044e-32, 1.068769e-32, 1.076068e-32, 1.076231e-32, 
    1.078581e-32, 1.085214e-32, 1.073822e-32, 1.109488e-32, 1.087327e-32, 
    1.055299e-32, 1.061666e-32, 1.062587e-32, 1.060113e-32, 1.077385e-32, 
    1.071041e-32, 1.088205e-32, 1.083543e-32, 1.091192e-32, 1.087385e-32, 
    1.086825e-32, 1.081956e-32, 1.078933e-32, 1.07133e-32, 1.065184e-32, 
    1.060472e-32, 1.061565e-32, 1.066792e-32, 1.076518e-32, 1.085797e-32, 
    1.083757e-32, 1.090609e-32, 1.072569e-32, 1.080097e-32, 1.07718e-32, 
    1.084803e-32, 1.068169e-32, 1.082299e-32, 1.0646e-32, 1.066126e-32, 
    1.070916e-32, 1.080605e-32, 1.082769e-32, 1.085072e-32, 1.083652e-32, 
    1.076767e-32, 1.075646e-32, 1.070801e-32, 1.069463e-32, 1.065791e-32, 
    1.062824e-32, 1.065527e-32, 1.068442e-32, 1.076773e-32, 1.084326e-32, 
    1.092618e-32, 1.094658e-32, 1.104418e-32, 1.096458e-32, 1.109611e-32, 
    1.098406e-32, 1.11793e-32, 1.083133e-32, 1.098091e-32, 1.071136e-32, 
    1.074013e-32, 1.079227e-32, 1.091285e-32, 1.084767e-32, 1.092396e-32, 
    1.075602e-32, 1.066973e-32, 1.064772e-32, 1.060756e-32, 1.064864e-32, 
    1.064529e-32, 1.068568e-32, 1.067262e-32, 1.07705e-32, 1.071783e-32, 
    1.086809e-32, 1.092338e-32, 1.108095e-32, 1.117905e-32, 1.128242e-32, 
    1.132893e-32, 1.134323e-32, 1.13492e-32,
  1.498526e-38, 1.514098e-38, 1.511058e-38, 1.523718e-38, 1.516684e-38, 
    1.524992e-38, 1.501668e-38, 1.514717e-38, 1.506375e-38, 1.49992e-38, 
    1.548883e-38, 1.524287e-38, 1.575538e-38, 1.559063e-38, 1.601476e-38, 
    1.57294e-38, 1.607332e-38, 1.60065e-38, 1.620879e-38, 1.615055e-38, 
    1.641223e-38, 1.623575e-38, 1.654992e-38, 1.636994e-38, 1.639791e-38, 
    1.622995e-38, 1.529155e-38, 1.545744e-38, 1.528188e-38, 1.530513e-38, 
    1.529471e-38, 1.516826e-38, 1.510491e-38, 1.497366e-38, 1.499722e-38, 
    1.509387e-38, 1.53156e-38, 1.524e-38, 1.543273e-38, 1.542826e-38, 
    1.565056e-38, 1.554987e-38, 1.59367e-38, 1.58236e-38, 1.615298e-38, 
    1.606942e-38, 1.614902e-38, 1.612485e-38, 1.614934e-38, 1.602699e-38, 
    1.607928e-38, 1.597211e-38, 1.556865e-38, 1.568389e-38, 1.534512e-38, 
    1.515016e-38, 1.502236e-38, 1.493344e-38, 1.494569e-38, 1.496953e-38, 
    1.509444e-38, 1.521327e-38, 1.530448e-38, 1.536581e-38, 1.542761e-38, 
    1.561796e-38, 1.572112e-38, 1.595964e-38, 1.591607e-38, 1.599002e-38, 
    1.606113e-38, 1.618122e-38, 1.61614e-38, 1.621453e-38, 1.598812e-38, 
    1.613817e-38, 1.589129e-38, 1.595838e-38, 1.544433e-38, 1.526037e-38, 
    1.51833e-38, 1.511641e-38, 1.49553e-38, 1.506618e-38, 1.502215e-38, 
    1.512719e-38, 1.51943e-38, 1.516108e-38, 1.536749e-38, 1.528687e-38, 
    1.572729e-38, 1.553397e-38, 1.605282e-38, 1.592501e-38, 1.608364e-38, 
    1.600249e-38, 1.614179e-38, 1.601636e-38, 1.623438e-38, 1.628226e-38, 
    1.624952e-38, 1.63758e-38, 1.600943e-38, 1.6149e-38, 1.516014e-38, 
    1.516555e-38, 1.519082e-38, 1.508007e-38, 1.507334e-38, 1.4973e-38, 
    1.506225e-38, 1.510051e-38, 1.519823e-38, 1.525629e-38, 1.531174e-38, 
    1.543573e-38, 1.557785e-38, 1.578127e-38, 1.593325e-38, 1.603625e-38, 
    1.597303e-38, 1.602883e-38, 1.596645e-38, 1.593732e-38, 1.626428e-38, 
    1.607975e-38, 1.635757e-38, 1.634207e-38, 1.621578e-38, 1.634381e-38, 
    1.516935e-38, 1.513823e-38, 1.50306e-38, 1.511476e-38, 1.496227e-38, 
    1.50472e-38, 1.509649e-38, 1.528849e-38, 1.53311e-38, 1.537063e-38, 
    1.545084e-38, 1.5555e-38, 1.57411e-38, 1.590905e-38, 1.606529e-38, 
    1.605379e-38, 1.605784e-38, 1.609293e-38, 1.600613e-38, 1.610723e-38, 
    1.612424e-38, 1.607976e-38, 1.633999e-38, 1.626517e-38, 1.634174e-38, 
    1.629298e-38, 1.514835e-38, 1.520081e-38, 1.517243e-38, 1.522583e-38, 
    1.518817e-38, 1.535633e-38, 1.54077e-38, 1.565484e-38, 1.555293e-38, 
    1.571655e-38, 1.556938e-38, 1.559513e-38, 1.572185e-38, 1.557725e-38, 
    1.589961e-38, 1.567856e-38, 1.609429e-38, 1.586776e-38, 1.61086e-38, 
    1.606461e-38, 1.613754e-38, 1.620314e-38, 1.628615e-38, 1.644049e-38, 
    1.640462e-38, 1.653469e-38, 1.527942e-38, 1.534812e-38, 1.534211e-38, 
    1.541513e-38, 1.547031e-38, 1.559071e-38, 1.578821e-38, 1.571325e-38, 
    1.58525e-38, 1.588097e-38, 1.566959e-38, 1.579785e-38, 1.539452e-38, 
    1.545846e-38, 1.54204e-38, 1.528479e-38, 1.573041e-38, 1.549781e-38, 
    1.593577e-38, 1.580312e-38, 1.619376e-38, 1.59981e-38, 1.638489e-38, 
    1.65533e-38, 1.671444e-38, 1.690976e-38, 1.538582e-38, 1.533897e-38, 
    1.542401e-38, 1.55443e-38, 1.56571e-38, 1.581117e-38, 1.582738e-38, 
    1.585704e-38, 1.593421e-38, 1.59994e-38, 1.586637e-38, 1.601579e-38, 
    1.547322e-38, 1.575104e-38, 1.532125e-38, 1.544743e-38, 1.553721e-38, 
    1.549781e-38, 1.570472e-38, 1.575453e-38, 1.596244e-38, 1.585414e-38, 
    1.65115e-38, 1.621696e-38, 1.70646e-38, 1.681471e-38, 1.532262e-38, 
    1.538568e-38, 1.561347e-38, 1.550462e-38, 1.582175e-38, 1.590318e-38, 
    1.596976e-38, 1.605523e-38, 1.606453e-38, 1.611546e-38, 1.60321e-38, 
    1.611218e-38, 1.58115e-38, 1.59451e-38, 1.558731e-38, 1.567191e-38, 
    1.563278e-38, 1.559028e-38, 1.572301e-38, 1.586844e-38, 1.587169e-38, 
    1.591917e-38, 1.605364e-38, 1.582309e-38, 1.654978e-38, 1.609652e-38, 
    1.545665e-38, 1.558284e-38, 1.560107e-38, 1.555197e-38, 1.589499e-38, 
    1.576772e-38, 1.611423e-38, 1.601959e-38, 1.6175e-38, 1.609756e-38, 
    1.608619e-38, 1.598744e-38, 1.592627e-38, 1.577341e-38, 1.56526e-38, 
    1.555909e-38, 1.558078e-38, 1.568419e-38, 1.587751e-38, 1.606533e-38, 
    1.602397e-38, 1.616313e-38, 1.579784e-38, 1.594984e-38, 1.589087e-38, 
    1.604515e-38, 1.571124e-38, 1.599452e-38, 1.564101e-38, 1.56711e-38, 
    1.576525e-38, 1.596014e-38, 1.600391e-38, 1.605063e-38, 1.60218e-38, 
    1.588253e-38, 1.585988e-38, 1.576298e-38, 1.573668e-38, 1.566451e-38, 
    1.560577e-38, 1.565934e-38, 1.571662e-38, 1.588263e-38, 1.603549e-38, 
    1.620406e-38, 1.624566e-38, 1.644548e-38, 1.628248e-38, 1.655233e-38, 
    1.632239e-38, 1.672361e-38, 1.601136e-38, 1.631587e-38, 1.576958e-38, 
    1.582693e-38, 1.593225e-38, 1.617695e-38, 1.604442e-38, 1.619958e-38, 
    1.5859e-38, 1.568776e-38, 1.564442e-38, 1.556474e-38, 1.564624e-38, 
    1.56396e-38, 1.571906e-38, 1.569341e-38, 1.588823e-38, 1.578231e-38, 
    1.608588e-38, 1.619837e-38, 1.652097e-38, 1.672301e-38, 1.693771e-38, 
    1.7036e-38, 1.706631e-38, 1.707899e-38,
  8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 9.809089e-45, 9.809089e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 9.809089e-45, 9.809089e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 9.809089e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 8.407791e-45, 
    8.407791e-45, 8.407791e-45, 8.407791e-45, 9.809089e-45, 9.809089e-45, 
    9.809089e-45, 9.809089e-45, 9.809089e-45,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  2.055999e-05, 2.037014e-05, 2.040709e-05, 2.025364e-05, 2.033882e-05, 
    2.023826e-05, 2.052155e-05, 2.036258e-05, 2.046412e-05, 2.054293e-05, 
    1.995479e-05, 2.024679e-05, 1.965022e-05, 1.983742e-05, 1.936624e-05, 
    1.967938e-05, 1.930293e-05, 1.937531e-05, 1.915729e-05, 1.921982e-05, 
    1.894021e-05, 1.912842e-05, 1.879488e-05, 1.898521e-05, 1.895546e-05, 
    1.913462e-05, 2.018814e-05, 1.999121e-05, 2.019979e-05, 2.017175e-05, 
    2.018434e-05, 2.033705e-05, 2.041386e-05, 2.057449e-05, 2.054536e-05, 
    2.042738e-05, 2.015914e-05, 2.025033e-05, 2.00203e-05, 2.002551e-05, 
    1.97685e-05, 1.98845e-05, 1.945109e-05, 1.957455e-05, 1.921721e-05, 
    1.930725e-05, 1.922144e-05, 1.924747e-05, 1.92211e-05, 1.93531e-05, 
    1.929657e-05, 1.941262e-05, 1.986278e-05, 1.973078e-05, 2.012371e-05, 
    2.035883e-05, 2.051459e-05, 2.062487e-05, 2.060929e-05, 2.057958e-05, 
    2.042669e-05, 2.028262e-05, 2.017262e-05, 2.009894e-05, 2.002625e-05, 
    1.980572e-05, 1.968875e-05, 1.942609e-05, 1.947358e-05, 1.939312e-05, 
    1.93162e-05, 1.918684e-05, 1.920815e-05, 1.915109e-05, 1.939526e-05, 
    1.923307e-05, 1.950061e-05, 1.942754e-05, 2.000642e-05, 2.022574e-05, 
    2.031869e-05, 2.039999e-05, 2.059731e-05, 2.04611e-05, 2.051483e-05, 
    2.038695e-05, 2.030556e-05, 2.034583e-05, 2.009692e-05, 2.01938e-05, 
    1.968181e-05, 1.990282e-05, 1.932517e-05, 1.946384e-05, 1.92919e-05, 
    1.937969e-05, 1.92292e-05, 1.936466e-05, 1.912985e-05, 1.907862e-05, 
    1.911363e-05, 1.897905e-05, 1.937216e-05, 1.922143e-05, 2.034696e-05, 
    2.034039e-05, 2.03098e-05, 2.044417e-05, 2.045239e-05, 2.057529e-05, 
    2.046595e-05, 2.041932e-05, 2.030085e-05, 2.023065e-05, 2.016386e-05, 
    2.001678e-05, 1.985211e-05, 1.962121e-05, 1.945486e-05, 1.934312e-05, 
    1.941166e-05, 1.935116e-05, 1.941879e-05, 1.945047e-05, 1.909781e-05, 
    1.929604e-05, 1.899843e-05, 1.901493e-05, 1.914973e-05, 1.901307e-05, 
    2.033578e-05, 2.037356e-05, 2.050454e-05, 2.040206e-05, 2.058866e-05, 
    2.048427e-05, 2.042416e-05, 2.019176e-05, 2.014061e-05, 2.009312e-05, 
    1.999924e-05, 1.987856e-05, 1.966635e-05, 1.948118e-05, 1.931172e-05, 
    1.932415e-05, 1.931978e-05, 1.928186e-05, 1.937573e-05, 1.926644e-05, 
    1.924808e-05, 1.929607e-05, 1.901714e-05, 1.909694e-05, 1.901528e-05, 
    1.906725e-05, 2.036128e-05, 2.029769e-05, 2.033206e-05, 2.026741e-05, 
    2.031296e-05, 2.011018e-05, 2.004926e-05, 1.97635e-05, 1.988094e-05, 
    1.969395e-05, 1.986197e-05, 1.983223e-05, 1.968782e-05, 1.985291e-05, 
    1.949139e-05, 1.973667e-05, 1.928039e-05, 1.952604e-05, 1.926497e-05, 
    1.931246e-05, 1.923382e-05, 1.916331e-05, 1.907452e-05, 1.891038e-05, 
    1.894843e-05, 1.881097e-05, 2.020279e-05, 2.012009e-05, 2.012739e-05, 
    2.004075e-05, 1.997661e-05, 1.983738e-05, 1.961347e-05, 1.969776e-05, 
    1.954295e-05, 1.951183e-05, 1.974699e-05, 1.960269e-05, 2.00647e-05, 
    1.999025e-05, 2.003459e-05, 2.019626e-05, 1.967833e-05, 1.994462e-05, 
    1.94521e-05, 1.959696e-05, 1.917336e-05, 1.938433e-05, 1.896936e-05, 
    1.879121e-05, 1.862321e-05, 1.842635e-05, 2.007493e-05, 2.013117e-05, 
    2.003045e-05, 1.989082e-05, 1.976106e-05, 1.958813e-05, 1.957042e-05, 
    1.953797e-05, 1.945385e-05, 1.938303e-05, 1.952769e-05, 1.936527e-05, 
    1.997295e-05, 1.965517e-05, 2.01524e-05, 2.000304e-05, 1.989907e-05, 
    1.994471e-05, 1.970739e-05, 1.965133e-05, 1.942306e-05, 1.954116e-05, 
    1.88352e-05, 1.914839e-05, 1.827616e-05, 1.852091e-05, 2.01508e-05, 
    2.007513e-05, 1.981107e-05, 1.993684e-05, 1.957658e-05, 1.948761e-05, 
    1.941521e-05, 1.932254e-05, 1.931253e-05, 1.925756e-05, 1.934762e-05, 
    1.926112e-05, 1.958776e-05, 1.944198e-05, 1.984132e-05, 1.974433e-05, 
    1.978897e-05, 1.983789e-05, 1.968679e-05, 1.952541e-05, 1.952198e-05, 
    1.947015e-05, 1.932386e-05, 1.957512e-05, 1.879465e-05, 1.927761e-05, 
    1.999251e-05, 1.98463e-05, 1.982542e-05, 1.98821e-05, 1.949653e-05, 
    1.963649e-05, 1.92589e-05, 1.936115e-05, 1.919355e-05, 1.927688e-05, 
    1.928913e-05, 1.939601e-05, 1.946246e-05, 1.963007e-05, 1.976616e-05, 
    1.987389e-05, 1.984885e-05, 1.973046e-05, 1.951553e-05, 1.931162e-05, 
    1.935633e-05, 1.92063e-05, 1.960276e-05, 1.943678e-05, 1.950097e-05, 
    1.933347e-05, 1.969999e-05, 1.938794e-05, 1.977953e-05, 1.974529e-05, 
    1.963926e-05, 1.942549e-05, 1.937814e-05, 1.932751e-05, 1.935876e-05, 
    1.951007e-05, 1.953484e-05, 1.964184e-05, 1.967135e-05, 1.975274e-05, 
    1.982005e-05, 1.975855e-05, 1.969391e-05, 1.951002e-05, 1.934388e-05, 
    1.91623e-05, 1.91178e-05, 1.890489e-05, 1.907823e-05, 1.879194e-05, 
    1.903537e-05, 1.861351e-05, 1.936984e-05, 1.904256e-05, 1.963444e-05, 
    1.957092e-05, 1.945585e-05, 1.919128e-05, 1.933426e-05, 1.916703e-05, 
    1.953581e-05, 1.972636e-05, 1.977561e-05, 1.986734e-05, 1.977351e-05, 
    1.978114e-05, 1.969124e-05, 1.972015e-05, 1.95039e-05, 1.962014e-05, 
    1.928943e-05, 1.916836e-05, 1.882538e-05, 1.861432e-05, 1.839891e-05, 
    1.830361e-05, 1.827459e-05, 1.826245e-05,
  1.428218e-05, 1.409153e-05, 1.412862e-05, 1.397467e-05, 1.40601e-05, 
    1.395925e-05, 1.424356e-05, 1.408394e-05, 1.418587e-05, 1.426504e-05, 
    1.367537e-05, 1.39678e-05, 1.337113e-05, 1.355805e-05, 1.308815e-05, 
    1.340021e-05, 1.302517e-05, 1.309719e-05, 1.288043e-05, 1.294255e-05, 
    1.2665e-05, 1.285175e-05, 1.252107e-05, 1.270963e-05, 1.268013e-05, 
    1.28579e-05, 1.390903e-05, 1.37118e-05, 1.39207e-05, 1.389259e-05, 
    1.390521e-05, 1.405833e-05, 1.41354e-05, 1.429676e-05, 1.426749e-05, 
    1.414898e-05, 1.387996e-05, 1.397136e-05, 1.374095e-05, 1.374615e-05, 
    1.34892e-05, 1.360511e-05, 1.317264e-05, 1.329567e-05, 1.293996e-05, 
    1.302947e-05, 1.294416e-05, 1.297003e-05, 1.294382e-05, 1.307509e-05, 
    1.301886e-05, 1.313433e-05, 1.35834e-05, 1.345154e-05, 1.384447e-05, 
    1.408017e-05, 1.423656e-05, 1.43474e-05, 1.433173e-05, 1.430186e-05, 
    1.414828e-05, 1.400374e-05, 1.389348e-05, 1.381966e-05, 1.37469e-05, 
    1.352636e-05, 1.340957e-05, 1.314774e-05, 1.319504e-05, 1.311492e-05, 
    1.303838e-05, 1.290977e-05, 1.293095e-05, 1.287426e-05, 1.311705e-05, 
    1.295571e-05, 1.322198e-05, 1.314919e-05, 1.372701e-05, 1.394671e-05, 
    1.40399e-05, 1.412149e-05, 1.431969e-05, 1.418284e-05, 1.42368e-05, 
    1.410841e-05, 1.402674e-05, 1.406715e-05, 1.381765e-05, 1.39147e-05, 
    1.340265e-05, 1.362342e-05, 1.30473e-05, 1.318534e-05, 1.301421e-05, 
    1.310156e-05, 1.295186e-05, 1.308659e-05, 1.285317e-05, 1.28023e-05, 
    1.283706e-05, 1.270353e-05, 1.309405e-05, 1.294415e-05, 1.406827e-05, 
    1.406168e-05, 1.4031e-05, 1.416584e-05, 1.417409e-05, 1.429756e-05, 
    1.418771e-05, 1.41409e-05, 1.402202e-05, 1.395163e-05, 1.38847e-05, 
    1.373741e-05, 1.357273e-05, 1.334219e-05, 1.317639e-05, 1.306517e-05, 
    1.313338e-05, 1.307316e-05, 1.314048e-05, 1.317203e-05, 1.282136e-05, 
    1.301832e-05, 1.272274e-05, 1.273911e-05, 1.287291e-05, 1.273727e-05, 
    1.405706e-05, 1.409497e-05, 1.422647e-05, 1.412357e-05, 1.431099e-05, 
    1.42061e-05, 1.414575e-05, 1.391265e-05, 1.38614e-05, 1.381383e-05, 
    1.371987e-05, 1.359918e-05, 1.338722e-05, 1.32026e-05, 1.303393e-05, 
    1.304629e-05, 1.304194e-05, 1.300423e-05, 1.309761e-05, 1.298889e-05, 
    1.297063e-05, 1.301836e-05, 1.27413e-05, 1.282049e-05, 1.273946e-05, 
    1.279103e-05, 1.408265e-05, 1.401885e-05, 1.405333e-05, 1.398849e-05, 
    1.403416e-05, 1.383091e-05, 1.376992e-05, 1.34842e-05, 1.360155e-05, 
    1.341477e-05, 1.358259e-05, 1.355286e-05, 1.340863e-05, 1.357353e-05, 
    1.321277e-05, 1.34574e-05, 1.300276e-05, 1.324729e-05, 1.298743e-05, 
    1.303466e-05, 1.295646e-05, 1.28864e-05, 1.279824e-05, 1.263546e-05, 
    1.267317e-05, 1.2537e-05, 1.39237e-05, 1.384084e-05, 1.384816e-05, 
    1.376141e-05, 1.369722e-05, 1.355802e-05, 1.333448e-05, 1.341858e-05, 
    1.326417e-05, 1.323315e-05, 1.346773e-05, 1.332372e-05, 1.378538e-05, 
    1.371086e-05, 1.375525e-05, 1.391716e-05, 1.339918e-05, 1.366521e-05, 
    1.317365e-05, 1.331801e-05, 1.289639e-05, 1.310616e-05, 1.269392e-05, 
    1.251742e-05, 1.235132e-05, 1.2157e-05, 1.379562e-05, 1.385194e-05, 
    1.37511e-05, 1.361142e-05, 1.348177e-05, 1.330921e-05, 1.329155e-05, 
    1.32592e-05, 1.317539e-05, 1.310488e-05, 1.324895e-05, 1.30872e-05, 
    1.369354e-05, 1.337607e-05, 1.387321e-05, 1.372366e-05, 1.361967e-05, 
    1.366531e-05, 1.342819e-05, 1.337225e-05, 1.314473e-05, 1.326239e-05, 
    1.256098e-05, 1.287157e-05, 1.200905e-05, 1.225029e-05, 1.387161e-05, 
    1.379582e-05, 1.353172e-05, 1.365744e-05, 1.329769e-05, 1.320902e-05, 
    1.313692e-05, 1.304468e-05, 1.303473e-05, 1.298006e-05, 1.306964e-05, 
    1.298361e-05, 1.330884e-05, 1.316357e-05, 1.356196e-05, 1.346507e-05, 
    1.350965e-05, 1.355853e-05, 1.340763e-05, 1.324668e-05, 1.324327e-05, 
    1.319162e-05, 1.304595e-05, 1.329624e-05, 1.252081e-05, 1.299996e-05, 
    1.371313e-05, 1.356692e-05, 1.354606e-05, 1.360272e-05, 1.321791e-05, 
    1.335743e-05, 1.29814e-05, 1.30831e-05, 1.291644e-05, 1.299927e-05, 
    1.301145e-05, 1.311779e-05, 1.318396e-05, 1.335103e-05, 1.348686e-05, 
    1.359451e-05, 1.356949e-05, 1.345122e-05, 1.323683e-05, 1.303381e-05, 
    1.30783e-05, 1.292911e-05, 1.33238e-05, 1.315838e-05, 1.322232e-05, 
    1.305556e-05, 1.342081e-05, 1.310972e-05, 1.350022e-05, 1.346603e-05, 
    1.33602e-05, 1.314714e-05, 1.310001e-05, 1.304962e-05, 1.308072e-05, 
    1.323139e-05, 1.325608e-05, 1.336278e-05, 1.339222e-05, 1.347347e-05, 
    1.35407e-05, 1.347927e-05, 1.341473e-05, 1.323134e-05, 1.306591e-05, 
    1.28854e-05, 1.284121e-05, 1.263e-05, 1.28019e-05, 1.251813e-05, 
    1.275934e-05, 1.23417e-05, 1.309173e-05, 1.27665e-05, 1.33554e-05, 
    1.329205e-05, 1.317737e-05, 1.291418e-05, 1.305634e-05, 1.289009e-05, 
    1.325705e-05, 1.344712e-05, 1.34963e-05, 1.358796e-05, 1.349421e-05, 
    1.350184e-05, 1.341208e-05, 1.344093e-05, 1.322525e-05, 1.334114e-05, 
    1.301175e-05, 1.289141e-05, 1.255126e-05, 1.234252e-05, 1.212997e-05, 
    1.203608e-05, 1.200751e-05, 1.199556e-05,
  6.640359e-06, 6.523288e-06, 6.546026e-06, 6.451778e-06, 6.50404e-06, 
    6.44236e-06, 6.616606e-06, 6.51864e-06, 6.581158e-06, 6.629817e-06, 
    6.269494e-06, 6.447581e-06, 6.0855e-06, 6.198387e-06, 5.91556e-06, 
    6.103031e-06, 5.877897e-06, 5.920971e-06, 5.791559e-06, 5.828577e-06, 
    5.663641e-06, 5.774491e-06, 5.578557e-06, 5.690084e-06, 5.672599e-06, 
    5.778152e-06, 6.411693e-06, 6.291615e-06, 6.418815e-06, 6.401667e-06, 
    6.409365e-06, 6.502953e-06, 6.550186e-06, 6.649332e-06, 6.631319e-06, 
    6.558514e-06, 6.393959e-06, 6.449754e-06, 6.309325e-06, 6.312491e-06, 
    6.156748e-06, 6.226885e-06, 5.966177e-06, 6.040071e-06, 5.827032e-06, 
    5.880467e-06, 5.829536e-06, 5.844973e-06, 5.829335e-06, 5.907744e-06, 
    5.874124e-06, 5.943216e-06, 6.213735e-06, 6.133999e-06, 6.372326e-06, 
    6.516329e-06, 6.612302e-06, 6.680521e-06, 6.67087e-06, 6.652474e-06, 
    6.558088e-06, 6.469552e-06, 6.402206e-06, 6.357218e-06, 6.312946e-06, 
    6.179213e-06, 6.108676e-06, 5.951248e-06, 5.979617e-06, 5.931584e-06, 
    5.885789e-06, 5.809037e-06, 5.821659e-06, 5.78789e-06, 5.932862e-06, 
    5.836429e-06, 5.995784e-06, 5.952115e-06, 6.300857e-06, 6.434697e-06, 
    6.491671e-06, 6.541652e-06, 6.66345e-06, 6.579299e-06, 6.612451e-06, 
    6.533635e-06, 6.483622e-06, 6.508353e-06, 6.355989e-06, 6.415151e-06, 
    6.1045e-06, 6.237982e-06, 5.891127e-06, 5.973793e-06, 5.871348e-06, 
    5.923584e-06, 5.834131e-06, 5.914626e-06, 5.775336e-06, 5.745087e-06, 
    5.765753e-06, 5.686468e-06, 5.919093e-06, 5.82953e-06, 6.509043e-06, 
    6.505008e-06, 6.486223e-06, 6.56886e-06, 6.573924e-06, 6.649823e-06, 
    6.582287e-06, 6.553555e-06, 6.48073e-06, 6.437704e-06, 6.39685e-06, 
    6.307177e-06, 6.207275e-06, 6.068069e-06, 5.968427e-06, 5.901808e-06, 
    5.942645e-06, 5.906588e-06, 5.946896e-06, 5.965809e-06, 5.756413e-06, 
    5.873807e-06, 5.697858e-06, 5.707568e-06, 5.787085e-06, 5.706474e-06, 
    6.502176e-06, 6.525397e-06, 6.606097e-06, 6.542929e-06, 6.658097e-06, 
    6.593586e-06, 6.556531e-06, 6.413901e-06, 6.382646e-06, 6.353669e-06, 
    6.296516e-06, 6.223291e-06, 6.095199e-06, 5.984154e-06, 5.883129e-06, 
    5.890521e-06, 5.887918e-06, 5.865385e-06, 5.921222e-06, 5.856229e-06, 
    5.845329e-06, 5.873828e-06, 5.708868e-06, 5.7559e-06, 5.707775e-06, 
    5.738389e-06, 6.517849e-06, 6.478795e-06, 6.499893e-06, 6.460225e-06, 
    6.488162e-06, 6.36407e-06, 6.326942e-06, 6.153725e-06, 6.224728e-06, 
    6.111811e-06, 6.213246e-06, 6.195247e-06, 6.108108e-06, 6.207761e-06, 
    5.990255e-06, 6.137541e-06, 5.86451e-06, 6.010987e-06, 5.855353e-06, 
    5.883565e-06, 5.836875e-06, 5.795115e-06, 5.742674e-06, 5.646151e-06, 
    5.668475e-06, 5.58796e-06, 6.420648e-06, 6.370118e-06, 6.374576e-06, 
    6.321769e-06, 6.282759e-06, 6.198367e-06, 6.063424e-06, 6.114109e-06, 
    6.021131e-06, 6.002493e-06, 6.143779e-06, 6.056949e-06, 6.336346e-06, 
    6.291045e-06, 6.318019e-06, 6.416653e-06, 6.102406e-06, 6.263332e-06, 
    5.966781e-06, 6.053514e-06, 5.801064e-06, 5.926342e-06, 5.680769e-06, 
    5.576409e-06, 5.478621e-06, 5.364763e-06, 6.34258e-06, 6.376882e-06, 
    6.315497e-06, 6.230712e-06, 6.152257e-06, 6.048215e-06, 6.037595e-06, 
    6.018142e-06, 5.967825e-06, 5.925575e-06, 6.011983e-06, 5.914994e-06, 
    6.280523e-06, 6.088479e-06, 6.389847e-06, 6.29882e-06, 6.235709e-06, 
    6.263393e-06, 6.11991e-06, 6.086175e-06, 5.949442e-06, 6.02006e-06, 
    5.602119e-06, 5.786285e-06, 5.278469e-06, 5.419351e-06, 6.388871e-06, 
    6.342704e-06, 6.182457e-06, 6.258616e-06, 6.041287e-06, 5.988003e-06, 
    5.944762e-06, 5.889555e-06, 5.88361e-06, 5.850955e-06, 5.904482e-06, 
    5.853072e-06, 6.047994e-06, 5.960739e-06, 6.200751e-06, 6.142169e-06, 
    6.16911e-06, 6.198678e-06, 6.107502e-06, 6.010618e-06, 6.00857e-06, 
    5.977563e-06, 5.890321e-06, 6.04041e-06, 5.578405e-06, 5.862838e-06, 
    6.292425e-06, 6.203755e-06, 6.191131e-06, 6.225437e-06, 5.99334e-06, 
    6.077249e-06, 5.851753e-06, 5.91254e-06, 5.813012e-06, 5.862426e-06, 
    5.869702e-06, 5.933307e-06, 5.972968e-06, 6.073394e-06, 6.155336e-06, 
    6.220462e-06, 6.205309e-06, 6.133807e-06, 6.004705e-06, 5.883063e-06, 
    5.909666e-06, 5.820564e-06, 6.056998e-06, 5.957628e-06, 5.995992e-06, 
    5.896062e-06, 6.115453e-06, 5.928477e-06, 6.163409e-06, 6.142748e-06, 
    6.078917e-06, 5.950887e-06, 5.922659e-06, 5.892514e-06, 5.911115e-06, 
    6.001438e-06, 6.016269e-06, 6.080472e-06, 6.098211e-06, 6.147246e-06, 
    6.187888e-06, 6.150749e-06, 6.111786e-06, 6.001408e-06, 5.902251e-06, 
    5.794518e-06, 5.76822e-06, 5.642922e-06, 5.744852e-06, 5.576826e-06, 
    5.719575e-06, 5.472972e-06, 5.917703e-06, 5.723823e-06, 6.076022e-06, 
    6.037891e-06, 5.969016e-06, 5.811663e-06, 5.896532e-06, 5.797312e-06, 
    6.016851e-06, 6.131334e-06, 6.16104e-06, 6.216495e-06, 6.159773e-06, 
    6.164384e-06, 6.110186e-06, 6.127595e-06, 5.99775e-06, 6.067434e-06, 
    5.86988e-06, 5.798099e-06, 5.59638e-06, 5.473455e-06, 5.348971e-06, 
    5.29421e-06, 5.277569e-06, 5.270615e-06,
  1.675916e-06, 1.632467e-06, 1.640877e-06, 1.606111e-06, 1.625359e-06, 
    1.602649e-06, 1.66707e-06, 1.63075e-06, 1.653898e-06, 1.671988e-06, 
    1.539561e-06, 1.604568e-06, 1.473319e-06, 1.513847e-06, 1.412986e-06, 
    1.47959e-06, 1.399726e-06, 1.414894e-06, 1.369484e-06, 1.382424e-06, 
    1.325075e-06, 1.36353e-06, 1.295802e-06, 1.334216e-06, 1.328169e-06, 
    1.364807e-06, 1.591397e-06, 1.547588e-06, 1.594008e-06, 1.587724e-06, 
    1.590544e-06, 1.624958e-06, 1.642417e-06, 1.679261e-06, 1.672547e-06, 
    1.645501e-06, 1.584902e-06, 1.605366e-06, 1.554022e-06, 1.555174e-06, 
    1.498856e-06, 1.524135e-06, 1.43087e-06, 1.45711e-06, 1.381883e-06, 
    1.400629e-06, 1.38276e-06, 1.388168e-06, 1.382689e-06, 1.410231e-06, 
    1.3984e-06, 1.422748e-06, 1.519385e-06, 1.490687e-06, 1.57699e-06, 
    1.629897e-06, 1.665469e-06, 1.690906e-06, 1.6873e-06, 1.680433e-06, 
    1.645344e-06, 1.612648e-06, 1.587921e-06, 1.571472e-06, 1.55534e-06, 
    1.506939e-06, 1.481611e-06, 1.425588e-06, 1.435631e-06, 1.41864e-06, 
    1.402501e-06, 1.375589e-06, 1.380002e-06, 1.368203e-06, 1.41909e-06, 
    1.385174e-06, 1.441364e-06, 1.425894e-06, 1.550946e-06, 1.599835e-06, 
    1.620797e-06, 1.639258e-06, 1.684529e-06, 1.653208e-06, 1.665525e-06, 
    1.636292e-06, 1.61783e-06, 1.62695e-06, 1.571024e-06, 1.592664e-06, 
    1.480115e-06, 1.528147e-06, 1.404379e-06, 1.433567e-06, 1.397424e-06, 
    1.415816e-06, 1.384369e-06, 1.412656e-06, 1.363825e-06, 1.353295e-06, 
    1.360487e-06, 1.332964e-06, 1.414231e-06, 1.382758e-06, 1.627205e-06, 
    1.625716e-06, 1.618788e-06, 1.649336e-06, 1.651214e-06, 1.679444e-06, 
    1.654317e-06, 1.643665e-06, 1.616764e-06, 1.600939e-06, 1.58596e-06, 
    1.553242e-06, 1.517053e-06, 1.467092e-06, 1.431667e-06, 1.408139e-06, 
    1.422546e-06, 1.409823e-06, 1.424049e-06, 1.430739e-06, 1.357235e-06, 
    1.398288e-06, 1.336907e-06, 1.340271e-06, 1.367922e-06, 1.339891e-06, 
    1.624671e-06, 1.633246e-06, 1.663162e-06, 1.63973e-06, 1.682531e-06, 
    1.658512e-06, 1.644767e-06, 1.592206e-06, 1.580763e-06, 1.570177e-06, 
    1.549367e-06, 1.522836e-06, 1.476787e-06, 1.437239e-06, 1.401565e-06, 
    1.404166e-06, 1.40325e-06, 1.39533e-06, 1.414982e-06, 1.392116e-06, 
    1.388293e-06, 1.398296e-06, 1.340721e-06, 1.357056e-06, 1.340342e-06, 
    1.350966e-06, 1.630457e-06, 1.616051e-06, 1.623828e-06, 1.609216e-06, 
    1.619503e-06, 1.573974e-06, 1.560434e-06, 1.49777e-06, 1.523355e-06, 
    1.482733e-06, 1.519208e-06, 1.512715e-06, 1.481408e-06, 1.517228e-06, 
    1.439403e-06, 1.491959e-06, 1.395023e-06, 1.446764e-06, 1.391808e-06, 
    1.401719e-06, 1.38533e-06, 1.370725e-06, 1.352456e-06, 1.31904e-06, 
    1.326744e-06, 1.299026e-06, 1.59468e-06, 1.576183e-06, 1.577812e-06, 
    1.55855e-06, 1.544371e-06, 1.51384e-06, 1.465434e-06, 1.483556e-06, 
    1.450369e-06, 1.443746e-06, 1.494197e-06, 1.463125e-06, 1.56386e-06, 
    1.54738e-06, 1.557186e-06, 1.593215e-06, 1.479366e-06, 1.537326e-06, 
    1.431084e-06, 1.4619e-06, 1.372802e-06, 1.416789e-06, 1.330993e-06, 
    1.295066e-06, 1.261692e-06, 1.223195e-06, 1.566133e-06, 1.578655e-06, 
    1.556268e-06, 1.525519e-06, 1.497243e-06, 1.460011e-06, 1.456228e-06, 
    1.449307e-06, 1.431453e-06, 1.416518e-06, 1.447118e-06, 1.412786e-06, 
    1.543561e-06, 1.474383e-06, 1.583397e-06, 1.550204e-06, 1.527325e-06, 
    1.537347e-06, 1.485634e-06, 1.47356e-06, 1.424949e-06, 1.449988e-06, 
    1.303887e-06, 1.367644e-06, 1.194278e-06, 1.241604e-06, 1.58304e-06, 
    1.566178e-06, 1.508106e-06, 1.535616e-06, 1.457543e-06, 1.438604e-06, 
    1.423294e-06, 1.403826e-06, 1.401734e-06, 1.390266e-06, 1.409081e-06, 
    1.391008e-06, 1.459932e-06, 1.428945e-06, 1.514699e-06, 1.493619e-06, 
    1.503302e-06, 1.513952e-06, 1.48119e-06, 1.446633e-06, 1.445904e-06, 
    1.434903e-06, 1.404097e-06, 1.45723e-06, 1.295751e-06, 1.394437e-06, 
    1.54788e-06, 1.515784e-06, 1.511231e-06, 1.523611e-06, 1.440497e-06, 
    1.47037e-06, 1.390546e-06, 1.411921e-06, 1.376978e-06, 1.394291e-06, 
    1.396846e-06, 1.419248e-06, 1.433275e-06, 1.468993e-06, 1.498349e-06, 
    1.521814e-06, 1.516344e-06, 1.490618e-06, 1.444532e-06, 1.401542e-06, 
    1.410908e-06, 1.379619e-06, 1.463142e-06, 1.427844e-06, 1.441439e-06, 
    1.406116e-06, 1.484037e-06, 1.417544e-06, 1.501251e-06, 1.493827e-06, 
    1.470966e-06, 1.42546e-06, 1.415489e-06, 1.404867e-06, 1.411419e-06, 
    1.443372e-06, 1.448641e-06, 1.471521e-06, 1.477864e-06, 1.495442e-06, 
    1.510062e-06, 1.4967e-06, 1.482724e-06, 1.443361e-06, 1.408296e-06, 
    1.370517e-06, 1.361346e-06, 1.317928e-06, 1.353214e-06, 1.29521e-06, 
    1.344437e-06, 1.259775e-06, 1.413742e-06, 1.345909e-06, 1.469932e-06, 
    1.456333e-06, 1.431876e-06, 1.376507e-06, 1.406281e-06, 1.371493e-06, 
    1.448848e-06, 1.489731e-06, 1.500399e-06, 1.520381e-06, 1.499944e-06, 
    1.501602e-06, 1.48215e-06, 1.488389e-06, 1.442062e-06, 1.466865e-06, 
    1.396909e-06, 1.371767e-06, 1.301916e-06, 1.259938e-06, 1.217886e-06, 
    1.199536e-06, 1.193977e-06, 1.191657e-06,
  1.527441e-07, 1.469319e-07, 1.480511e-07, 1.434419e-07, 1.459879e-07, 
    1.429856e-07, 1.515549e-07, 1.467037e-07, 1.497896e-07, 1.522157e-07, 
    1.347517e-07, 1.432384e-07, 1.262781e-07, 1.314413e-07, 1.18717e-07, 
    1.270727e-07, 1.170755e-07, 1.189537e-07, 1.133594e-07, 1.149447e-07, 
    1.079736e-07, 1.126325e-07, 1.044697e-07, 1.090752e-07, 1.083461e-07, 
    1.127882e-07, 1.415054e-07, 1.357906e-07, 1.418484e-07, 1.410233e-07, 
    1.413933e-07, 1.459348e-07, 1.482565e-07, 1.531946e-07, 1.522909e-07, 
    1.486678e-07, 1.406533e-07, 1.433437e-07, 1.36625e-07, 1.367746e-07, 
    1.295236e-07, 1.327624e-07, 1.209425e-07, 1.242318e-07, 1.148783e-07, 
    1.17187e-07, 1.14986e-07, 1.156507e-07, 1.149773e-07, 1.183752e-07, 
    1.169117e-07, 1.199301e-07, 1.321519e-07, 1.284825e-07, 1.396176e-07, 
    1.465904e-07, 1.5134e-07, 1.547663e-07, 1.54279e-07, 1.533526e-07, 
    1.486468e-07, 1.443049e-07, 1.410491e-07, 1.388967e-07, 1.367961e-07, 
    1.305566e-07, 1.27329e-07, 1.202837e-07, 1.215371e-07, 1.194191e-07, 
    1.174183e-07, 1.141065e-07, 1.146475e-07, 1.13203e-07, 1.194751e-07, 
    1.152826e-07, 1.222546e-07, 1.203219e-07, 1.36226e-07, 1.426149e-07, 
    1.453833e-07, 1.478355e-07, 1.53905e-07, 1.496974e-07, 1.513475e-07, 
    1.474405e-07, 1.449903e-07, 1.461991e-07, 1.388381e-07, 1.416718e-07, 
    1.271393e-07, 1.332789e-07, 1.176506e-07, 1.212792e-07, 1.167912e-07, 
    1.190681e-07, 1.151836e-07, 1.18676e-07, 1.126685e-07, 1.113863e-07, 
    1.122615e-07, 1.089241e-07, 1.188714e-07, 1.149858e-07, 1.462329e-07, 
    1.460353e-07, 1.451171e-07, 1.491799e-07, 1.494308e-07, 1.532193e-07, 
    1.498456e-07, 1.484228e-07, 1.448492e-07, 1.427602e-07, 1.407919e-07, 
    1.365237e-07, 1.318526e-07, 1.254908e-07, 1.210419e-07, 1.18116e-07, 
    1.199049e-07, 1.183247e-07, 1.20092e-07, 1.209261e-07, 1.118655e-07, 
    1.16898e-07, 1.094002e-07, 1.098069e-07, 1.131687e-07, 1.09761e-07, 
    1.458967e-07, 1.470354e-07, 1.510304e-07, 1.478983e-07, 1.536354e-07, 
    1.504072e-07, 1.485699e-07, 1.416117e-07, 1.401111e-07, 1.387277e-07, 
    1.36021e-07, 1.325954e-07, 1.267172e-07, 1.217383e-07, 1.173027e-07, 
    1.176242e-07, 1.175109e-07, 1.165329e-07, 1.189647e-07, 1.161367e-07, 
    1.156661e-07, 1.168988e-07, 1.098614e-07, 1.118437e-07, 1.098156e-07, 
    1.111034e-07, 1.466647e-07, 1.447549e-07, 1.457849e-07, 1.438517e-07, 
    1.452118e-07, 1.392235e-07, 1.374584e-07, 1.293851e-07, 1.326622e-07, 
    1.274714e-07, 1.321292e-07, 1.312961e-07, 1.273033e-07, 1.31875e-07, 
    1.220091e-07, 1.286444e-07, 1.16495e-07, 1.229317e-07, 1.160988e-07, 
    1.173216e-07, 1.153017e-07, 1.135112e-07, 1.112843e-07, 1.072481e-07, 
    1.081744e-07, 1.048538e-07, 1.419367e-07, 1.395121e-07, 1.39725e-07, 
    1.372133e-07, 1.353738e-07, 1.314403e-07, 1.252814e-07, 1.275758e-07, 
    1.233841e-07, 1.225531e-07, 1.289295e-07, 1.2499e-07, 1.379043e-07, 
    1.357635e-07, 1.37036e-07, 1.417442e-07, 1.270442e-07, 1.344628e-07, 
    1.209691e-07, 1.248354e-07, 1.137654e-07, 1.191891e-07, 1.086864e-07, 
    1.043822e-07, 1.004344e-07, 9.594218e-08, 1.382003e-07, 1.398353e-07, 
    1.369166e-07, 1.329406e-07, 1.293178e-07, 1.245973e-07, 1.241208e-07, 
    1.232507e-07, 1.210152e-07, 1.191554e-07, 1.229759e-07, 1.186921e-07, 
    1.352691e-07, 1.264128e-07, 1.404561e-07, 1.361297e-07, 1.331731e-07, 
    1.344656e-07, 1.278398e-07, 1.263085e-07, 1.202042e-07, 1.233362e-07, 
    1.054339e-07, 1.131347e-07, 9.261151e-08, 9.808201e-08, 1.404093e-07, 
    1.382061e-07, 1.307058e-07, 1.342421e-07, 1.242864e-07, 1.21909e-07, 
    1.19998e-07, 1.175822e-07, 1.173236e-07, 1.159089e-07, 1.182327e-07, 
    1.160003e-07, 1.245874e-07, 1.207022e-07, 1.315505e-07, 1.288558e-07, 
    1.300913e-07, 1.314546e-07, 1.272755e-07, 1.229151e-07, 1.228237e-07, 
    1.214462e-07, 1.17616e-07, 1.24247e-07, 1.044639e-07, 1.16423e-07, 
    1.358283e-07, 1.316897e-07, 1.31106e-07, 1.326951e-07, 1.22146e-07, 
    1.25905e-07, 1.159433e-07, 1.185848e-07, 1.142767e-07, 1.164047e-07, 
    1.167199e-07, 1.194946e-07, 1.212427e-07, 1.25731e-07, 1.294589e-07, 
    1.32464e-07, 1.317614e-07, 1.284737e-07, 1.226516e-07, 1.172999e-07, 
    1.184592e-07, 1.146005e-07, 1.249921e-07, 1.20565e-07, 1.22264e-07, 
    1.178655e-07, 1.27637e-07, 1.19283e-07, 1.298293e-07, 1.288823e-07, 
    1.259804e-07, 1.202679e-07, 1.190276e-07, 1.17711e-07, 1.185225e-07, 
    1.225062e-07, 1.231671e-07, 1.260506e-07, 1.268538e-07, 1.290882e-07, 
    1.309562e-07, 1.292486e-07, 1.274702e-07, 1.225048e-07, 1.181355e-07, 
    1.134858e-07, 1.123661e-07, 1.071147e-07, 1.113765e-07, 1.043995e-07, 
    1.103115e-07, 1.002092e-07, 1.188108e-07, 1.104899e-07, 1.258495e-07, 
    1.241341e-07, 1.210681e-07, 1.142191e-07, 1.17886e-07, 1.136052e-07, 
    1.23193e-07, 1.283609e-07, 1.297206e-07, 1.322799e-07, 1.296624e-07, 
    1.298741e-07, 1.273974e-07, 1.281901e-07, 1.22342e-07, 1.254621e-07, 
    1.167277e-07, 1.136387e-07, 1.051985e-07, 1.002283e-07, 9.532775e-08, 
    9.321421e-08, 9.257705e-08, 9.23115e-08,
  4.410179e-09, 4.173248e-09, 4.218586e-09, 4.03276e-09, 4.135114e-09, 
    4.014493e-09, 4.361402e-09, 4.164022e-09, 4.28928e-09, 4.388484e-09, 
    3.688907e-09, 4.024612e-09, 3.362072e-09, 3.560203e-09, 3.077783e-09, 
    3.392355e-09, 3.01701e-09, 3.086574e-09, 2.8807e-09, 2.938631e-09, 
    2.686346e-09, 2.854244e-09, 2.561989e-09, 2.725783e-09, 2.699663e-09, 
    2.859906e-09, 3.955392e-09, 3.729558e-09, 3.969065e-09, 3.936199e-09, 
    3.950928e-09, 4.132972e-09, 4.226924e-09, 4.428692e-09, 4.391568e-09, 
    4.243628e-09, 3.921485e-09, 4.028824e-09, 3.762295e-09, 3.768171e-09, 
    3.486244e-09, 3.611411e-09, 3.16072e-09, 3.284437e-09, 2.936196e-09, 
    3.021126e-09, 2.940143e-09, 2.964534e-09, 2.939826e-09, 3.0651e-09, 
    3.010961e-09, 3.122914e-09, 3.587723e-09, 3.446273e-09, 3.880378e-09, 
    4.159445e-09, 4.352603e-09, 4.493462e-09, 4.473355e-09, 4.435194e-09, 
    4.242772e-09, 4.067375e-09, 3.937224e-09, 3.851839e-09, 3.769016e-09, 
    3.526032e-09, 3.40214e-09, 3.136107e-09, 3.182986e-09, 3.10388e-09, 
    3.029672e-09, 2.907959e-09, 2.927747e-09, 2.875e-09, 3.105963e-09, 
    2.95102e-09, 3.20991e-09, 3.13753e-09, 3.746633e-09, 3.999666e-09, 
    4.110747e-09, 4.20984e-09, 4.457936e-09, 4.285522e-09, 4.35291e-09, 
    4.193835e-09, 4.094922e-09, 4.143636e-09, 3.849523e-09, 3.962026e-09, 
    3.394896e-09, 3.631488e-09, 3.038261e-09, 3.173325e-09, 3.006519e-09, 
    3.090826e-09, 2.947391e-09, 3.076259e-09, 2.855552e-09, 2.809052e-09, 
    2.840767e-09, 2.720365e-09, 3.083518e-09, 2.940136e-09, 4.145003e-09, 
    4.137027e-09, 4.100026e-09, 4.264449e-09, 4.274662e-09, 4.429708e-09, 
    4.291565e-09, 4.233672e-09, 4.089248e-09, 4.005478e-09, 3.926995e-09, 
    3.758315e-09, 3.576124e-09, 3.332141e-09, 3.16444e-09, 3.055493e-09, 
    3.121976e-09, 3.063227e-09, 3.128952e-09, 3.160108e-09, 2.826406e-09, 
    3.010455e-09, 2.73745e-09, 2.75207e-09, 2.873751e-09, 2.75042e-09, 
    4.131435e-09, 4.177433e-09, 4.339939e-09, 4.212389e-09, 4.446832e-09, 
    4.314476e-09, 4.239649e-09, 3.959631e-09, 3.899949e-09, 3.845157e-09, 
    3.738585e-09, 3.604927e-09, 3.378798e-09, 3.19053e-09, 3.025398e-09, 
    3.037284e-09, 3.033095e-09, 2.996994e-09, 3.086982e-09, 2.982405e-09, 
    2.965101e-09, 3.010487e-09, 2.754032e-09, 2.825615e-09, 2.752381e-09, 
    2.798819e-09, 4.162444e-09, 4.085456e-09, 4.126929e-09, 4.049184e-09, 
    4.103838e-09, 3.864771e-09, 3.79508e-09, 3.48092e-09, 3.60752e-09, 
    3.407581e-09, 3.586841e-09, 3.55459e-09, 3.401161e-09, 3.57699e-09, 
    3.200693e-09, 3.452483e-09, 2.995597e-09, 3.23538e-09, 2.981011e-09, 
    3.026099e-09, 2.951721e-09, 2.886232e-09, 2.805362e-09, 2.660461e-09, 
    2.693521e-09, 2.575538e-09, 3.972588e-09, 3.8762e-09, 3.884636e-09, 
    3.785427e-09, 3.71323e-09, 3.560164e-09, 3.324194e-09, 3.411569e-09, 
    3.252426e-09, 3.221129e-09, 3.463415e-09, 3.313142e-09, 3.812648e-09, 
    3.728495e-09, 3.77845e-09, 3.964913e-09, 3.391267e-09, 3.677622e-09, 
    3.161718e-09, 3.307284e-09, 2.895503e-09, 3.095327e-09, 2.711845e-09, 
    2.558906e-09, 2.420862e-09, 2.266462e-09, 3.824326e-09, 3.889008e-09, 
    3.773756e-09, 3.618332e-09, 3.478329e-09, 3.298267e-09, 3.280239e-09, 
    3.247395e-09, 3.163442e-09, 3.094071e-09, 3.237045e-09, 3.076856e-09, 
    3.709136e-09, 3.367201e-09, 3.913649e-09, 3.74285e-09, 3.627372e-09, 
    3.677726e-09, 3.421663e-09, 3.363227e-09, 3.133138e-09, 3.250621e-09, 
    2.596042e-09, 2.872515e-09, 2.15387e-09, 2.339649e-09, 3.911786e-09, 
    3.824555e-09, 3.531788e-09, 3.669004e-09, 3.286499e-09, 3.196934e-09, 
    3.125447e-09, 3.035733e-09, 3.026171e-09, 2.974024e-09, 3.059818e-09, 
    2.977385e-09, 3.297891e-09, 3.151737e-09, 3.564428e-09, 3.460591e-09, 
    3.508091e-09, 3.56072e-09, 3.400094e-09, 3.234754e-09, 3.231311e-09, 
    3.17958e-09, 3.036986e-09, 3.285011e-09, 2.561788e-09, 2.992949e-09, 
    3.731031e-09, 3.569818e-09, 3.547239e-09, 3.608796e-09, 3.205832e-09, 
    3.347878e-09, 2.975291e-09, 3.072873e-09, 2.914178e-09, 2.992273e-09, 
    3.003888e-09, 3.106691e-09, 3.171958e-09, 3.341263e-09, 3.483753e-09, 
    3.599824e-09, 3.572593e-09, 3.445936e-09, 3.224838e-09, 3.025295e-09, 
    3.068216e-09, 2.926026e-09, 3.313221e-09, 3.14661e-09, 3.210263e-09, 
    3.046215e-09, 3.413907e-09, 3.098823e-09, 3.498002e-09, 3.461605e-09, 
    3.350743e-09, 3.135517e-09, 3.08932e-09, 3.040497e-09, 3.070562e-09, 
    3.219367e-09, 3.244244e-09, 3.353413e-09, 3.384003e-09, 3.469508e-09, 
    3.541453e-09, 3.475672e-09, 3.407535e-09, 3.219313e-09, 3.056213e-09, 
    2.885304e-09, 2.844567e-09, 2.655709e-09, 2.8087e-09, 2.559517e-09, 
    2.770246e-09, 2.413057e-09, 3.08127e-09, 2.776673e-09, 3.345769e-09, 
    3.280741e-09, 3.165421e-09, 2.912075e-09, 3.046972e-09, 2.889659e-09, 
    3.245223e-09, 3.441611e-09, 3.493818e-09, 3.592685e-09, 3.491581e-09, 
    3.499727e-09, 3.404752e-09, 3.435069e-09, 3.213196e-09, 3.331049e-09, 
    3.004174e-09, 2.890883e-09, 2.587716e-09, 2.413716e-09, 2.245568e-09, 
    2.174122e-09, 2.152713e-09, 2.143808e-09,
  3.553785e-11, 3.277706e-11, 3.330075e-11, 3.116849e-11, 3.233831e-11, 
    3.096093e-11, 3.496466e-11, 3.267078e-11, 3.41217e-11, 3.528259e-11, 
    2.732496e-11, 3.107586e-11, 2.38018e-11, 2.592189e-11, 2.084808e-11, 
    2.412266e-11, 2.023076e-11, 2.093778e-11, 1.886499e-11, 1.944221e-11, 
    1.696436e-11, 1.8603e-11, 1.577828e-11, 1.734546e-11, 1.709278e-11, 
    1.865898e-11, 3.029191e-11, 2.777222e-11, 3.044635e-11, 3.007552e-11, 
    3.024156e-11, 3.231371e-11, 3.339732e-11, 3.575603e-11, 3.531886e-11, 
    3.359095e-11, 2.990989e-11, 3.112373e-11, 2.813378e-11, 2.819882e-11, 
    2.512476e-11, 2.647772e-11, 2.169867e-11, 2.298461e-11, 1.941786e-11, 
    2.02724e-11, 1.945734e-11, 1.970185e-11, 1.945417e-11, 2.071882e-11, 
    2.01696e-11, 2.130977e-11, 2.62202e-11, 2.469678e-11, 2.944846e-11, 
    3.261809e-11, 3.486153e-11, 3.652217e-11, 3.628387e-11, 3.583276e-11, 
    3.358102e-11, 3.156281e-11, 3.008705e-11, 2.912924e-11, 2.820817e-11, 
    2.555278e-11, 2.422657e-11, 2.144528e-11, 2.192861e-11, 2.111472e-11, 
    2.035895e-11, 1.9136e-11, 1.93334e-11, 1.880847e-11, 2.113604e-11, 
    1.956628e-11, 2.220753e-11, 2.145989e-11, 2.796067e-11, 3.079272e-11, 
    3.205878e-11, 3.319956e-11, 3.610142e-11, 3.407793e-11, 3.486512e-11, 
    3.301457e-11, 3.187757e-11, 3.243621e-11, 2.910338e-11, 3.036682e-11, 
    2.414963e-11, 2.669651e-11, 2.044604e-11, 2.182876e-11, 2.01247e-11, 
    2.098122e-11, 1.952991e-11, 2.083252e-11, 1.861593e-11, 1.815782e-11, 
    1.846993e-11, 1.729295e-11, 2.090658e-11, 1.945727e-11, 3.245192e-11, 
    3.236027e-11, 3.193598e-11, 3.383274e-11, 3.395152e-11, 3.576802e-11, 
    3.414832e-11, 3.34755e-11, 3.181266e-11, 3.085861e-11, 2.997188e-11, 
    2.808975e-11, 2.609436e-11, 2.348583e-11, 2.173704e-11, 2.062106e-11, 
    2.130014e-11, 2.069974e-11, 2.137175e-11, 2.169236e-11, 1.832842e-11, 
    2.016449e-11, 1.745865e-11, 1.760079e-11, 1.879609e-11, 1.758473e-11, 
    3.229605e-11, 3.28253e-11, 3.471323e-11, 3.322903e-11, 3.597017e-11, 
    3.441557e-11, 3.35448e-11, 3.033979e-11, 2.96679e-11, 2.905464e-11, 
    2.787176e-11, 2.640716e-11, 2.397886e-11, 2.200667e-11, 2.031565e-11, 
    2.043612e-11, 2.039364e-11, 2.002856e-11, 2.094195e-11, 1.988154e-11, 
    1.970755e-11, 2.01648e-11, 1.761988e-11, 1.832063e-11, 1.760381e-11, 
    1.805743e-11, 3.265259e-11, 3.176932e-11, 3.224432e-11, 3.135542e-11, 
    3.197963e-11, 2.927379e-11, 2.849719e-11, 2.506765e-11, 2.643537e-11, 
    2.42844e-11, 2.621063e-11, 2.586115e-11, 2.421618e-11, 2.610375e-11, 
    2.211195e-11, 2.476315e-11, 2.001447e-11, 2.24723e-11, 1.986751e-11, 
    2.032275e-11, 1.95733e-11, 1.891991e-11, 1.812159e-11, 1.671549e-11, 
    1.703351e-11, 1.590633e-11, 3.048617e-11, 2.940168e-11, 2.949616e-11, 
    2.839005e-11, 2.759229e-11, 2.592145e-11, 2.340211e-11, 2.432681e-11, 
    2.264994e-11, 2.232405e-11, 2.488007e-11, 2.328585e-11, 2.869242e-11, 
    2.776047e-11, 2.831269e-11, 3.039943e-11, 2.41111e-11, 2.720111e-11, 
    2.170896e-11, 2.322429e-11, 1.901203e-11, 2.102722e-11, 1.721049e-11, 
    1.574919e-11, 1.446201e-11, 1.305985e-11, 2.882239e-11, 2.954516e-11, 
    2.826067e-11, 2.65531e-11, 2.503985e-11, 2.312961e-11, 2.294065e-11, 
    2.259747e-11, 2.172674e-11, 2.101438e-11, 2.248962e-11, 2.083861e-11, 
    2.754728e-11, 2.385605e-11, 2.982177e-11, 2.791887e-11, 2.665162e-11, 
    2.720224e-11, 2.443426e-11, 2.3814e-11, 2.141476e-11, 2.263111e-11, 
    1.610067e-11, 1.878384e-11, 1.20635e-11, 1.371943e-11, 2.980084e-11, 
    2.882495e-11, 2.561483e-11, 2.710665e-11, 2.300621e-11, 2.207299e-11, 
    2.133577e-11, 2.042039e-11, 2.032348e-11, 1.979722e-11, 2.066505e-11, 
    1.983102e-11, 2.312567e-11, 2.160609e-11, 2.596762e-11, 2.484985e-11, 
    2.535952e-11, 2.592747e-11, 2.420482e-11, 2.246577e-11, 2.242992e-11, 
    2.18934e-11, 2.043314e-11, 2.299062e-11, 1.577641e-11, 1.998781e-11, 
    2.778841e-11, 2.602602e-11, 2.578167e-11, 2.644926e-11, 2.216523e-11, 
    2.365181e-11, 1.980996e-11, 2.0798e-11, 1.919798e-11, 1.998095e-11, 
    2.009814e-11, 2.114348e-11, 2.181464e-11, 2.3582e-11, 2.509803e-11, 
    2.635167e-11, 2.605607e-11, 2.469318e-11, 2.236261e-11, 2.031461e-11, 
    2.075056e-11, 1.931621e-11, 2.328668e-11, 2.155331e-11, 2.22112e-11, 
    2.052678e-11, 2.435169e-11, 2.1063e-11, 2.525103e-11, 2.48607e-11, 
    2.368206e-11, 2.143921e-11, 2.096583e-11, 2.046872e-11, 2.077445e-11, 
    2.230574e-11, 2.256462e-11, 2.371026e-11, 2.403403e-11, 2.494531e-11, 
    2.571916e-11, 2.501136e-11, 2.428391e-11, 2.230518e-11, 2.062839e-11, 
    1.89107e-11, 1.850741e-11, 1.666993e-11, 1.815438e-11, 1.575498e-11, 
    1.777798e-11, 1.439018e-11, 2.088366e-11, 1.784072e-11, 2.362953e-11, 
    2.29459e-11, 2.174717e-11, 1.917703e-11, 2.053447e-11, 1.895395e-11, 
    2.257483e-11, 2.4647e-11, 2.520607e-11, 2.627408e-11, 2.518205e-11, 
    2.526957e-11, 2.425431e-11, 2.457716e-11, 2.224164e-11, 2.347431e-11, 
    2.010103e-11, 1.896612e-11, 1.602166e-11, 1.439623e-11, 1.287324e-11, 
    1.224104e-11, 1.205337e-11, 1.197556e-11,
  4.488108e-14, 3.797916e-14, 3.925928e-14, 3.413617e-14, 3.691747e-14, 
    3.365031e-14, 4.341745e-14, 3.772108e-14, 4.129379e-14, 4.422734e-14, 
    2.553412e-14, 3.391904e-14, 1.844821e-14, 2.261447e-14, 1.318213e-14, 
    1.905897e-14, 1.216764e-14, 1.333211e-14, 1.003749e-14, 1.091808e-14, 
    7.353243e-15, 9.647567e-15, 5.856841e-15, 7.863999e-15, 7.523763e-15, 
    9.730375e-15, 3.210029e-14, 2.649063e-14, 3.24559e-14, 3.160424e-14, 
    3.198461e-14, 3.685826e-14, 3.949688e-14, 4.544227e-14, 4.432002e-14, 
    3.997463e-14, 3.122633e-14, 3.403117e-14, 2.727261e-14, 2.741412e-14, 
    2.101234e-14, 2.375612e-14, 1.46303e-14, 1.692585e-14, 1.088034e-14, 
    1.223507e-14, 1.094157e-14, 1.132366e-14, 1.093665e-14, 1.296711e-14, 
    1.206883e-14, 1.396105e-14, 2.322472e-14, 2.016968e-14, 3.018166e-14, 
    3.75934e-14, 4.315579e-14, 4.743062e-14, 4.680923e-14, 4.564018e-14, 
    3.995009e-14, 3.506556e-14, 3.163058e-14, 2.946604e-14, 2.743451e-14, 
    2.186744e-14, 1.92583e-14, 1.419291e-14, 1.503154e-14, 1.36299e-14, 
    1.237571e-14, 1.044729e-14, 1.074985e-14, 9.952853e-15, 1.366593e-14, 
    1.111118e-14, 1.552369e-14, 1.421798e-14, 2.689728e-14, 3.325826e-14, 
    3.624638e-14, 3.901085e-14, 4.633527e-14, 4.11845e-14, 4.316492e-14, 
    3.855799e-14, 3.581339e-14, 3.71535e-14, 2.940832e-14, 3.227261e-14, 
    1.911063e-14, 2.421096e-14, 1.251784e-14, 1.48568e-14, 1.19965e-14, 
    1.340497e-14, 1.105444e-14, 1.315616e-14, 9.666678e-15, 8.999314e-15, 
    9.451905e-15, 7.792776e-15, 1.327986e-14, 1.094147e-14, 3.719143e-14, 
    3.697039e-14, 3.595274e-14, 4.057387e-14, 4.08693e-14, 4.547318e-14, 
    4.136033e-14, 3.968952e-14, 3.565873e-14, 3.341166e-14, 3.136756e-14, 
    2.717697e-14, 2.296661e-14, 1.785387e-14, 1.469696e-14, 1.280539e-14, 
    1.394463e-14, 1.293548e-14, 1.40669e-14, 1.461933e-14, 9.24559e-15, 
    1.206059e-14, 8.018409e-15, 8.214065e-15, 9.934358e-15, 8.191863e-15, 
    3.681575e-14, 3.809648e-14, 4.278043e-14, 3.908311e-14, 4.599526e-14, 
    4.203023e-14, 3.986059e-14, 3.22104e-14, 3.067693e-14, 2.929966e-14, 
    2.670505e-14, 2.36101e-14, 1.878433e-14, 1.516868e-14, 1.230526e-14, 
    1.250162e-14, 1.243225e-14, 1.184219e-14, 1.33391e-14, 1.160773e-14, 
    1.133264e-14, 1.206108e-14, 8.240502e-15, 9.234273e-15, 8.218258e-15, 
    8.855635e-15, 3.767692e-14, 3.55556e-14, 3.669135e-14, 3.457571e-14, 
    3.605701e-14, 2.978938e-14, 2.806663e-14, 2.089922e-14, 2.366845e-14, 
    1.936956e-14, 2.320505e-14, 2.249092e-14, 1.923836e-14, 2.298579e-14, 
    1.535441e-14, 2.029959e-14, 1.181964e-14, 1.599643e-14, 1.158546e-14, 
    1.23168e-14, 1.112214e-14, 1.012002e-14, 8.947353e-15, 7.027411e-15, 
    7.444849e-15, 6.011403e-15, 3.25478e-14, 3.007642e-14, 3.028906e-14, 
    2.78317e-14, 2.610427e-14, 2.261357e-14, 1.76976e-14, 1.945128e-14, 
    1.631645e-14, 1.573107e-14, 2.052904e-14, 1.748143e-14, 2.849638e-14, 
    2.646527e-14, 2.766252e-14, 3.234773e-14, 1.903683e-14, 2.527136e-14, 
    1.464817e-14, 1.736735e-14, 1.025903e-14, 1.348234e-14, 7.681476e-15, 
    5.821982e-15, 4.370629e-15, 3.004993e-15, 2.878373e-14, 3.039956e-14, 
    2.754895e-14, 2.39125e-14, 2.084418e-14, 1.719245e-14, 1.684533e-14, 
    1.622167e-14, 1.467905e-14, 1.34607e-14, 1.602751e-14, 1.316631e-14, 
    2.600802e-14, 1.855095e-14, 3.102589e-14, 2.680683e-14, 2.411738e-14, 
    2.527374e-14, 1.965895e-14, 1.847126e-14, 1.414057e-14, 1.628241e-14, 
    6.249308e-15, 9.916089e-15, 2.180953e-15, 3.618328e-15, 3.097832e-14, 
    2.878937e-14, 2.199237e-14, 2.507162e-14, 1.696548e-14, 1.528557e-14, 
    1.400541e-14, 1.247593e-14, 1.231798e-14, 1.14741e-14, 1.287806e-14, 
    1.152759e-14, 1.718518e-14, 1.44699e-14, 2.270762e-14, 2.046964e-14, 
    2.14798e-14, 2.262581e-14, 1.921647e-14, 1.598469e-14, 1.592037e-14, 
    1.496984e-14, 1.249684e-14, 1.693688e-14, 5.854638e-15, 1.177709e-14, 
    2.652538e-14, 2.282686e-14, 2.232961e-14, 2.369717e-14, 1.544869e-14, 
    1.816517e-14, 1.149424e-14, 1.309865e-14, 1.054192e-14, 1.176607e-14, 
    1.195379e-14, 1.367853e-14, 1.483215e-14, 1.8034e-14, 2.095936e-14, 
    2.349547e-14, 2.288823e-14, 2.016264e-14, 1.579993e-14, 1.230358e-14, 
    1.301978e-14, 1.072337e-14, 1.748295e-14, 1.437876e-14, 1.553024e-14, 
    1.265018e-14, 1.949931e-14, 1.354266e-14, 2.126331e-14, 2.049095e-14, 
    1.822212e-14, 1.418251e-14, 1.337915e-14, 1.255498e-14, 1.305947e-14, 
    1.569842e-14, 1.616244e-14, 1.827526e-14, 1.888951e-14, 2.065751e-14, 
    2.220301e-14, 2.078785e-14, 1.93686e-14, 1.569741e-14, 1.281749e-14, 
    1.010616e-14, 9.506854e-15, 6.968465e-15, 8.994401e-15, 5.828946e-15, 
    8.460761e-15, 4.295109e-15, 1.324157e-14, 8.54876e-15, 1.812327e-14, 
    1.685495e-14, 1.47146e-14, 1.050993e-14, 1.266281e-14, 1.017132e-14, 
    1.618083e-14, 2.007249e-14, 2.117383e-14, 2.333555e-14, 2.112606e-14, 
    2.130026e-14, 1.931161e-14, 1.993636e-14, 1.558431e-14, 1.783233e-14, 
    1.195844e-14, 1.018967e-14, 6.152106e-15, 4.301424e-15, 2.841109e-15, 
    2.318504e-15, 2.173228e-15, 2.114337e-15,
  1.518248e-19, 1.28757e-19, 1.330399e-19, 1.158864e-19, 1.252033e-19, 
    1.142577e-19, 1.469378e-19, 1.278933e-19, 1.398425e-19, 1.496423e-19, 
    8.699569e-20, 1.151586e-19, 6.309223e-20, 7.715978e-20, 4.524835e-20, 
    6.515706e-20, 4.180048e-20, 4.575776e-20, 3.454754e-20, 3.754819e-20, 
    2.537725e-20, 3.321771e-20, 2.024644e-20, 2.71252e-20, 2.596099e-20, 
    3.350018e-20, 1.090595e-19, 9.021444e-20, 1.102524e-19, 1.073951e-19, 
    1.086714e-19, 1.250051e-19, 1.338346e-19, 1.53698e-19, 1.499517e-19, 
    1.354323e-19, 1.061269e-19, 1.155344e-19, 9.284465e-20, 9.332052e-20, 
    7.175487e-20, 8.100791e-20, 5.016379e-20, 5.794173e-20, 3.741965e-20, 
    4.202974e-20, 3.762816e-20, 3.892908e-20, 3.76114e-20, 4.451787e-20, 
    4.146443e-20, 4.789308e-20, 7.921706e-20, 6.890975e-20, 1.026199e-19, 
    1.27466e-19, 1.460638e-19, 1.60332e-19, 1.582592e-19, 1.543585e-19, 
    1.353503e-19, 1.190009e-19, 1.074835e-19, 1.002165e-19, 9.338907e-20, 
    7.464031e-20, 6.583076e-20, 4.867992e-20, 5.152446e-20, 4.676895e-20, 
    4.250792e-20, 3.594436e-20, 3.697519e-20, 3.425894e-20, 4.689129e-20, 
    3.820572e-20, 5.319275e-20, 4.876501e-20, 9.158235e-20, 1.129433e-19, 
    1.229562e-19, 1.322089e-19, 1.566779e-19, 1.394772e-19, 1.460943e-19, 
    1.306939e-19, 1.215061e-19, 1.259935e-19, 1.000226e-19, 1.096376e-19, 
    6.533165e-20, 8.254024e-20, 4.299109e-20, 5.093195e-20, 4.121845e-20, 
    4.600519e-20, 3.801254e-20, 4.516011e-20, 3.328291e-20, 3.100526e-20, 
    3.255015e-20, 2.688155e-20, 4.55803e-20, 3.762783e-20, 1.261205e-19, 
    1.253805e-19, 1.219728e-19, 1.374359e-19, 1.384236e-19, 1.538011e-19, 
    1.400649e-19, 1.344789e-19, 1.209881e-19, 1.134576e-19, 1.066009e-19, 
    9.252301e-20, 7.834702e-20, 6.108199e-20, 5.03899e-20, 4.396839e-20, 
    4.783734e-20, 4.441042e-20, 4.825233e-20, 5.012659e-20, 3.184603e-20, 
    4.143641e-20, 2.765333e-20, 2.832234e-20, 3.419587e-20, 2.824644e-20, 
    1.248628e-19, 1.291496e-19, 1.4481e-19, 1.324506e-19, 1.555434e-19, 
    1.423036e-19, 1.35051e-19, 1.094289e-19, 1.042828e-19, 9.965765e-20, 
    9.093576e-20, 8.051587e-20, 6.422867e-20, 5.198944e-20, 4.226843e-20, 
    4.293597e-20, 4.270014e-20, 4.069356e-20, 4.578147e-20, 3.989586e-20, 
    3.895965e-20, 4.143809e-20, 2.841272e-20, 3.18074e-20, 2.833667e-20, 
    3.051461e-20, 1.277455e-19, 1.206426e-19, 1.244462e-19, 1.173595e-19, 
    1.223221e-19, 1.013026e-19, 9.551425e-20, 7.137301e-20, 8.071248e-20, 
    6.620674e-20, 7.915075e-20, 7.674318e-20, 6.576338e-20, 7.841169e-20, 
    5.261901e-20, 6.934848e-20, 4.061686e-20, 5.47945e-20, 3.982006e-20, 
    4.230763e-20, 3.824303e-20, 3.482888e-20, 3.082783e-20, 2.426133e-20, 
    2.569087e-20, 2.077713e-20, 1.105606e-19, 1.022665e-19, 1.029805e-19, 
    9.472449e-20, 8.891452e-20, 7.715674e-20, 6.055328e-20, 6.648289e-20, 
    5.587846e-20, 5.389547e-20, 7.012328e-20, 5.982184e-20, 9.695863e-20, 
    9.012913e-20, 9.41557e-20, 1.098896e-19, 6.508224e-20, 8.61112e-20, 
    5.022439e-20, 5.943584e-20, 3.530276e-20, 4.626793e-20, 2.650074e-20, 
    2.012672e-20, 1.513347e-20, 1.041586e-20, 9.792425e-20, 1.033516e-19, 
    9.377386e-20, 8.15348e-20, 7.118723e-20, 5.884402e-20, 5.766916e-20, 
    5.555746e-20, 5.032915e-20, 4.619445e-20, 5.48998e-20, 4.519461e-20, 
    8.859064e-20, 6.343964e-20, 1.054541e-19, 9.127813e-20, 8.222503e-20, 
    8.61192e-20, 6.718457e-20, 6.317016e-20, 4.850233e-20, 5.576317e-20, 
    2.159362e-20, 3.413357e-20, 7.557001e-21, 1.253726e-20, 1.052945e-19, 
    9.794322e-20, 7.506176e-20, 8.543874e-20, 5.807583e-20, 5.238565e-20, 
    4.804365e-20, 4.284863e-20, 4.231166e-20, 3.94411e-20, 4.421532e-20, 
    3.962315e-20, 5.881941e-20, 4.961971e-20, 7.747387e-20, 6.992271e-20, 
    7.333246e-20, 7.719803e-20, 6.568939e-20, 5.475473e-20, 5.453684e-20, 
    5.131527e-20, 4.29197e-20, 5.797904e-20, 2.023887e-20, 4.047208e-20, 
    9.033135e-20, 7.787588e-20, 7.619921e-20, 8.080926e-20, 5.293856e-20, 
    6.2135e-20, 3.950964e-20, 4.496476e-20, 3.626683e-20, 4.043459e-20, 
    4.107316e-20, 4.693406e-20, 5.084838e-20, 6.169132e-20, 7.157604e-20, 
    8.012956e-20, 7.808279e-20, 6.888597e-20, 5.41288e-20, 4.226271e-20, 
    4.469683e-20, 3.688497e-20, 5.982696e-20, 4.931053e-20, 5.321494e-20, 
    4.344091e-20, 6.664518e-20, 4.647276e-20, 7.260191e-20, 6.999469e-20, 
    6.232762e-20, 4.864466e-20, 4.591749e-20, 4.311734e-20, 4.483166e-20, 
    5.378487e-20, 5.535683e-20, 6.250734e-20, 6.458426e-20, 7.055702e-20, 
    7.577224e-20, 7.099708e-20, 6.62035e-20, 5.378144e-20, 4.400952e-20, 
    3.478164e-20, 3.273764e-20, 2.405938e-20, 3.098848e-20, 2.015064e-20, 
    2.916557e-20, 1.487312e-20, 4.545022e-20, 2.946628e-20, 6.199328e-20, 
    5.770171e-20, 5.044972e-20, 3.615781e-20, 4.348384e-20, 3.500378e-20, 
    5.541914e-20, 6.858152e-20, 7.229992e-20, 7.959061e-20, 7.213871e-20, 
    7.27266e-20, 6.60109e-20, 6.812171e-20, 5.339817e-20, 6.100909e-20, 
    4.108898e-20, 3.506632e-20, 2.126007e-20, 1.48949e-20, 9.848162e-21, 
    8.035011e-21, 7.530147e-21, 7.325373e-21,
  1.114744e-25, 9.461627e-26, 9.774716e-26, 8.520466e-26, 9.201808e-26, 
    8.401338e-26, 1.079039e-25, 9.398483e-26, 1.027191e-25, 1.098799e-25, 
    6.406004e-26, 8.467233e-26, 4.653991e-26, 5.685412e-26, 3.343759e-26, 
    4.805451e-26, 3.090297e-26, 3.381198e-26, 2.556723e-26, 2.77754e-26, 
    1.881149e-26, 2.458828e-26, 1.502547e-26, 2.010018e-26, 1.924192e-26, 
    2.479624e-26, 8.021063e-26, 6.641725e-26, 8.108338e-26, 7.89929e-26, 
    7.992668e-26, 9.187313e-26, 9.832805e-26, 1.128429e-25, 1.10106e-25, 
    9.949588e-26, 7.806494e-26, 8.494724e-26, 6.834315e-26, 6.869157e-26, 
    5.289253e-26, 5.967382e-26, 3.70493e-26, 4.276053e-26, 2.768083e-26, 
    3.107154e-26, 2.783423e-26, 2.879125e-26, 2.78219e-26, 3.290069e-26, 
    3.065587e-26, 3.53811e-26, 5.836167e-26, 5.080656e-26, 7.549863e-26, 
    9.367238e-26, 1.072654e-25, 1.176887e-25, 1.161747e-25, 1.133254e-25, 
    9.943592e-26, 8.748255e-26, 7.905756e-26, 7.373967e-26, 6.874175e-26, 
    5.500763e-26, 4.854862e-26, 3.59592e-26, 3.804873e-26, 3.455509e-26, 
    3.142312e-26, 2.659528e-26, 2.735381e-26, 2.53548e-26, 3.464499e-26, 
    2.825914e-26, 3.927393e-26, 3.602172e-26, 6.74189e-26, 8.305187e-26, 
    9.037501e-26, 9.713971e-26, 1.150197e-25, 1.024521e-25, 1.072876e-25, 
    9.60322e-26, 8.931462e-26, 9.259583e-26, 7.359776e-26, 8.063355e-26, 
    4.818256e-26, 6.079644e-26, 3.177834e-26, 3.761354e-26, 3.047499e-26, 
    3.399383e-26, 2.811702e-26, 3.337274e-26, 2.463628e-26, 2.295906e-26, 
    2.409676e-26, 1.992058e-26, 3.368156e-26, 2.783399e-26, 9.268865e-26, 
    9.214761e-26, 8.96559e-26, 1.009603e-25, 1.016821e-25, 1.129182e-25, 
    1.028816e-25, 9.879899e-26, 8.893578e-26, 8.342809e-26, 7.841176e-26, 
    6.810766e-26, 5.772414e-26, 4.506511e-26, 3.721539e-26, 3.249678e-26, 
    3.534014e-26, 3.28217e-26, 3.564505e-26, 3.702197e-26, 2.357827e-26, 
    3.063526e-26, 2.048945e-26, 2.09825e-26, 2.530837e-26, 2.092656e-26, 
    9.176907e-26, 9.490328e-26, 1.063492e-25, 9.731641e-26, 1.14191e-25, 
    1.045177e-25, 9.921716e-26, 8.048087e-26, 7.671552e-26, 7.333061e-26, 
    6.694545e-26, 5.931332e-26, 4.737355e-26, 3.839023e-26, 3.124704e-26, 
    3.173782e-26, 3.156444e-26, 3.0089e-26, 3.382941e-26, 2.950234e-26, 
    2.881374e-26, 3.06365e-26, 2.10491e-26, 2.354982e-26, 2.099306e-26, 
    2.259766e-26, 9.387677e-26, 8.868316e-26, 9.146451e-26, 8.628209e-26, 
    8.991127e-26, 7.453453e-26, 7.029763e-26, 5.261258e-26, 5.945738e-26, 
    4.882437e-26, 5.831309e-26, 5.654883e-26, 4.849921e-26, 5.777153e-26, 
    3.885259e-26, 5.112824e-26, 3.00326e-26, 4.045007e-26, 2.94466e-26, 
    3.127586e-26, 2.828658e-26, 2.577432e-26, 2.282838e-26, 1.798849e-26, 
    1.904275e-26, 1.541732e-26, 8.130888e-26, 7.524001e-26, 7.576254e-26, 
    6.971946e-26, 6.546532e-26, 5.68519e-26, 4.467718e-26, 4.90269e-26, 
    4.124591e-26, 3.978995e-26, 5.169634e-26, 4.414046e-26, 7.135499e-26, 
    6.635478e-26, 6.930304e-26, 8.081792e-26, 4.799963e-26, 6.341222e-26, 
    3.709381e-26, 4.385717e-26, 2.61231e-26, 3.418691e-26, 1.963985e-26, 
    1.493707e-26, 1.124652e-26, 7.752129e-27, 7.206183e-26, 7.603406e-26, 
    6.902348e-26, 6.005984e-26, 5.247638e-26, 4.342281e-26, 4.256045e-26, 
    4.101024e-26, 3.717076e-26, 3.413291e-26, 4.052739e-26, 3.339809e-26, 
    6.522813e-26, 4.679476e-26, 7.757267e-26, 6.719614e-26, 6.056552e-26, 
    6.341808e-26, 4.954148e-26, 4.659708e-26, 3.582872e-26, 4.116126e-26, 
    1.602008e-26, 2.526251e-26, 5.629368e-27, 9.324627e-27, 7.745584e-26, 
    7.207572e-26, 5.531652e-26, 6.291967e-26, 4.285897e-26, 3.868122e-26, 
    3.549172e-26, 3.167361e-26, 3.127882e-26, 2.916787e-26, 3.26783e-26, 
    2.930177e-26, 4.340474e-26, 3.664962e-26, 5.70843e-26, 5.154928e-26, 
    5.404898e-26, 5.688215e-26, 4.844494e-26, 4.042087e-26, 4.026089e-26, 
    3.789508e-26, 3.172586e-26, 4.278792e-26, 1.501988e-26, 2.992613e-26, 
    6.650286e-26, 5.73789e-26, 5.615016e-26, 5.952828e-26, 3.908726e-26, 
    4.583768e-26, 2.921828e-26, 3.322916e-26, 2.683258e-26, 2.989855e-26, 
    3.036815e-26, 3.467642e-26, 3.755215e-26, 4.551217e-26, 5.276141e-26, 
    5.903028e-26, 5.753052e-26, 5.078912e-26, 3.996128e-26, 3.124283e-26, 
    3.303223e-26, 2.728743e-26, 4.414422e-26, 3.642248e-26, 3.929023e-26, 
    3.210903e-26, 4.914592e-26, 3.433743e-26, 5.351347e-26, 5.160205e-26, 
    4.597899e-26, 3.59333e-26, 3.392938e-26, 3.187116e-26, 3.313133e-26, 
    3.970873e-26, 4.086294e-26, 4.611083e-26, 4.763437e-26, 5.201434e-26, 
    5.583725e-26, 5.233697e-26, 4.8822e-26, 3.970621e-26, 3.252702e-26, 
    2.573954e-26, 2.423482e-26, 1.783953e-26, 2.29467e-26, 1.495473e-26, 
    2.160384e-26, 1.10539e-26, 3.358596e-26, 2.182539e-26, 4.573371e-26, 
    4.258435e-26, 3.725933e-26, 2.675235e-26, 3.214059e-26, 2.590305e-26, 
    4.090868e-26, 5.056588e-26, 5.329209e-26, 5.863538e-26, 5.317391e-26, 
    5.360487e-26, 4.868074e-26, 5.022871e-26, 3.942477e-26, 4.501162e-26, 
    3.037979e-26, 2.594908e-26, 1.577386e-26, 1.107001e-26, 7.330961e-27, 
    5.98464e-27, 5.609405e-27, 5.457159e-27,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.004712567, 0.004712572, 0.004712572, 0.004712573, 0.004712574, 
    0.004712573, 0.00471257, 0.00471257, 0.004712572, 0.00471257, 
    0.004712562, 0.004712573, 0.004712561, 0.004712572, 0.004712542, 
    0.00471256, 0.004712538, 0.004712547, 0.004712529, 0.004712535, 
    0.004712495, 0.004712526, 0.004712479, 0.004712506, 0.0047125, 
    0.004712526, 0.004712576, 0.004712563, 0.004712576, 0.004712574, 
    0.004712576, 0.004712573, 0.004712568, 0.00471257, 0.00471257, 
    0.00471257, 0.004712574, 0.004712576, 0.004712577, 0.004712578, 
    0.00471257, 0.004712575, 0.004712553, 0.004712563, 0.004712535, 
    0.004712542, 0.004712534, 0.004712537, 0.004712534, 0.004712545, 
    0.004712541, 0.004712551, 0.004712573, 0.004712568, 0.004712575, 
    0.004712566, 0.00471257, 0.004712568, 0.004712568, 0.004712568, 
    0.00471257, 0.004712576, 0.004712577, 0.004712577, 0.004712577, 
    0.004712563, 0.004712563, 0.004712549, 0.004712556, 0.004712547, 
    0.004712543, 0.00471253, 0.004712533, 0.004712526, 0.00471255, 
    0.004712533, 0.004712559, 0.004712552, 0.004712562, 0.004712576, 
    0.004712568, 0.004712572, 0.004712568, 0.00471257, 0.004712569, 
    0.004712574, 0.004712575, 0.004712576, 0.004712577, 0.004712577, 
    0.004712563, 0.004712572, 0.004712543, 0.004712555, 0.004712541, 
    0.004712549, 0.004712534, 0.004712548, 0.004712525, 0.004712517, 
    0.004712522, 0.004712508, 0.004712548, 0.004712533, 0.004712575, 
    0.004712575, 0.004712576, 0.00471257, 0.00471257, 0.004712569, 
    0.004712572, 0.004712571, 0.004712577, 0.004712576, 0.004712577, 
    0.004712576, 0.00471257, 0.004712562, 0.004712554, 0.004712546, 
    0.004712552, 0.004712547, 0.004712552, 0.004712555, 0.004712519, 
    0.004712539, 0.00471251, 0.004712513, 0.004712525, 0.004712512, 
    0.004712575, 0.004712575, 0.00471257, 0.004712574, 0.004712569, 
    0.00471257, 0.00471257, 0.004712573, 0.004712577, 0.004712576, 
    0.004712577, 0.004712574, 0.004712564, 0.004712554, 0.004712543, 
    0.004712545, 0.004712544, 0.00471254, 0.004712548, 0.004712539, 
    0.004712536, 0.004712542, 0.004712513, 0.004712522, 0.004712513, 
    0.004712519, 0.004712576, 0.004712576, 0.004712575, 0.004712575, 
    0.004712574, 0.004712573, 0.004712571, 0.004712566, 0.004712573, 
    0.004712565, 0.004712574, 0.004712572, 0.004712558, 0.004712575, 
    0.004712551, 0.004712563, 0.00471254, 0.00471255, 0.004712538, 
    0.004712544, 0.004712536, 0.004712528, 0.004712519, 0.004712496, 
    0.004712502, 0.004712484, 0.004712577, 0.004712575, 0.004712577, 
    0.004712577, 0.004712575, 0.004712574, 0.004712563, 0.004712569, 
    0.004712561, 0.004712558, 0.004712571, 0.004712561, 0.004712575, 
    0.004712571, 0.004712576, 0.004712575, 0.004712563, 0.004712571, 
    0.004712553, 0.004712563, 0.004712529, 0.004712545, 0.004712505, 
    0.004712474, 0.004712456, 0.004712414, 0.004712577, 0.004712578, 
    0.004712578, 0.00471257, 0.00471257, 0.004712562, 0.004712562, 
    0.004712559, 0.004712555, 0.00471255, 0.004712556, 0.004712548, 
    0.004712564, 0.004712563, 0.004712576, 0.004712571, 0.004712572, 
    0.004712575, 0.00471257, 0.004712567, 0.004712549, 0.004712561, 
    0.004712479, 0.004712522, 0.004712389, 0.004712433, 0.004712577, 
    0.004712578, 0.00471257, 0.004712575, 0.004712563, 0.004712556, 
    0.004712552, 0.004712542, 0.004712543, 0.004712537, 0.004712547, 
    0.004712539, 0.004712562, 0.004712553, 0.004712575, 0.00471257, 
    0.004712573, 0.004712575, 0.004712569, 0.004712555, 0.004712559, 
    0.004712553, 0.004712526, 0.004712563, 0.004712464, 0.004712524, 
    0.004712577, 0.004712569, 0.004712573, 0.004712576, 0.004712556, 
    0.004712565, 0.004712538, 0.004712548, 0.004712532, 0.00471254, 
    0.004712541, 0.00471255, 0.004712555, 0.004712563, 0.00471257, 
    0.004712576, 0.004712575, 0.004712568, 0.004712555, 0.004712541, 
    0.004712544, 0.004712534, 0.004712564, 0.00471255, 0.004712555, 
    0.004712544, 0.004712568, 0.004712534, 0.004712573, 0.004712571, 
    0.004712565, 0.004712546, 0.004712549, 0.004712543, 0.004712548, 
    0.004712555, 0.004712558, 0.004712566, 0.004712566, 0.004712572, 
    0.004712575, 0.004712571, 0.004712566, 0.004712557, 0.004712543, 
    0.004712527, 0.004712524, 0.004712487, 0.004712511, 0.004712462, 
    0.004712494, 0.004712441, 0.004712539, 0.004712505, 0.004712566, 
    0.004712563, 0.00471255, 0.004712525, 0.004712544, 0.004712524, 
    0.004712559, 0.004712565, 0.004712573, 0.004712575, 0.004712572, 
    0.004712573, 0.00471257, 0.004712571, 0.004712557, 0.004712565, 
    0.004712539, 0.004712526, 0.004712484, 0.004712449, 0.004712416, 
    0.004712397, 0.004712392, 0.004712389,
  9.379945e-06, 9.388586e-06, 9.386914e-06, 9.393862e-06, 9.390018e-06, 
    9.394558e-06, 9.381709e-06, 9.38892e-06, 9.384325e-06, 9.380738e-06, 
    9.407278e-06, 9.394174e-06, 9.421875e-06, 9.412604e-06, 9.436173e-06, 
    9.420389e-06, 9.439352e-06, 9.435744e-06, 9.446652e-06, 9.443533e-06, 
    9.457394e-06, 9.448092e-06, 9.464598e-06, 9.455189e-06, 9.456653e-06, 
    9.447781e-06, 9.396837e-06, 9.405642e-06, 9.39631e-06, 9.397568e-06, 
    9.397008e-06, 9.390089e-06, 9.386582e-06, 9.379301e-06, 9.380627e-06, 
    9.385984e-06, 9.398134e-06, 9.39403e-06, 9.404413e-06, 9.404179e-06, 
    9.41591e-06, 9.410503e-06, 9.431938e-06, 9.425728e-06, 9.443664e-06, 
    9.439158e-06, 9.443447e-06, 9.44215e-06, 9.443464e-06, 9.436855e-06, 
    9.439687e-06, 9.433874e-06, 9.41147e-06, 9.417816e-06, 9.399741e-06, 
    9.389067e-06, 9.382022e-06, 9.376998e-06, 9.377708e-06, 9.379058e-06, 
    9.386015e-06, 9.392567e-06, 9.397546e-06, 9.40087e-06, 9.404145e-06, 
    9.413979e-06, 9.419927e-06, 9.43318e-06, 9.430812e-06, 9.434839e-06, 
    9.438711e-06, 9.445173e-06, 9.444112e-06, 9.446951e-06, 9.434748e-06, 
    9.442855e-06, 9.429459e-06, 9.433125e-06, 9.404954e-06, 9.395141e-06, 
    9.390893e-06, 9.387232e-06, 9.378253e-06, 9.384452e-06, 9.382007e-06, 
    9.387837e-06, 9.391527e-06, 9.389706e-06, 9.400961e-06, 9.396585e-06, 
    9.42028e-06, 9.409669e-06, 9.438259e-06, 9.431301e-06, 9.439927e-06, 
    9.435533e-06, 9.443053e-06, 9.436286e-06, 9.448014e-06, 9.450553e-06, 
    9.448816e-06, 9.455511e-06, 9.435907e-06, 9.443439e-06, 9.389651e-06, 
    9.389947e-06, 9.391339e-06, 9.38522e-06, 9.38485e-06, 9.379261e-06, 
    9.384242e-06, 9.386355e-06, 9.391747e-06, 9.394917e-06, 9.397935e-06, 
    9.404563e-06, 9.411937e-06, 9.423355e-06, 9.431751e-06, 9.437365e-06, 
    9.433929e-06, 9.436963e-06, 9.433568e-06, 9.43198e-06, 9.449596e-06, 
    9.439708e-06, 9.454548e-06, 9.453733e-06, 9.447015e-06, 9.453825e-06, 
    9.390157e-06, 9.388447e-06, 9.382482e-06, 9.387151e-06, 9.378652e-06, 
    9.383401e-06, 9.386124e-06, 9.396659e-06, 9.39899e-06, 9.401125e-06, 
    9.405356e-06, 9.410768e-06, 9.421076e-06, 9.430419e-06, 9.438939e-06, 
    9.438317e-06, 9.438535e-06, 9.440427e-06, 9.435727e-06, 9.441199e-06, 
    9.442108e-06, 9.439717e-06, 9.453623e-06, 9.449656e-06, 9.453714e-06, 
    9.451135e-06, 9.389006e-06, 9.391884e-06, 9.390328e-06, 9.39325e-06, 
    9.391185e-06, 9.400337e-06, 9.403077e-06, 9.416142e-06, 9.410657e-06, 
    9.419676e-06, 9.411513e-06, 9.412837e-06, 9.419949e-06, 9.411923e-06, 
    9.429888e-06, 9.417491e-06, 9.4405e-06, 9.428123e-06, 9.441273e-06, 
    9.438902e-06, 9.442835e-06, 9.446345e-06, 9.45077e-06, 9.458897e-06, 
    9.45702e-06, 9.463818e-06, 9.396181e-06, 9.399901e-06, 9.399589e-06, 
    9.403489e-06, 9.406367e-06, 9.412617e-06, 9.423756e-06, 9.419503e-06, 
    9.427324e-06, 9.428886e-06, 9.417013e-06, 9.424292e-06, 9.4024e-06, 
    9.405732e-06, 9.40376e-06, 9.396465e-06, 9.420462e-06, 9.407783e-06, 
    9.431887e-06, 9.424592e-06, 9.445842e-06, 9.435274e-06, 9.455983e-06, 
    9.464755e-06, 9.473065e-06, 9.48266e-06, 9.401946e-06, 9.399419e-06, 
    9.403956e-06, 9.410198e-06, 9.41629e-06, 9.425035e-06, 9.425938e-06, 
    9.427568e-06, 9.431809e-06, 9.435364e-06, 9.428069e-06, 9.436256e-06, 
    9.406474e-06, 9.42164e-06, 9.398448e-06, 9.405153e-06, 9.409837e-06, 
    9.407799e-06, 9.419021e-06, 9.421853e-06, 9.433336e-06, 9.427415e-06, 
    9.462578e-06, 9.447062e-06, 9.490002e-06, 9.478049e-06, 9.398531e-06, 
    9.401944e-06, 9.413777e-06, 9.408154e-06, 9.425627e-06, 9.430103e-06, 
    9.433751e-06, 9.438384e-06, 9.438895e-06, 9.441639e-06, 9.43714e-06, 
    9.441467e-06, 9.425054e-06, 9.4324e-06, 9.412445e-06, 9.417138e-06, 
    9.414885e-06, 9.412598e-06, 9.420061e-06, 9.42818e-06, 9.428379e-06, 
    9.430973e-06, 9.438229e-06, 9.425701e-06, 9.464527e-06, 9.440557e-06, 
    9.405661e-06, 9.412187e-06, 9.413148e-06, 9.410617e-06, 9.429654e-06, 
    9.422596e-06, 9.441575e-06, 9.436461e-06, 9.444844e-06, 9.440679e-06, 
    9.440065e-06, 9.434712e-06, 9.43137e-06, 9.422915e-06, 9.416029e-06, 
    9.410987e-06, 9.412107e-06, 9.417836e-06, 9.428682e-06, 9.438931e-06, 
    9.436684e-06, 9.444208e-06, 9.424304e-06, 9.432651e-06, 9.429418e-06, 
    9.437844e-06, 9.419384e-06, 9.435033e-06, 9.415365e-06, 9.417098e-06, 
    9.422456e-06, 9.433198e-06, 9.435609e-06, 9.438135e-06, 9.436581e-06, 
    9.428962e-06, 9.427723e-06, 9.422332e-06, 9.42083e-06, 9.416723e-06, 
    9.413397e-06, 9.416422e-06, 9.419684e-06, 9.428975e-06, 9.437314e-06, 
    9.44639e-06, 9.448619e-06, 9.459122e-06, 9.450539e-06, 9.464656e-06, 
    9.452604e-06, 9.473465e-06, 9.435975e-06, 9.452301e-06, 9.422708e-06, 
    9.425915e-06, 9.431679e-06, 9.44492e-06, 9.437805e-06, 9.446137e-06, 
    9.427677e-06, 9.41803e-06, 9.415561e-06, 9.411275e-06, 9.415668e-06, 
    9.415281e-06, 9.419838e-06, 9.418375e-06, 9.429284e-06, 9.423429e-06, 
    9.440042e-06, 9.446077e-06, 9.463097e-06, 9.473471e-06, 9.484038e-06, 
    9.488677e-06, 9.490091e-06, 9.49068e-06,
  1.936e-10, 1.938759e-10, 1.938224e-10, 1.940449e-10, 1.939217e-10, 
    1.940672e-10, 1.936562e-10, 1.938866e-10, 1.937397e-10, 1.936253e-10, 
    1.944769e-10, 1.940549e-10, 1.949454e-10, 1.946491e-10, 1.954033e-10, 
    1.94898e-10, 1.955055e-10, 1.953895e-10, 1.957406e-10, 1.9564e-10, 
    1.96088e-10, 1.957871e-10, 1.963219e-10, 1.960166e-10, 1.96064e-10, 
    1.95777e-10, 1.941404e-10, 1.94424e-10, 1.941235e-10, 1.941639e-10, 
    1.941459e-10, 1.93924e-10, 1.938118e-10, 1.935795e-10, 1.936218e-10, 
    1.937927e-10, 1.941821e-10, 1.940503e-10, 1.943843e-10, 1.943768e-10, 
    1.947552e-10, 1.945811e-10, 1.952674e-10, 1.950686e-10, 1.956443e-10, 
    1.954992e-10, 1.956373e-10, 1.955955e-10, 1.956379e-10, 1.954252e-10, 
    1.955163e-10, 1.953295e-10, 1.946124e-10, 1.948159e-10, 1.942338e-10, 
    1.938913e-10, 1.936662e-10, 1.935062e-10, 1.935288e-10, 1.935717e-10, 
    1.937937e-10, 1.940034e-10, 1.941632e-10, 1.942701e-10, 1.943757e-10, 
    1.946937e-10, 1.948832e-10, 1.953072e-10, 1.952313e-10, 1.953604e-10, 
    1.954848e-10, 1.956929e-10, 1.956587e-10, 1.957503e-10, 1.953575e-10, 
    1.956182e-10, 1.951879e-10, 1.953055e-10, 1.944018e-10, 1.94086e-10, 
    1.939497e-10, 1.938326e-10, 1.935461e-10, 1.937437e-10, 1.936657e-10, 
    1.938519e-10, 1.9397e-10, 1.939117e-10, 1.942731e-10, 1.941323e-10, 
    1.948945e-10, 1.945541e-10, 1.954703e-10, 1.95247e-10, 1.95524e-10, 
    1.953827e-10, 1.956246e-10, 1.954069e-10, 1.957846e-10, 1.958666e-10, 
    1.958105e-10, 1.96027e-10, 1.953948e-10, 1.95637e-10, 1.9391e-10, 
    1.939194e-10, 1.93964e-10, 1.937683e-10, 1.937565e-10, 1.935782e-10, 
    1.93737e-10, 1.938045e-10, 1.939771e-10, 1.940788e-10, 1.941757e-10, 
    1.943892e-10, 1.946275e-10, 1.949927e-10, 1.952614e-10, 1.954416e-10, 
    1.953313e-10, 1.954286e-10, 1.953197e-10, 1.952687e-10, 1.958357e-10, 
    1.955169e-10, 1.959958e-10, 1.959694e-10, 1.957524e-10, 1.959724e-10, 
    1.939262e-10, 1.938714e-10, 1.936809e-10, 1.9383e-10, 1.935588e-10, 
    1.937102e-10, 1.937971e-10, 1.941347e-10, 1.942096e-10, 1.942783e-10, 
    1.944147e-10, 1.945897e-10, 1.949199e-10, 1.952187e-10, 1.954922e-10, 
    1.954722e-10, 1.954792e-10, 1.955401e-10, 1.95389e-10, 1.955649e-10, 
    1.955942e-10, 1.955172e-10, 1.959659e-10, 1.958376e-10, 1.959688e-10, 
    1.958854e-10, 1.938893e-10, 1.939815e-10, 1.939316e-10, 1.940253e-10, 
    1.939591e-10, 1.94253e-10, 1.943412e-10, 1.947626e-10, 1.945861e-10, 
    1.948752e-10, 1.946138e-10, 1.946567e-10, 1.94884e-10, 1.946271e-10, 
    1.952017e-10, 1.948056e-10, 1.955424e-10, 1.951452e-10, 1.955673e-10, 
    1.95491e-10, 1.956176e-10, 1.957307e-10, 1.958736e-10, 1.961367e-10, 
    1.960759e-10, 1.962965e-10, 1.941193e-10, 1.942389e-10, 1.942289e-10, 
    1.943545e-10, 1.944474e-10, 1.946495e-10, 1.950055e-10, 1.948697e-10, 
    1.951196e-10, 1.951696e-10, 1.947903e-10, 1.950226e-10, 1.943194e-10, 
    1.944269e-10, 1.943633e-10, 1.941285e-10, 1.949003e-10, 1.944932e-10, 
    1.952657e-10, 1.950322e-10, 1.957145e-10, 1.953744e-10, 1.960423e-10, 
    1.96327e-10, 1.965976e-10, 1.969114e-10, 1.943048e-10, 1.942234e-10, 
    1.943696e-10, 1.945712e-10, 1.947673e-10, 1.950464e-10, 1.950752e-10, 
    1.951274e-10, 1.952633e-10, 1.953773e-10, 1.951434e-10, 1.954059e-10, 
    1.944509e-10, 1.949379e-10, 1.941922e-10, 1.944082e-10, 1.945596e-10, 
    1.944937e-10, 1.948543e-10, 1.949447e-10, 1.953123e-10, 1.951225e-10, 
    1.962562e-10, 1.957539e-10, 1.971523e-10, 1.967604e-10, 1.941949e-10, 
    1.943048e-10, 1.946872e-10, 1.945051e-10, 1.950653e-10, 1.952086e-10, 
    1.953255e-10, 1.954743e-10, 1.954908e-10, 1.955791e-10, 1.954344e-10, 
    1.955735e-10, 1.95047e-10, 1.952822e-10, 1.94644e-10, 1.947943e-10, 
    1.947226e-10, 1.946489e-10, 1.948875e-10, 1.95147e-10, 1.951534e-10, 
    1.952365e-10, 1.954694e-10, 1.950677e-10, 1.963196e-10, 1.955443e-10, 
    1.944246e-10, 1.946356e-10, 1.946668e-10, 1.945848e-10, 1.951942e-10, 
    1.949684e-10, 1.95577e-10, 1.954126e-10, 1.956823e-10, 1.955482e-10, 
    1.955284e-10, 1.953564e-10, 1.952492e-10, 1.949786e-10, 1.94759e-10, 
    1.945968e-10, 1.94633e-10, 1.948166e-10, 1.951631e-10, 1.954919e-10, 
    1.954197e-10, 1.956618e-10, 1.95023e-10, 1.952902e-10, 1.951866e-10, 
    1.95457e-10, 1.948659e-10, 1.953667e-10, 1.947378e-10, 1.947931e-10, 
    1.94964e-10, 1.953078e-10, 1.953852e-10, 1.954663e-10, 1.954164e-10, 
    1.95172e-10, 1.951324e-10, 1.9496e-10, 1.94912e-10, 1.947811e-10, 
    1.946748e-10, 1.947715e-10, 1.948755e-10, 1.951724e-10, 1.954399e-10, 
    1.957322e-10, 1.958041e-10, 1.961441e-10, 1.958662e-10, 1.963238e-10, 
    1.95933e-10, 1.966107e-10, 1.953969e-10, 1.959231e-10, 1.94972e-10, 
    1.950745e-10, 1.952591e-10, 1.956848e-10, 1.954557e-10, 1.95724e-10, 
    1.951309e-10, 1.948227e-10, 1.947441e-10, 1.946061e-10, 1.947475e-10, 
    1.947352e-10, 1.948804e-10, 1.948338e-10, 1.951823e-10, 1.949951e-10, 
    1.955277e-10, 1.957221e-10, 1.962731e-10, 1.966109e-10, 1.969565e-10, 
    1.971088e-10, 1.971552e-10, 1.971746e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  2.450547, 2.427437, 2.431935, 2.413259, 2.423625, 2.411387, 2.445868, 
    2.426517, 2.438876, 2.448471, 2.376895, 2.412425, 2.339849, 2.362617, 
    2.305317, 2.343394, 2.297621, 2.306421, 2.279918, 2.287519, 2.253536, 
    2.276409, 2.235877, 2.259004, 2.255389, 2.277162, 2.405288, 2.381326, 
    2.406706, 2.403293, 2.404825, 2.42341, 2.432759, 2.452312, 2.448766, 
    2.434404, 2.401758, 2.412856, 2.384866, 2.385499, 2.354234, 2.368344, 
    2.315634, 2.330647, 2.287201, 2.298146, 2.287715, 2.29088, 2.287674, 
    2.303721, 2.296849, 2.310957, 2.365703, 2.349647, 2.397447, 2.426061, 
    2.44502, 2.458446, 2.456549, 2.452931, 2.43432, 2.416786, 2.4034, 
    2.394433, 2.38559, 2.358761, 2.344534, 2.312595, 2.318369, 2.308586, 
    2.299234, 2.283509, 2.286099, 2.279165, 2.308846, 2.289129, 2.321656, 
    2.312771, 2.383176, 2.409864, 2.421175, 2.431071, 2.45509, 2.438509, 
    2.445049, 2.429484, 2.419578, 2.424479, 2.394188, 2.405977, 2.343691, 
    2.370573, 2.300325, 2.317184, 2.29628, 2.306953, 2.288658, 2.305125, 
    2.276583, 2.270356, 2.274611, 2.258256, 2.306037, 2.287715, 2.424616, 
    2.423817, 2.420093, 2.436448, 2.437448, 2.452409, 2.439099, 2.433424, 
    2.419004, 2.410461, 2.402333, 2.384437, 2.364405, 2.336321, 2.316092, 
    2.302508, 2.310841, 2.303484, 2.311707, 2.315559, 2.272689, 2.296784, 
    2.26061, 2.262616, 2.278999, 2.26239, 2.423256, 2.427854, 2.443796, 
    2.431322, 2.454037, 2.441329, 2.434013, 2.405729, 2.399504, 2.393725, 
    2.382303, 2.367623, 2.34181, 2.319292, 2.29869, 2.300201, 2.299669, 
    2.29506, 2.306472, 2.293186, 2.290953, 2.296788, 2.262884, 2.272583, 
    2.262658, 2.268975, 2.42636, 2.41862, 2.422803, 2.414935, 2.420478, 
    2.395801, 2.388389, 2.353626, 2.367911, 2.345167, 2.365604, 2.361986, 
    2.344421, 2.364501, 2.320534, 2.350363, 2.294881, 2.324747, 2.293006, 
    2.298779, 2.28922, 2.280649, 2.269858, 2.249912, 2.254535, 2.237832, 
    2.40707, 2.397007, 2.397895, 2.387354, 2.37955, 2.362613, 2.33538, 
    2.345631, 2.326804, 2.32302, 2.351619, 2.334069, 2.390267, 2.38121, 
    2.386605, 2.406276, 2.343267, 2.375658, 2.315757, 2.333372, 2.281872, 
    2.307517, 2.257078, 2.235431, 2.215024, 2.191114, 2.391512, 2.398355, 
    2.3861, 2.369114, 2.353329, 2.332298, 2.330145, 2.326198, 2.315969, 
    2.30736, 2.324948, 2.3052, 2.379105, 2.340451, 2.400939, 2.382766, 
    2.370117, 2.375669, 2.346802, 2.339984, 2.312227, 2.326587, 2.240777, 
    2.278836, 2.172877, 2.202598, 2.400744, 2.391536, 2.359412, 2.374712, 
    2.330894, 2.320075, 2.311272, 2.300005, 2.298789, 2.292106, 2.303054, 
    2.292539, 2.332253, 2.314527, 2.363092, 2.351295, 2.356724, 2.362675, 
    2.344296, 2.324671, 2.324254, 2.317952, 2.300165, 2.330716, 2.235849, 
    2.294543, 2.381485, 2.363698, 2.361158, 2.368053, 2.32116, 2.338178, 
    2.292269, 2.304699, 2.284325, 2.294455, 2.295944, 2.308937, 2.317016, 
    2.337398, 2.353949, 2.367054, 2.364009, 2.349608, 2.32347, 2.298677, 
    2.304113, 2.285875, 2.334078, 2.313894, 2.321699, 2.301334, 2.345902, 
    2.307955, 2.355576, 2.351411, 2.338516, 2.312522, 2.306765, 2.300609, 
    2.304409, 2.322806, 2.325818, 2.33883, 2.342418, 2.352318, 2.360505, 
    2.353024, 2.345162, 2.322799, 2.302599, 2.280527, 2.275119, 2.249244, 
    2.270309, 2.235521, 2.265099, 2.213844, 2.305756, 2.265973, 2.33793, 
    2.330205, 2.316213, 2.28405, 2.30143, 2.281102, 2.325936, 2.349109, 
    2.355098, 2.366257, 2.354843, 2.355772, 2.344838, 2.348353, 2.322056, 
    2.336191, 2.29598, 2.281263, 2.239583, 2.213943, 2.187782, 2.17621, 
    2.172686, 2.171212,
  1.699967, 1.676936, 1.681416, 1.662822, 1.67314, 1.66096, 1.695302, 
    1.676019, 1.688332, 1.697897, 1.626684, 1.661992, 1.589966, 1.612523, 
    1.55583, 1.593475, 1.548234, 1.55692, 1.530781, 1.538271, 1.504813, 
    1.527324, 1.487466, 1.510192, 1.506636, 1.528065, 1.654895, 1.631081, 
    1.656304, 1.65291, 1.654434, 1.672926, 1.682235, 1.701729, 1.698192, 
    1.683875, 1.651384, 1.662422, 1.6346, 1.635229, 1.604214, 1.618203, 
    1.56602, 1.580862, 1.537959, 1.548753, 1.538465, 1.541586, 1.538425, 
    1.554254, 1.547473, 1.5614, 1.615583, 1.599669, 1.647099, 1.675563, 
    1.694456, 1.707848, 1.705955, 1.702346, 1.683791, 1.666333, 1.653017, 
    1.644104, 1.635319, 1.608698, 1.594605, 1.563017, 1.568723, 1.559058, 
    1.549827, 1.534319, 1.536872, 1.530038, 1.559315, 1.539859, 1.571972, 
    1.563191, 1.632918, 1.659445, 1.670699, 1.680555, 1.704499, 1.687966, 
    1.694485, 1.678975, 1.669111, 1.673991, 1.64386, 1.655579, 1.593769, 
    1.620413, 1.550904, 1.567552, 1.546912, 1.557446, 1.539394, 1.555641, 
    1.527495, 1.521362, 1.525553, 1.509457, 1.556542, 1.538464, 1.674127, 
    1.673331, 1.669624, 1.685912, 1.686909, 1.701825, 1.688554, 1.682899, 
    1.66854, 1.66004, 1.651956, 1.634174, 1.614295, 1.586475, 1.566473, 
    1.553058, 1.561285, 1.554021, 1.562141, 1.565946, 1.523659, 1.547409, 
    1.511772, 1.513745, 1.529875, 1.513523, 1.672772, 1.677351, 1.693237, 
    1.680806, 1.703449, 1.690777, 1.683485, 1.655331, 1.649144, 1.6434, 
    1.632056, 1.617487, 1.591908, 1.569635, 1.54929, 1.550781, 1.550256, 
    1.545709, 1.556971, 1.54386, 1.541657, 1.547413, 1.514009, 1.523555, 
    1.513787, 1.520003, 1.675863, 1.668158, 1.672322, 1.664491, 1.670007, 
    1.645462, 1.638098, 1.60361, 1.617773, 1.595232, 1.615485, 1.611897, 
    1.594491, 1.614392, 1.570861, 1.600376, 1.545532, 1.575025, 1.543683, 
    1.549378, 1.539949, 1.531501, 1.520873, 1.501252, 1.505797, 1.489387, 
    1.656667, 1.646661, 1.647545, 1.637071, 1.629321, 1.612519, 1.585544, 
    1.595692, 1.577062, 1.57332, 1.601623, 1.584246, 1.639964, 1.630968, 
    1.636327, 1.655876, 1.59335, 1.625458, 1.566142, 1.583558, 1.532705, 
    1.558002, 1.508298, 1.487028, 1.467015, 1.44361, 1.641201, 1.648002, 
    1.635826, 1.618965, 1.603317, 1.582495, 1.580365, 1.576462, 1.566352, 
    1.557847, 1.575225, 1.555716, 1.628877, 1.590562, 1.65057, 1.632513, 
    1.61996, 1.62547, 1.596852, 1.590101, 1.562653, 1.576847, 1.492276, 
    1.529713, 1.425796, 1.454845, 1.650377, 1.641226, 1.609345, 1.62452, 
    1.581106, 1.570408, 1.561711, 1.550587, 1.549387, 1.542794, 1.553597, 
    1.543222, 1.582451, 1.564926, 1.612994, 1.601301, 1.606682, 1.612581, 
    1.59437, 1.574951, 1.57454, 1.56831, 1.550741, 1.58093, 1.487435, 
    1.545194, 1.631243, 1.613593, 1.611076, 1.617914, 1.571481, 1.588314, 
    1.542956, 1.555221, 1.535123, 1.545111, 1.54658, 1.559405, 1.567386, 
    1.587541, 1.603931, 1.616923, 1.613903, 1.59963, 1.573764, 1.549277, 
    1.554642, 1.536651, 1.584256, 1.5643, 1.572013, 1.551899, 1.59596, 
    1.558432, 1.605544, 1.601417, 1.588648, 1.562944, 1.55726, 1.551183, 
    1.554934, 1.573108, 1.576086, 1.588959, 1.592511, 1.602316, 1.610429, 
    1.603015, 1.595227, 1.573102, 1.553147, 1.53138, 1.526053, 1.500594, 
    1.521314, 1.487113, 1.516184, 1.465856, 1.556261, 1.517046, 1.588068, 
    1.580425, 1.566591, 1.53485, 1.551994, 1.531946, 1.576203, 1.599136, 
    1.605071, 1.616133, 1.604818, 1.605738, 1.594907, 1.598388, 1.572367, 
    1.586347, 1.546616, 1.532105, 1.491105, 1.465955, 1.440355, 1.42905, 
    1.42561, 1.424171,
  0.7771534, 0.7632287, 0.7659328, 0.7547256, 0.7609397, 0.7536058, 
    0.7743278, 0.7626759, 0.7701113, 0.7758994, 0.7330593, 0.7542265, 
    0.7112027, 0.7246109, 0.6910276, 0.7132847, 0.6865579, 0.6916698, 
    0.6763138, 0.6807056, 0.6611418, 0.6742889, 0.651054, 0.6642774, 
    0.6622041, 0.6747233, 0.7499599, 0.7356879, 0.7508066, 0.748768, 
    0.7496831, 0.7608105, 0.7664275, 0.778221, 0.776078, 0.767418, 0.7478517, 
    0.7544849, 0.7377924, 0.7381686, 0.7196646, 0.7279965, 0.6970356, 
    0.7058083, 0.6805222, 0.6868628, 0.6808194, 0.682651, 0.6807956, 0.6901, 
    0.6861101, 0.6943101, 0.7264342, 0.7169626, 0.7452802, 0.762401, 
    0.7738158, 0.7819316, 0.7807834, 0.7785949, 0.7673673, 0.7568388, 
    0.748832, 0.7434845, 0.7382227, 0.7223333, 0.713955, 0.6952634, 0.698631, 
    0.6929295, 0.6874944, 0.6783873, 0.6798848, 0.6758784, 0.6930811, 
    0.6816372, 0.7005503, 0.6953664, 0.7367862, 0.7526947, 0.7594689, 
    0.7654126, 0.7799006, 0.7698901, 0.7738336, 0.7644591, 0.7585118, 
    0.7614526, 0.7433383, 0.750371, 0.7134591, 0.729315, 0.6881279, 
    0.6979397, 0.6857807, 0.6919799, 0.6813646, 0.6909168, 0.6743892, 
    0.670801, 0.6732525, 0.6638488, 0.6914469, 0.6808187, 0.7615346, 
    0.7610548, 0.7588211, 0.7686486, 0.7692509, 0.7782794, 0.7702456, 
    0.7668282, 0.7581679, 0.7530521, 0.7481954, 0.7375372, 0.7256667, 
    0.7091327, 0.6973027, 0.6893955, 0.6942424, 0.6899628, 0.6947469, 
    0.6969919, 0.6721445, 0.6860725, 0.6651995, 0.666351, 0.6757829, 
    0.6662213, 0.760718, 0.7634794, 0.7730778, 0.7655644, 0.7792637, 
    0.7715895, 0.7671822, 0.7502224, 0.746507, 0.7430626, 0.7362702, 
    0.7275696, 0.7123545, 0.6991696, 0.6871788, 0.688056, 0.6877471, 
    0.6850731, 0.6916996, 0.6839867, 0.6826933, 0.686075, 0.6665053, 
    0.6720837, 0.6663755, 0.6700065, 0.7625818, 0.7579378, 0.7604465, 
    0.7557298, 0.7590516, 0.7442989, 0.739886, 0.7193056, 0.7277402, 
    0.7143274, 0.7263761, 0.7242379, 0.7138877, 0.7257245, 0.6998939, 
    0.7173833, 0.6849693, 0.7023552, 0.6838827, 0.6872305, 0.6816902, 
    0.6767356, 0.6705148, 0.6590679, 0.661715, 0.6521686, 0.7510245, 
    0.7450178, 0.7455477, 0.7392712, 0.7346355, 0.7246085, 0.7085811, 
    0.7146003, 0.7035595, 0.7013468, 0.7181242, 0.7078124, 0.7410038, 
    0.7356201, 0.7388256, 0.7505496, 0.7132105, 0.732327, 0.6971073, 
    0.7074045, 0.6774414, 0.6923073, 0.6631728, 0.6507995, 0.6392093, 
    0.6257198, 0.7417448, 0.7458218, 0.7385259, 0.7284513, 0.7191312, 
    0.7067752, 0.7055143, 0.7032047, 0.6972312, 0.6922162, 0.7024735, 
    0.6909604, 0.7343699, 0.7115564, 0.747363, 0.736544, 0.729045, 0.7323342, 
    0.7152892, 0.7112828, 0.6950492, 0.7034323, 0.6538472, 0.6756881, 
    0.6154998, 0.6321864, 0.7472469, 0.7417594, 0.7227184, 0.7317666, 
    0.7059527, 0.6996265, 0.6944935, 0.6879414, 0.6872358, 0.6833609, 
    0.6897129, 0.683612, 0.706749, 0.69639, 0.7248917, 0.7179329, 0.7211331, 
    0.7246455, 0.7138156, 0.7023114, 0.7020682, 0.6983872, 0.6880323, 
    0.7058485, 0.6510361, 0.6847709, 0.7357841, 0.7252487, 0.7237489, 
    0.7278245, 0.7002601, 0.7102229, 0.6834556, 0.6906692, 0.6788588, 
    0.684722, 0.6855854, 0.693134, 0.6978418, 0.7097651, 0.7194968, 
    0.7272334, 0.7254332, 0.7169397, 0.7016094, 0.6871709, 0.6903281, 
    0.6797549, 0.7078182, 0.6960208, 0.700575, 0.6887136, 0.7147598, 
    0.6925607, 0.7204558, 0.7180017, 0.710421, 0.6952206, 0.6918702, 
    0.6882925, 0.6905001, 0.7012215, 0.7029822, 0.7106056, 0.7127122, 
    0.718536, 0.7233636, 0.7189521, 0.7143244, 0.7012179, 0.6894481, 
    0.6766648, 0.6735451, 0.658685, 0.6707732, 0.6508488, 0.6677752, 0.63854, 
    0.691282, 0.6682789, 0.7100772, 0.7055495, 0.6973727, 0.678699, 
    0.6887693, 0.6769963, 0.7030514, 0.716646, 0.7201744, 0.7267622, 
    0.720024, 0.7205716, 0.7141343, 0.7162019, 0.7007836, 0.7090573, 
    0.6856065, 0.6770896, 0.6531668, 0.6385971, 0.6238493, 0.6173637, 
    0.6153932, 0.6145698,
  0.1899293, 0.1849349, 0.1859014, 0.1819064, 0.184118, 0.1815088, 0.1889123, 
    0.1847376, 0.1873981, 0.1894777, 0.1742636, 0.1817292, 0.1666619, 
    0.1713121, 0.1597438, 0.1673813, 0.158224, 0.1599624, 0.1547587, 
    0.1562412, 0.1496727, 0.1540767, 0.1463216, 0.1507193, 0.150027, 
    0.1542229, 0.1802161, 0.1751851, 0.180516, 0.1797942, 0.1801181, 
    0.184072, 0.1860785, 0.1903139, 0.189542, 0.186433, 0.1794701, 0.1818209, 
    0.1759239, 0.1760561, 0.1695918, 0.1724928, 0.1617939, 0.1648028, 
    0.1561792, 0.1583275, 0.1562797, 0.1568994, 0.1562717, 0.1594279, 
    0.158072, 0.1608628, 0.1719476, 0.1686544, 0.1785614, 0.1846395, 
    0.1887283, 0.191653, 0.1912383, 0.1904488, 0.1864148, 0.1826575, 
    0.1798168, 0.1779277, 0.1760751, 0.1705194, 0.1676131, 0.1611883, 
    0.1623397, 0.1603918, 0.158542, 0.1554581, 0.1559638, 0.154612, 
    0.1604435, 0.1565564, 0.1629972, 0.1612234, 0.1755707, 0.1811855, 
    0.1835939, 0.1857154, 0.1909197, 0.1873188, 0.1887347, 0.1853745, 
    0.1832529, 0.1843009, 0.1778761, 0.1803617, 0.1674416, 0.1729534, 
    0.1587572, 0.1621031, 0.1579602, 0.1600681, 0.1564641, 0.1597059, 
    0.1541105, 0.1529043, 0.153728, 0.150576, 0.1598865, 0.1562795, 
    0.1843302, 0.1841591, 0.183363, 0.1868738, 0.1870896, 0.190335, 
    0.1874463, 0.1862218, 0.1831304, 0.1813123, 0.1795916, 0.1758342, 
    0.17168, 0.1659478, 0.1618852, 0.1591882, 0.1608396, 0.1593812, 
    0.1610119, 0.1617789, 0.1533556, 0.1580592, 0.1510274, 0.1514126, 
    0.1545798, 0.1513692, 0.184039, 0.1850244, 0.188463, 0.1857696, 
    0.1906899, 0.1879285, 0.1863486, 0.1803091, 0.1789947, 0.1777789, 
    0.1753893, 0.1723438, 0.1670597, 0.1625242, 0.1584347, 0.1587328, 
    0.1586278, 0.1577202, 0.1599726, 0.1573518, 0.1569138, 0.15806, 
    0.1514643, 0.1533351, 0.1514208, 0.1526376, 0.1847039, 0.1830485, 
    0.1839422, 0.1822632, 0.1834452, 0.178215, 0.1766602, 0.1694672, 
    0.1724034, 0.1677419, 0.1719274, 0.1711822, 0.1675899, 0.1717001, 
    0.1627723, 0.1688003, 0.1576849, 0.1636164, 0.1573166, 0.1584523, 
    0.1565742, 0.1549009, 0.1528082, 0.1489817, 0.1498638, 0.1466907, 
    0.1805933, 0.1784687, 0.1786558, 0.1764438, 0.1748158, 0.1713112, 
    0.1657576, 0.1678363, 0.1640298, 0.1632703, 0.1690571, 0.1654927, 
    0.1770535, 0.1751612, 0.1762871, 0.180425, 0.1673556, 0.174007, 
    0.1618184, 0.1653522, 0.1551389, 0.1601797, 0.1503503, 0.1462375, 
    0.1424187, 0.1380159, 0.1773145, 0.1787526, 0.1761817, 0.1726516, 
    0.1694066, 0.1651355, 0.1647016, 0.1639079, 0.1618608, 0.1601486, 
    0.1636569, 0.1597208, 0.1747228, 0.1667841, 0.1792972, 0.1754855, 
    0.172859, 0.1740094, 0.1680747, 0.1666895, 0.1611151, 0.1639861, 
    0.1472471, 0.1545479, 0.1347103, 0.1401209, 0.1792562, 0.1773196, 
    0.1706533, 0.1738107, 0.1648524, 0.1626807, 0.1609254, 0.1586939, 
    0.1584541, 0.1571398, 0.1592962, 0.1572249, 0.1651265, 0.1615732, 
    0.1714099, 0.1689909, 0.1701019, 0.1713241, 0.1675648, 0.1636013, 
    0.1635178, 0.1622563, 0.158725, 0.1648166, 0.1463159, 0.1576179, 
    0.1752187, 0.1715344, 0.1710119, 0.1724327, 0.1628978, 0.1663237, 
    0.1571719, 0.1596216, 0.1556173, 0.1576011, 0.1578939, 0.1604615, 
    0.1620696, 0.1661658, 0.1695335, 0.1722264, 0.1715986, 0.1686465, 
    0.1633604, 0.1584321, 0.1595056, 0.1559199, 0.1654947, 0.161447, 
    0.1630057, 0.1589563, 0.1678915, 0.1602663, 0.1698665, 0.1690147, 
    0.1663921, 0.1611737, 0.1600307, 0.1588132, 0.1595641, 0.1632274, 
    0.1638315, 0.1664557, 0.1671833, 0.1692, 0.1708777, 0.1693444, 0.1677408, 
    0.1632261, 0.1592061, 0.154877, 0.1538264, 0.1488543, 0.152895, 0.146254, 
    0.1518898, 0.1421993, 0.1598304, 0.1520584, 0.1662734, 0.1647137, 
    0.1619092, 0.1555634, 0.1589752, 0.1549888, 0.1638553, 0.1685448, 
    0.1697688, 0.172062, 0.1697166, 0.1699068, 0.1676751, 0.1683908, 
    0.1630772, 0.1659217, 0.1579011, 0.1550203, 0.1470215, 0.142218, 
    0.1374089, 0.1353112, 0.1346759, 0.1344107,
  0.01658138, 0.01594443, 0.01606706, 0.01556211, 0.01584101, 0.01551213, 
    0.01645103, 0.01591943, 0.01625756, 0.01652345, 0.01461064, 0.01553983, 
    0.01368358, 0.01424837, 0.01285697, 0.01377047, 0.0126776, 0.01288283, 
    0.01227163, 0.01244479, 0.01168352, 0.01219223, 0.01130109, 0.01180378, 
    0.01172418, 0.01220924, 0.01535002, 0.01472434, 0.01538759, 0.01529723, 
    0.01533775, 0.01583518, 0.01608957, 0.01663076, 0.01653169, 0.01613463, 
    0.01525672, 0.01555135, 0.01481568, 0.01483205, 0.01403857, 0.01439293, 
    0.0131002, 0.01345981, 0.01243754, 0.01268978, 0.0124493, 0.01252192, 
    0.01244836, 0.01281962, 0.01265969, 0.01298955, 0.01432613, 0.01392468, 
    0.0151433, 0.01590702, 0.01642747, 0.01680305, 0.01674964, 0.01664808, 
    0.01613233, 0.01565664, 0.01530006, 0.01506437, 0.0148344, 0.01415158, 
    0.01379851, 0.0130282, 0.0131652, 0.0129337, 0.01271505, 0.01235323, 
    0.01241233, 0.01225454, 0.01293981, 0.0124817, 0.01324364, 0.01303237, 
    0.014772, 0.01547153, 0.01577477, 0.01604343, 0.01670863, 0.01624745, 
    0.01642829, 0.01600016, 0.01573172, 0.01586414, 0.01505796, 0.01536825, 
    0.01377776, 0.01444945, 0.01274043, 0.01313701, 0.01264654, 0.01289534, 
    0.0124709, 0.01285249, 0.01219616, 0.01205613, 0.01215171, 0.01178729, 
    0.01287385, 0.01244928, 0.01586785, 0.0158462, 0.01574561, 0.01619074, 
    0.01621824, 0.01663346, 0.0162637, 0.01610778, 0.01571626, 0.01548745, 
    0.01527189, 0.01480459, 0.01429337, 0.01359748, 0.01311107, 0.0127913, 
    0.0129868, 0.0128141, 0.01300724, 0.01309841, 0.01210847, 0.01265819, 
    0.01183927, 0.01188367, 0.0122508, 0.01187866, 0.01583101, 0.01595576, 
    0.01639354, 0.01605032, 0.01667908, 0.01632525, 0.0161239, 0.01536167, 
    0.01519734, 0.01504587, 0.01474956, 0.01437466, 0.0137316, 0.0131872, 
    0.01270242, 0.01273755, 0.01272517, 0.01261831, 0.01288404, 0.01257502, 
    0.0125236, 0.01265829, 0.01188963, 0.01210608, 0.01188462, 0.01202524, 
    0.01591515, 0.01570594, 0.01581877, 0.01560699, 0.01575598, 0.01510016, 
    0.01490691, 0.01402342, 0.01438196, 0.01381409, 0.01432364, 0.01423249, 
    0.0137957, 0.01429582, 0.0132168, 0.01394239, 0.01261416, 0.01331766, 
    0.01257088, 0.01270449, 0.01248379, 0.01228821, 0.012045, 0.01160433, 
    0.01170544, 0.01134301, 0.01539726, 0.01513176, 0.01515507, 0.01488008, 
    0.01467872, 0.01424826, 0.01357458, 0.01382551, 0.01336712, 0.01327627, 
    0.01397357, 0.01354271, 0.01495572, 0.01472138, 0.01486066, 0.01537618, 
    0.01376736, 0.01457902, 0.01310312, 0.01352581, 0.01231597, 0.01290857, 
    0.01176133, 0.01129155, 0.01086084, 0.01037097, 0.01498813, 0.01516714, 
    0.0148476, 0.01441242, 0.01401605, 0.01349978, 0.01344767, 0.01335253, 
    0.01310816, 0.01290488, 0.0133225, 0.01285424, 0.01466727, 0.01369831, 
    0.01523512, 0.01476146, 0.01443787, 0.01457931, 0.01385438, 0.0136869, 
    0.01301951, 0.01336189, 0.01140631, 0.01224708, 0.01000793, 0.01060428, 
    0.01522999, 0.01498877, 0.0141679, 0.01455485, 0.01346577, 0.01320586, 
    0.01299697, 0.01273296, 0.0127047, 0.01255013, 0.01280405, 0.01256011, 
    0.01349869, 0.01307394, 0.01426032, 0.01396552, 0.01410067, 0.01424983, 
    0.01379266, 0.01331585, 0.01330585, 0.01315527, 0.01273665, 0.01346147, 
    0.01130046, 0.0126063, 0.01472847, 0.01427555, 0.01421168, 0.01438556, 
    0.01323177, 0.01364277, 0.01255389, 0.01284252, 0.01237182, 0.01260431, 
    0.01263874, 0.01294195, 0.01313302, 0.01362374, 0.01403148, 0.01436027, 
    0.0142834, 0.01392372, 0.01328704, 0.01270211, 0.0128288, 0.0124072, 
    0.01354294, 0.01305894, 0.01324466, 0.01276392, 0.0138322, 0.01291883, 
    0.01407201, 0.01396841, 0.01365101, 0.01302647, 0.01289091, 0.01274704, 
    0.01283571, 0.01327114, 0.01334339, 0.01365869, 0.01374653, 0.01399093, 
    0.0141953, 0.01400848, 0.01381396, 0.01327098, 0.01279342, 0.01228543, 
    0.01216314, 0.01158976, 0.01205507, 0.01129343, 0.01193877, 0.01083628, 
    0.01286723, 0.01195825, 0.01363671, 0.01344912, 0.01311393, 0.01236553, 
    0.01276616, 0.01229847, 0.01334623, 0.01391137, 0.01406011, 0.01434013, 
    0.01405375, 0.01407691, 0.01380599, 0.01389269, 0.01325319, 0.01359433, 
    0.01263959, 0.01230214, 0.01138062, 0.01083835, 0.01030398, 0.01007361, 
    0.01000417, 0.009975231,
  0.0004568995, 0.0004322279, 0.0004369482, 0.0004176034, 0.0004282579, 
    0.0004157022, 0.0004518195, 0.0004312674, 0.0004443091, 0.00045464, 
    0.0003818243, 0.0004167554, 0.0003478366, 0.0003684378, 0.0003182909, 
    0.0003509849, 0.000311977, 0.0003192042, 0.0002978184, 0.0003038352, 
    0.0002776381, 0.000295071, 0.0002647305, 0.0002817323, 0.0002790206, 
    0.0002956589, 0.0004095511, 0.0003860531, 0.0004109741, 0.0004075538, 
    0.0004090866, 0.0004280349, 0.0004378163, 0.0004588276, 0.0004549612, 
    0.0004395555, 0.0004060225, 0.0004171938, 0.0003894587, 0.00039007, 
    0.0003607468, 0.0003737635, 0.0003269086, 0.0003397664, 0.0003035824, 
    0.0003124046, 0.0003039923, 0.0003065258, 0.0003039594, 0.0003169731, 
    0.0003113487, 0.0003229801, 0.0003712998, 0.0003565906, 0.0004017449, 
    0.0004307909, 0.0004509032, 0.000465574, 0.0004634795, 0.0004595049, 
    0.0004394664, 0.0004212065, 0.0004076604, 0.0003987752, 0.0003901579, 
    0.0003648842, 0.0003520021, 0.000324351, 0.0003292225, 0.0003210024, 
    0.0003132925, 0.0003006495, 0.0003027047, 0.0002972265, 0.0003212188, 
    0.0003051221, 0.0003320205, 0.0003244988, 0.0003878294, 0.000414159, 
    0.0004257213, 0.0004360376, 0.0004618736, 0.0004439178, 0.0004509352, 
    0.0004343712, 0.0004240739, 0.0004291451, 0.0003985342, 0.0004102416, 
    0.0003512491, 0.0003758517, 0.0003141847, 0.0003282185, 0.0003108871, 
    0.000319646, 0.0003047451, 0.0003181325, 0.0002952068, 0.0002903781, 
    0.0002936714, 0.0002811698, 0.0003188867, 0.0003039916, 0.0004292873, 
    0.000428457, 0.0004246052, 0.0004417235, 0.000442787, 0.0004589335, 
    0.000444547, 0.0004385189, 0.0004234832, 0.0004147638, 0.0004065959, 
    0.0003890446, 0.0003700936, 0.0003447252, 0.0003272952, 0.000315975, 
    0.0003228826, 0.0003167785, 0.0003236074, 0.0003268451, 0.00029218, 
    0.0003112961, 0.0002829436, 0.0002844615, 0.0002970968, 0.0002842901, 
    0.0004278749, 0.0004326636, 0.0004495844, 0.0004363029, 0.000460717, 
    0.0004469328, 0.0004391412, 0.0004099923, 0.0004037814, 0.0003980799, 
    0.0003869921, 0.0003730892, 0.0003495754, 0.0003300064, 0.0003128485, 
    0.0003140832, 0.0003136481, 0.0003098977, 0.0003192466, 0.0003083822, 
    0.0003065847, 0.0003112994, 0.0002846651, 0.0002920979, 0.0002844938, 
    0.0002893155, 0.000431103, 0.0004230886, 0.0004274058, 0.000419313, 
    0.0004250021, 0.0004001209, 0.0003928696, 0.0003601932, 0.0003733588, 
    0.0003525678, 0.0003712082, 0.0003678541, 0.0003519004, 0.0003701837, 
    0.0003310626, 0.0003572364, 0.0003097526, 0.0003346676, 0.0003082374, 
    0.0003129212, 0.0003051949, 0.000298393, 0.0002899948, 0.000274951, 
    0.000278383, 0.0002661366, 0.0004113408, 0.0004013102, 0.0004021879, 
    0.0003918653, 0.0003843544, 0.0003684337, 0.000343899, 0.0003529824, 
    0.0003364392, 0.0003331865, 0.000358373, 0.0003427502, 0.0003946974, 
    0.0003859424, 0.0003911394, 0.000410542, 0.0003508718, 0.0003806503, 
    0.0003270123, 0.0003421413, 0.0002993558, 0.0003201136, 0.0002802853, 
    0.0002644106, 0.0002500868, 0.0002340716, 0.0003959125, 0.0004026429, 
    0.0003906511, 0.0003744834, 0.0003599238, 0.0003412039, 0.0003393301, 
    0.0003359164, 0.0003271915, 0.0003199832, 0.0003348406, 0.0003181946, 
    0.0003839286, 0.0003483698, 0.000405207, 0.0003874358, 0.0003754236, 
    0.0003806612, 0.0003540319, 0.0003479566, 0.0003240425, 0.0003362516, 
    0.0002682647, 0.0002969685, 0.000222397, 0.0002416622, 0.0004050132, 
    0.0003959364, 0.0003654828, 0.0003797539, 0.0003399808, 0.000330672, 
    0.0003232434, 0.0003139221, 0.0003129287, 0.0003075116, 0.0003164243, 
    0.0003078608, 0.0003411649, 0.0003259752, 0.0003688772, 0.0003580794, 
    0.0003630186, 0.0003684915, 0.0003517894, 0.0003346025, 0.0003342446, 
    0.0003288685, 0.0003140523, 0.0003398261, 0.0002647096, 0.0003094776, 
    0.0003862062, 0.0003694378, 0.0003670896, 0.0003734916, 0.0003315968, 
    0.0003463611, 0.0003076432, 0.0003177807, 0.0003012955, 0.0003094073, 
    0.0003106139, 0.0003212944, 0.0003280765, 0.0003456734, 0.0003604878, 
    0.0003725585, 0.0003697263, 0.0003565556, 0.000333572, 0.0003128377, 
    0.0003172969, 0.000302526, 0.0003427584, 0.0003254424, 0.0003320572, 
    0.0003150111, 0.0003532256, 0.0003204769, 0.0003619694, 0.0003581848, 
    0.0003466589, 0.0003242897, 0.0003194896, 0.000314417, 0.0003175406, 
    0.0003330033, 0.0003355888, 0.0003469365, 0.0003501165, 0.0003590066, 
    0.0003664879, 0.0003596474, 0.000352563, 0.0003329977, 0.0003160498, 
    0.0002982966, 0.000294066, 0.0002744578, 0.0002903416, 0.000264474, 
    0.0002863487, 0.0002492771, 0.0003186531, 0.000287016, 0.0003461418, 
    0.0003393823, 0.0003273971, 0.0003010771, 0.0003150898, 0.0002987489, 
    0.0003356906, 0.000356106, 0.0003615343, 0.0003718159, 0.0003613017, 
    0.0003621488, 0.0003522736, 0.0003554257, 0.000332362, 0.0003446116, 
    0.0003106436, 0.0002988761, 0.0002674005, 0.0002493454, 0.0002319048, 
    0.0002244967, 0.0002222771, 0.0002213539,
  3.512436e-06, 3.239124e-06, 3.290964e-06, 3.07991e-06, 3.195695e-06, 
    3.059367e-06, 3.455686e-06, 3.228604e-06, 3.372232e-06, 3.487164e-06, 
    2.699576e-06, 3.070742e-06, 2.351069e-06, 2.560771e-06, 2.058988e-06, 
    2.382802e-06, 1.997956e-06, 2.067856e-06, 1.862941e-06, 1.92e-06, 
    1.675088e-06, 1.837044e-06, 1.557881e-06, 1.712752e-06, 1.68778e-06, 
    1.842578e-06, 2.993157e-06, 2.743828e-06, 3.00844e-06, 2.971742e-06, 
    2.988173e-06, 3.19326e-06, 3.300523e-06, 3.534039e-06, 3.490754e-06, 
    3.319691e-06, 2.955351e-06, 3.07548e-06, 2.779601e-06, 2.786036e-06, 
    2.48192e-06, 2.615757e-06, 2.14309e-06, 2.270251e-06, 1.917592e-06, 
    2.002072e-06, 1.921496e-06, 1.945667e-06, 1.921182e-06, 2.046208e-06, 
    1.991909e-06, 2.104636e-06, 2.590281e-06, 2.439587e-06, 2.909689e-06, 
    3.223389e-06, 3.445476e-06, 3.609898e-06, 3.586302e-06, 3.541636e-06, 
    3.318708e-06, 3.118937e-06, 2.972883e-06, 2.8781e-06, 2.786962e-06, 
    2.524258e-06, 2.39308e-06, 2.118035e-06, 2.165826e-06, 2.085351e-06, 
    2.010629e-06, 1.88973e-06, 1.909243e-06, 1.857354e-06, 2.087458e-06, 
    1.932265e-06, 2.193406e-06, 2.11948e-06, 2.762473e-06, 3.04272e-06, 
    3.168027e-06, 3.280947e-06, 3.568236e-06, 3.367899e-06, 3.445832e-06, 
    3.262635e-06, 3.150091e-06, 3.205386e-06, 2.875541e-06, 3.00057e-06, 
    2.38547e-06, 2.637402e-06, 2.019238e-06, 2.155953e-06, 1.98747e-06, 
    2.072151e-06, 1.92867e-06, 2.05745e-06, 1.838323e-06, 1.793042e-06, 
    1.823891e-06, 1.707563e-06, 2.064772e-06, 1.921489e-06, 3.206941e-06, 
    3.197869e-06, 3.155872e-06, 3.343627e-06, 3.355385e-06, 3.535226e-06, 
    3.374868e-06, 3.308262e-06, 3.143666e-06, 3.049241e-06, 2.961485e-06, 
    2.775245e-06, 2.577833e-06, 2.319819e-06, 2.146883e-06, 2.036542e-06, 
    2.103684e-06, 2.044321e-06, 2.110764e-06, 2.142465e-06, 1.809904e-06, 
    1.991403e-06, 1.723938e-06, 1.737986e-06, 1.85613e-06, 1.736399e-06, 
    3.191512e-06, 3.2439e-06, 3.430794e-06, 3.283864e-06, 3.555241e-06, 
    3.401326e-06, 3.315122e-06, 2.997894e-06, 2.931404e-06, 2.870718e-06, 
    2.753676e-06, 2.608777e-06, 2.36858e-06, 2.173545e-06, 2.006348e-06, 
    2.018258e-06, 2.014059e-06, 1.977965e-06, 2.068269e-06, 1.963431e-06, 
    1.946231e-06, 1.991434e-06, 1.739874e-06, 1.809133e-06, 1.738286e-06, 
    1.783119e-06, 3.226803e-06, 3.139377e-06, 3.186392e-06, 3.098411e-06, 
    3.160193e-06, 2.892404e-06, 2.815559e-06, 2.476272e-06, 2.611567e-06, 
    2.3988e-06, 2.589335e-06, 2.554763e-06, 2.392052e-06, 2.578761e-06, 
    2.183956e-06, 2.446153e-06, 1.976573e-06, 2.219589e-06, 1.962044e-06, 
    2.007049e-06, 1.932959e-06, 1.86837e-06, 1.789461e-06, 1.650494e-06, 
    1.681922e-06, 1.570534e-06, 3.012381e-06, 2.905059e-06, 2.914408e-06, 
    2.804958e-06, 2.726025e-06, 2.560728e-06, 2.31154e-06, 2.402994e-06, 
    2.237155e-06, 2.204928e-06, 2.457717e-06, 2.300042e-06, 2.834876e-06, 
    2.742665e-06, 2.797303e-06, 3.003797e-06, 2.38166e-06, 2.687323e-06, 
    2.144107e-06, 2.293954e-06, 1.877476e-06, 2.0767e-06, 1.699413e-06, 
    1.555007e-06, 1.427829e-06, 1.289315e-06, 2.847737e-06, 2.919258e-06, 
    2.792156e-06, 2.623214e-06, 2.473522e-06, 2.284591e-06, 2.265904e-06, 
    2.231966e-06, 2.145865e-06, 2.075429e-06, 2.221302e-06, 2.058052e-06, 
    2.721572e-06, 2.356435e-06, 2.946631e-06, 2.758337e-06, 2.632961e-06, 
    2.687435e-06, 2.413622e-06, 2.352275e-06, 2.115017e-06, 2.235293e-06, 
    1.589739e-06, 1.85492e-06, 1.190905e-06, 1.35447e-06, 2.944559e-06, 
    2.84799e-06, 2.530397e-06, 2.677978e-06, 2.272388e-06, 2.180103e-06, 
    2.107207e-06, 2.016703e-06, 2.007122e-06, 1.955095e-06, 2.040892e-06, 
    1.958437e-06, 2.284201e-06, 2.133935e-06, 2.565295e-06, 2.454728e-06, 
    2.505142e-06, 2.561323e-06, 2.390928e-06, 2.218943e-06, 2.215398e-06, 
    2.162344e-06, 2.017964e-06, 2.270846e-06, 1.557697e-06, 1.973937e-06, 
    2.74543e-06, 2.571072e-06, 2.546901e-06, 2.612941e-06, 2.189224e-06, 
    2.336234e-06, 1.956354e-06, 2.054036e-06, 1.895857e-06, 1.973259e-06, 
    1.984844e-06, 2.088195e-06, 2.154557e-06, 2.32933e-06, 2.479276e-06, 
    2.603287e-06, 2.574045e-06, 2.439231e-06, 2.208742e-06, 2.006245e-06, 
    2.049346e-06, 1.907544e-06, 2.300124e-06, 2.128716e-06, 2.19377e-06, 
    2.027221e-06, 2.405456e-06, 2.080238e-06, 2.49441e-06, 2.455801e-06, 
    2.339226e-06, 2.117435e-06, 2.07063e-06, 2.021482e-06, 2.051708e-06, 
    2.203118e-06, 2.228718e-06, 2.342015e-06, 2.374037e-06, 2.464171e-06, 
    2.540716e-06, 2.470703e-06, 2.398751e-06, 2.203062e-06, 2.037267e-06, 
    1.867459e-06, 1.827596e-06, 1.645992e-06, 1.792702e-06, 1.555579e-06, 
    1.7555e-06, 1.420733e-06, 2.062505e-06, 1.761701e-06, 2.334031e-06, 
    2.266423e-06, 2.147885e-06, 1.893786e-06, 2.027981e-06, 1.871735e-06, 
    2.229727e-06, 2.434664e-06, 2.489963e-06, 2.595612e-06, 2.487587e-06, 
    2.496244e-06, 2.395824e-06, 2.427756e-06, 2.19678e-06, 2.31868e-06, 
    1.98513e-06, 1.872938e-06, 1.581931e-06, 1.42133e-06, 1.270882e-06, 
    1.208439e-06, 1.189905e-06, 1.18222e-06,
  4.243282e-09, 3.591658e-09, 3.712521e-09, 3.228801e-09, 3.491416e-09, 
    3.182924e-09, 4.105103e-09, 3.567291e-09, 3.904607e-09, 4.181563e-09, 
    2.416473e-09, 3.208299e-09, 1.747137e-09, 2.140708e-09, 1.249524e-09, 
    1.804838e-09, 1.153636e-09, 1.2637e-09, 9.522626e-10, 1.035516e-09, 
    6.984192e-10, 9.153948e-10, 5.568496e-10, 7.467294e-10, 7.145485e-10, 
    9.232246e-10, 3.036561e-09, 2.506811e-09, 3.070141e-09, 2.98972e-09, 
    3.025638e-09, 3.485825e-09, 3.734955e-09, 4.296262e-09, 4.190313e-09, 
    3.78006e-09, 2.954033e-09, 3.218886e-09, 2.580662e-09, 2.594027e-09, 
    1.989371e-09, 2.248543e-09, 1.386387e-09, 1.603302e-09, 1.031948e-09, 
    1.16001e-09, 1.037735e-09, 1.073857e-09, 1.03727e-09, 1.229201e-09, 
    1.144296e-09, 1.32314e-09, 2.19835e-09, 1.909767e-09, 2.855384e-09, 
    3.555235e-09, 4.0804e-09, 4.483974e-09, 4.425312e-09, 4.314946e-09, 
    3.777744e-09, 3.316557e-09, 2.992207e-09, 2.787805e-09, 2.595952e-09, 
    2.070145e-09, 1.82367e-09, 1.345052e-09, 1.424304e-09, 1.291844e-09, 
    1.173303e-09, 9.910067e-10, 1.019611e-09, 9.442599e-10, 1.295249e-09, 
    1.05377e-09, 1.470812e-09, 1.347422e-09, 2.545216e-09, 3.145905e-09, 
    3.428051e-09, 3.689066e-09, 4.380567e-09, 3.894288e-09, 4.081261e-09, 
    3.646308e-09, 3.387169e-09, 3.513702e-09, 2.782354e-09, 3.052833e-09, 
    1.809718e-09, 2.291503e-09, 1.186737e-09, 1.407792e-09, 1.137459e-09, 
    1.270586e-09, 1.048406e-09, 1.247069e-09, 9.172019e-10, 8.540977e-10, 
    8.968942e-10, 7.39993e-10, 1.258761e-09, 1.037726e-09, 3.517282e-09, 
    3.496412e-09, 3.400326e-09, 3.836637e-09, 3.864529e-09, 4.29918e-09, 
    3.910889e-09, 3.753143e-09, 3.372565e-09, 3.160389e-09, 2.96737e-09, 
    2.57163e-09, 2.17397e-09, 1.690984e-09, 1.392687e-09, 1.213916e-09, 
    1.321588e-09, 1.226212e-09, 1.333144e-09, 1.385351e-09, 8.773857e-10, 
    1.143517e-09, 7.613334e-10, 7.798379e-10, 9.425113e-10, 7.777382e-10, 
    3.481811e-09, 3.602734e-09, 4.044962e-09, 3.695888e-09, 4.348468e-09, 
    3.974135e-09, 3.769294e-09, 3.046959e-09, 2.902153e-09, 2.772093e-09, 
    2.527061e-09, 2.234751e-09, 1.778891e-09, 1.437265e-09, 1.166645e-09, 
    1.185205e-09, 1.178647e-09, 1.122873e-09, 1.26436e-09, 1.10071e-09, 
    1.074706e-09, 1.143564e-09, 7.823382e-10, 8.763154e-10, 7.802344e-10, 
    8.405109e-10, 3.563121e-09, 3.362828e-09, 3.470065e-09, 3.270304e-09, 
    3.410171e-09, 2.81834e-09, 2.65565e-09, 1.978684e-09, 2.240262e-09, 
    1.83418e-09, 2.196492e-09, 2.129038e-09, 1.821786e-09, 2.175782e-09, 
    1.454815e-09, 1.92204e-09, 1.120742e-09, 1.515482e-09, 1.098604e-09, 
    1.167735e-09, 1.054806e-09, 9.600648e-10, 8.491841e-10, 6.675975e-10, 
    7.070842e-10, 5.714746e-10, 3.078819e-09, 2.845446e-09, 2.865526e-09, 
    2.633463e-09, 2.470322e-09, 2.140623e-09, 1.67622e-09, 1.841901e-09, 
    1.545722e-09, 1.490407e-09, 1.943715e-09, 1.655796e-09, 2.696234e-09, 
    2.504416e-09, 2.617486e-09, 3.059927e-09, 1.802747e-09, 2.391657e-09, 
    1.388076e-09, 1.645016e-09, 9.732082e-10, 1.277898e-09, 7.294659e-10, 
    5.535511e-10, 4.161848e-10, 2.868559e-10, 2.723371e-09, 2.875961e-09, 
    2.60676e-09, 2.263313e-09, 1.973485e-09, 1.628492e-09, 1.595694e-09, 
    1.536766e-09, 1.390995e-09, 1.275853e-09, 1.518419e-09, 1.248029e-09, 
    2.461231e-09, 1.756843e-09, 2.935106e-09, 2.536674e-09, 2.282665e-09, 
    2.391882e-09, 1.861519e-09, 1.749314e-09, 1.340106e-09, 1.542505e-09, 
    5.939846e-10, 9.40784e-10, 2.087635e-10, 3.449514e-10, 2.930614e-09, 
    2.723904e-09, 2.081946e-09, 2.372792e-09, 1.607046e-09, 1.44831e-09, 
    1.327333e-09, 1.182776e-09, 1.167847e-09, 1.088077e-09, 1.220785e-09, 
    1.093134e-09, 1.627805e-09, 1.371229e-09, 2.149507e-09, 1.938104e-09, 
    2.033528e-09, 2.141779e-09, 1.819718e-09, 1.514373e-09, 1.508295e-09, 
    1.418474e-09, 1.184752e-09, 1.604344e-09, 5.566412e-10, 1.116719e-09, 
    2.510092e-09, 2.16077e-09, 2.113801e-09, 2.242974e-09, 1.463724e-09, 
    1.720395e-09, 1.089981e-09, 1.241634e-09, 9.999538e-10, 1.115677e-09, 
    1.133422e-09, 1.29644e-09, 1.405463e-09, 1.708002e-09, 1.984366e-09, 
    2.223923e-09, 2.166567e-09, 1.909102e-09, 1.496914e-09, 1.166486e-09, 
    1.23418e-09, 1.017107e-09, 1.655939e-09, 1.362617e-09, 1.47143e-09, 
    1.199246e-09, 1.846438e-09, 1.283599e-09, 2.013078e-09, 1.940117e-09, 
    1.725776e-09, 1.34407e-09, 1.268145e-09, 1.190248e-09, 1.237931e-09, 
    1.487323e-09, 1.531168e-09, 1.730796e-09, 1.788829e-09, 1.955851e-09, 
    2.101843e-09, 1.968164e-09, 1.83409e-09, 1.487227e-09, 1.215061e-09, 
    9.587545e-10, 9.020898e-10, 6.620214e-10, 8.53633e-10, 5.542101e-10, 
    8.031686e-10, 4.090351e-10, 1.255142e-09, 8.114907e-10, 1.716437e-09, 
    1.596603e-09, 1.394354e-09, 9.969288e-10, 1.20044e-09, 9.649155e-10, 
    1.532907e-09, 1.900587e-09, 2.004625e-09, 2.208818e-09, 2.000113e-09, 
    2.016568e-09, 1.828705e-09, 1.887726e-09, 1.476539e-09, 1.688948e-09, 
    1.133861e-09, 9.6665e-10, 5.847878e-10, 4.096329e-10, 2.71329e-10, 
    2.218027e-10, 2.080312e-10, 2.02448e-10,
  4.175814e-13, 4.150199e-13, 4.154954e-13, 4.135916e-13, 4.146255e-13, 
    4.134109e-13, 4.170386e-13, 4.149241e-13, 4.162507e-13, 4.17339e-13, 
    4.103881e-13, 4.135108e-13, 4.077413e-13, 4.092984e-13, 4.057686e-13, 
    4.079697e-13, 4.053879e-13, 4.058249e-13, 4.045875e-13, 4.049186e-13, 
    4.03577e-13, 4.044409e-13, 4.030126e-13, 4.037695e-13, 4.036413e-13, 
    4.04472e-13, 4.128342e-13, 4.107447e-13, 4.129665e-13, 4.126496e-13, 
    4.127912e-13, 4.146035e-13, 4.155836e-13, 4.177895e-13, 4.173734e-13, 
    4.15761e-13, 4.125089e-13, 4.135525e-13, 4.110362e-13, 4.11089e-13, 
    4.087e-13, 4.097247e-13, 4.063116e-13, 4.071715e-13, 4.049044e-13, 
    4.054132e-13, 4.049274e-13, 4.050709e-13, 4.049255e-13, 4.056879e-13, 
    4.053508e-13, 4.060608e-13, 4.095263e-13, 4.08385e-13, 4.1212e-13, 
    4.148766e-13, 4.169415e-13, 4.185265e-13, 4.182962e-13, 4.178629e-13, 
    4.157519e-13, 4.139371e-13, 4.126594e-13, 4.118535e-13, 4.110966e-13, 
    4.090194e-13, 4.080443e-13, 4.061477e-13, 4.06462e-13, 4.059366e-13, 
    4.05466e-13, 4.047416e-13, 4.048553e-13, 4.045557e-13, 4.059501e-13, 
    4.049911e-13, 4.066465e-13, 4.061571e-13, 4.108964e-13, 4.13265e-13, 
    4.143761e-13, 4.154031e-13, 4.181206e-13, 4.162101e-13, 4.169449e-13, 
    4.152349e-13, 4.142152e-13, 4.147132e-13, 4.11832e-13, 4.128983e-13, 
    4.07989e-13, 4.098944e-13, 4.055193e-13, 4.063965e-13, 4.053236e-13, 
    4.058522e-13, 4.049698e-13, 4.057589e-13, 4.044481e-13, 4.04197e-13, 
    4.043673e-13, 4.037427e-13, 4.058053e-13, 4.049273e-13, 4.147273e-13, 
    4.146452e-13, 4.14267e-13, 4.159834e-13, 4.160931e-13, 4.17801e-13, 
    4.162754e-13, 4.156551e-13, 4.141577e-13, 4.133221e-13, 4.125615e-13, 
    4.110006e-13, 4.094299e-13, 4.075189e-13, 4.063366e-13, 4.056272e-13, 
    4.060546e-13, 4.056761e-13, 4.061004e-13, 4.063076e-13, 4.042897e-13, 
    4.053477e-13, 4.038277e-13, 4.039014e-13, 4.045488e-13, 4.03893e-13, 
    4.145877e-13, 4.150635e-13, 4.168023e-13, 4.1543e-13, 4.179945e-13, 
    4.165239e-13, 4.157186e-13, 4.128752e-13, 4.123044e-13, 4.117916e-13, 
    4.108247e-13, 4.096702e-13, 4.07867e-13, 4.065134e-13, 4.054395e-13, 
    4.055132e-13, 4.054872e-13, 4.052657e-13, 4.058275e-13, 4.051776e-13, 
    4.050743e-13, 4.053479e-13, 4.039113e-13, 4.042854e-13, 4.039029e-13, 
    4.041429e-13, 4.149076e-13, 4.141193e-13, 4.145414e-13, 4.13755e-13, 
    4.143057e-13, 4.119739e-13, 4.113322e-13, 4.086577e-13, 4.096919e-13, 
    4.080859e-13, 4.095189e-13, 4.092523e-13, 4.080368e-13, 4.094371e-13, 
    4.06583e-13, 4.084336e-13, 4.052572e-13, 4.068235e-13, 4.051693e-13, 
    4.054439e-13, 4.049952e-13, 4.046186e-13, 4.041774e-13, 4.034542e-13, 
    4.036116e-13, 4.030709e-13, 4.130007e-13, 4.120808e-13, 4.1216e-13, 
    4.112446e-13, 4.106007e-13, 4.092981e-13, 4.074604e-13, 4.081164e-13, 
    4.069434e-13, 4.067241e-13, 4.085194e-13, 4.073795e-13, 4.114923e-13, 
    4.107353e-13, 4.111816e-13, 4.129263e-13, 4.079614e-13, 4.1029e-13, 
    4.063184e-13, 4.073368e-13, 4.046708e-13, 4.058812e-13, 4.037007e-13, 
    4.029994e-13, 4.02451e-13, 4.019339e-13, 4.115994e-13, 4.122011e-13, 
    4.111392e-13, 4.09783e-13, 4.086371e-13, 4.072713e-13, 4.071414e-13, 
    4.069079e-13, 4.063299e-13, 4.058731e-13, 4.068352e-13, 4.057627e-13, 
    4.105648e-13, 4.077797e-13, 4.124343e-13, 4.108626e-13, 4.098595e-13, 
    4.102909e-13, 4.081941e-13, 4.077499e-13, 4.061281e-13, 4.069306e-13, 
    4.031607e-13, 4.045419e-13, 4.016214e-13, 4.021663e-13, 4.124166e-13, 
    4.116015e-13, 4.090661e-13, 4.102155e-13, 4.071864e-13, 4.065572e-13, 
    4.060774e-13, 4.055036e-13, 4.054443e-13, 4.051274e-13, 4.056545e-13, 
    4.051475e-13, 4.072686e-13, 4.062515e-13, 4.093332e-13, 4.084972e-13, 
    4.088746e-13, 4.093027e-13, 4.080286e-13, 4.068191e-13, 4.06795e-13, 
    4.064389e-13, 4.055115e-13, 4.071756e-13, 4.030117e-13, 4.052412e-13, 
    4.107577e-13, 4.093777e-13, 4.091921e-13, 4.097027e-13, 4.066183e-13, 
    4.076353e-13, 4.05135e-13, 4.057373e-13, 4.047772e-13, 4.052371e-13, 
    4.053076e-13, 4.059548e-13, 4.063873e-13, 4.075863e-13, 4.086802e-13, 
    4.096274e-13, 4.094007e-13, 4.083824e-13, 4.067499e-13, 4.054389e-13, 
    4.057077e-13, 4.048454e-13, 4.0738e-13, 4.062174e-13, 4.066489e-13, 
    4.05569e-13, 4.081344e-13, 4.059039e-13, 4.087937e-13, 4.085051e-13, 
    4.076567e-13, 4.061438e-13, 4.058425e-13, 4.055333e-13, 4.057226e-13, 
    4.067119e-13, 4.068857e-13, 4.076765e-13, 4.079063e-13, 4.085674e-13, 
    4.091448e-13, 4.086161e-13, 4.080855e-13, 4.067115e-13, 4.056318e-13, 
    4.046134e-13, 4.043879e-13, 4.03432e-13, 4.041952e-13, 4.03002e-13, 
    4.039942e-13, 4.024224e-13, 4.057909e-13, 4.040274e-13, 4.076197e-13, 
    4.07145e-13, 4.063433e-13, 4.047651e-13, 4.055737e-13, 4.046379e-13, 
    4.068926e-13, 4.083487e-13, 4.087603e-13, 4.095677e-13, 4.087425e-13, 
    4.088076e-13, 4.080642e-13, 4.082978e-13, 4.066691e-13, 4.075108e-13, 
    4.053093e-13, 4.046447e-13, 4.03124e-13, 4.024248e-13, 4.018718e-13, 
    4.016736e-13, 4.016184e-13, 4.015961e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 
    8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949653e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949653e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 
    8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949651e-07, 8.949652e-07, 8.94965e-07, 8.94965e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949654e-07, 8.949651e-07, 8.949652e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949653e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949654e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.780541e-16, 6.798939e-16, 6.795365e-16, 6.810191e-16, 6.80197e-16, 
    6.811675e-16, 6.784274e-16, 6.799667e-16, 6.789844e-16, 6.782201e-16, 
    6.838921e-16, 6.810853e-16, 6.868051e-16, 6.850182e-16, 6.895041e-16, 
    6.865268e-16, 6.901038e-16, 6.894189e-16, 6.914811e-16, 6.908906e-16, 
    6.935243e-16, 6.917535e-16, 6.948888e-16, 6.931019e-16, 6.933813e-16, 
    6.91695e-16, 6.81651e-16, 6.835427e-16, 6.815388e-16, 6.818087e-16, 
    6.816877e-16, 6.802138e-16, 6.794703e-16, 6.779137e-16, 6.781965e-16, 
    6.793399e-16, 6.819301e-16, 6.810516e-16, 6.832658e-16, 6.832158e-16, 
    6.856772e-16, 6.845678e-16, 6.886999e-16, 6.875267e-16, 6.909152e-16, 
    6.900637e-16, 6.908752e-16, 6.906292e-16, 6.908783e-16, 6.896292e-16, 
    6.901645e-16, 6.890651e-16, 6.847755e-16, 6.860371e-16, 6.822713e-16, 
    6.800023e-16, 6.784949e-16, 6.774241e-16, 6.775755e-16, 6.77864e-16, 
    6.793466e-16, 6.807399e-16, 6.818008e-16, 6.8251e-16, 6.832086e-16, 
    6.853201e-16, 6.864378e-16, 6.889368e-16, 6.884866e-16, 6.892496e-16, 
    6.899789e-16, 6.91202e-16, 6.910008e-16, 6.915393e-16, 6.892299e-16, 
    6.907649e-16, 6.882299e-16, 6.889236e-16, 6.833967e-16, 6.812887e-16, 
    6.803904e-16, 6.796052e-16, 6.776918e-16, 6.790133e-16, 6.784924e-16, 
    6.797317e-16, 6.805184e-16, 6.801294e-16, 6.825295e-16, 6.815967e-16, 
    6.86504e-16, 6.84392e-16, 6.898939e-16, 6.88579e-16, 6.902089e-16, 
    6.893775e-16, 6.908017e-16, 6.8952e-16, 6.917398e-16, 6.922226e-16, 
    6.918927e-16, 6.931603e-16, 6.894489e-16, 6.90875e-16, 6.801184e-16, 
    6.801819e-16, 6.804776e-16, 6.791773e-16, 6.790978e-16, 6.779059e-16, 
    6.789667e-16, 6.79418e-16, 6.805641e-16, 6.812413e-16, 6.81885e-16, 
    6.832994e-16, 6.848773e-16, 6.870819e-16, 6.886643e-16, 6.89724e-16, 
    6.890744e-16, 6.896479e-16, 6.890067e-16, 6.887062e-16, 6.920416e-16, 
    6.901694e-16, 6.92978e-16, 6.928228e-16, 6.915521e-16, 6.928403e-16, 
    6.802264e-16, 6.798613e-16, 6.785925e-16, 6.795855e-16, 6.777761e-16, 
    6.787889e-16, 6.793709e-16, 6.816158e-16, 6.82109e-16, 6.825658e-16, 
    6.834679e-16, 6.846246e-16, 6.866519e-16, 6.884141e-16, 6.900214e-16, 
    6.899037e-16, 6.899451e-16, 6.903038e-16, 6.89415e-16, 6.904497e-16, 
    6.906231e-16, 6.901694e-16, 6.92802e-16, 6.920503e-16, 6.928195e-16, 
    6.923302e-16, 6.799801e-16, 6.805944e-16, 6.802624e-16, 6.808865e-16, 
    6.804468e-16, 6.824011e-16, 6.829866e-16, 6.857243e-16, 6.846018e-16, 
    6.863885e-16, 6.847835e-16, 6.850679e-16, 6.864459e-16, 6.848704e-16, 
    6.883166e-16, 6.859802e-16, 6.903178e-16, 6.879867e-16, 6.904637e-16, 
    6.900145e-16, 6.907583e-16, 6.914241e-16, 6.922616e-16, 6.938052e-16, 
    6.93448e-16, 6.947383e-16, 6.815101e-16, 6.823061e-16, 6.822363e-16, 
    6.830692e-16, 6.836849e-16, 6.850189e-16, 6.87156e-16, 6.863527e-16, 
    6.878274e-16, 6.881231e-16, 6.858829e-16, 6.872584e-16, 6.828389e-16, 
    6.835533e-16, 6.831282e-16, 6.815727e-16, 6.865374e-16, 6.839911e-16, 
    6.886904e-16, 6.873133e-16, 6.913291e-16, 6.893328e-16, 6.932512e-16, 
    6.949225e-16, 6.964954e-16, 6.983296e-16, 6.827407e-16, 6.822e-16, 
    6.831684e-16, 6.845066e-16, 6.857483e-16, 6.873972e-16, 6.87566e-16, 
    6.878746e-16, 6.886741e-16, 6.893458e-16, 6.879718e-16, 6.895142e-16, 
    6.837183e-16, 6.867584e-16, 6.819952e-16, 6.834304e-16, 6.844279e-16, 
    6.839908e-16, 6.86261e-16, 6.867955e-16, 6.889657e-16, 6.878444e-16, 
    6.945098e-16, 6.915642e-16, 6.99726e-16, 6.974492e-16, 6.820109e-16, 
    6.82739e-16, 6.8527e-16, 6.840663e-16, 6.875074e-16, 6.883532e-16, 
    6.890408e-16, 6.899187e-16, 6.900137e-16, 6.905336e-16, 6.896814e-16, 
    6.905001e-16, 6.874007e-16, 6.887865e-16, 6.849814e-16, 6.859081e-16, 
    6.854819e-16, 6.850141e-16, 6.864575e-16, 6.879934e-16, 6.880268e-16, 
    6.885188e-16, 6.899036e-16, 6.875214e-16, 6.948885e-16, 6.903418e-16, 
    6.835326e-16, 6.849327e-16, 6.851332e-16, 6.845909e-16, 6.882684e-16, 
    6.869368e-16, 6.90521e-16, 6.895532e-16, 6.911388e-16, 6.90351e-16, 
    6.902351e-16, 6.892228e-16, 6.885922e-16, 6.869978e-16, 6.856995e-16, 
    6.846696e-16, 6.849093e-16, 6.860403e-16, 6.880874e-16, 6.90022e-16, 
    6.895984e-16, 6.910184e-16, 6.872581e-16, 6.888356e-16, 6.882259e-16, 
    6.898153e-16, 6.863313e-16, 6.892969e-16, 6.855722e-16, 6.858992e-16, 
    6.869104e-16, 6.889422e-16, 6.893922e-16, 6.898715e-16, 6.895759e-16, 
    6.881395e-16, 6.879043e-16, 6.868859e-16, 6.866043e-16, 6.85828e-16, 
    6.851848e-16, 6.857724e-16, 6.863891e-16, 6.881403e-16, 6.897165e-16, 
    6.914335e-16, 6.918536e-16, 6.938555e-16, 6.922253e-16, 6.949137e-16, 
    6.926272e-16, 6.965839e-16, 6.894694e-16, 6.92561e-16, 6.869565e-16, 
    6.875614e-16, 6.886542e-16, 6.911591e-16, 6.898079e-16, 6.913883e-16, 
    6.878951e-16, 6.860791e-16, 6.856096e-16, 6.847322e-16, 6.856297e-16, 
    6.855567e-16, 6.86415e-16, 6.861393e-16, 6.881984e-16, 6.870927e-16, 
    6.90232e-16, 6.91376e-16, 6.94603e-16, 6.965776e-16, 6.98586e-16, 
    6.994715e-16, 6.99741e-16, 6.998536e-16 ;

 CWDC_TO_LITR2C =
  5.153211e-16, 5.167194e-16, 5.164477e-16, 5.175746e-16, 5.169498e-16, 
    5.176873e-16, 5.156049e-16, 5.167747e-16, 5.160281e-16, 5.154473e-16, 
    5.19758e-16, 5.176249e-16, 5.219719e-16, 5.206138e-16, 5.240231e-16, 
    5.217604e-16, 5.244789e-16, 5.239583e-16, 5.255256e-16, 5.250768e-16, 
    5.270785e-16, 5.257327e-16, 5.281155e-16, 5.267575e-16, 5.269698e-16, 
    5.256882e-16, 5.180548e-16, 5.194925e-16, 5.179695e-16, 5.181746e-16, 
    5.180826e-16, 5.169625e-16, 5.163974e-16, 5.152144e-16, 5.154293e-16, 
    5.162983e-16, 5.182668e-16, 5.175992e-16, 5.19282e-16, 5.192441e-16, 
    5.211146e-16, 5.202716e-16, 5.234119e-16, 5.225203e-16, 5.250956e-16, 
    5.244484e-16, 5.250651e-16, 5.248782e-16, 5.250676e-16, 5.241182e-16, 
    5.24525e-16, 5.236895e-16, 5.204294e-16, 5.213882e-16, 5.185262e-16, 
    5.168017e-16, 5.156561e-16, 5.148423e-16, 5.149574e-16, 5.151767e-16, 
    5.163034e-16, 5.173623e-16, 5.181686e-16, 5.187076e-16, 5.192386e-16, 
    5.208433e-16, 5.216927e-16, 5.23592e-16, 5.232498e-16, 5.238297e-16, 
    5.24384e-16, 5.253135e-16, 5.251606e-16, 5.255699e-16, 5.238147e-16, 
    5.249813e-16, 5.230548e-16, 5.235819e-16, 5.193814e-16, 5.177794e-16, 
    5.170967e-16, 5.164999e-16, 5.150458e-16, 5.160501e-16, 5.156542e-16, 
    5.165961e-16, 5.17194e-16, 5.168984e-16, 5.187224e-16, 5.180135e-16, 
    5.21743e-16, 5.201379e-16, 5.243193e-16, 5.233201e-16, 5.245588e-16, 
    5.239269e-16, 5.250093e-16, 5.240352e-16, 5.257223e-16, 5.260891e-16, 
    5.258384e-16, 5.268018e-16, 5.239811e-16, 5.25065e-16, 5.1689e-16, 
    5.169382e-16, 5.17163e-16, 5.161747e-16, 5.161143e-16, 5.152085e-16, 
    5.160146e-16, 5.163577e-16, 5.172288e-16, 5.177434e-16, 5.182326e-16, 
    5.193075e-16, 5.205068e-16, 5.221823e-16, 5.233848e-16, 5.241903e-16, 
    5.236965e-16, 5.241324e-16, 5.236451e-16, 5.234167e-16, 5.259516e-16, 
    5.245288e-16, 5.266633e-16, 5.265453e-16, 5.255795e-16, 5.265586e-16, 
    5.169721e-16, 5.166946e-16, 5.157303e-16, 5.16485e-16, 5.151098e-16, 
    5.158795e-16, 5.163219e-16, 5.18028e-16, 5.184029e-16, 5.1875e-16, 
    5.194356e-16, 5.203147e-16, 5.218555e-16, 5.231947e-16, 5.244163e-16, 
    5.243268e-16, 5.243583e-16, 5.246309e-16, 5.239554e-16, 5.247418e-16, 
    5.248736e-16, 5.245288e-16, 5.265295e-16, 5.259583e-16, 5.265428e-16, 
    5.261709e-16, 5.167849e-16, 5.172517e-16, 5.169994e-16, 5.174738e-16, 
    5.171395e-16, 5.186249e-16, 5.190698e-16, 5.211505e-16, 5.202973e-16, 
    5.216552e-16, 5.204355e-16, 5.206516e-16, 5.216989e-16, 5.205015e-16, 
    5.231206e-16, 5.21345e-16, 5.246415e-16, 5.228699e-16, 5.247524e-16, 
    5.24411e-16, 5.249764e-16, 5.254823e-16, 5.261188e-16, 5.272919e-16, 
    5.270205e-16, 5.280011e-16, 5.179477e-16, 5.185526e-16, 5.184996e-16, 
    5.191326e-16, 5.196005e-16, 5.206143e-16, 5.222385e-16, 5.216281e-16, 
    5.227488e-16, 5.229735e-16, 5.21271e-16, 5.223164e-16, 5.189576e-16, 
    5.195005e-16, 5.191775e-16, 5.179953e-16, 5.217684e-16, 5.198332e-16, 
    5.234047e-16, 5.223581e-16, 5.254101e-16, 5.238929e-16, 5.268709e-16, 
    5.281411e-16, 5.293365e-16, 5.307305e-16, 5.18883e-16, 5.18472e-16, 
    5.19208e-16, 5.20225e-16, 5.211687e-16, 5.224219e-16, 5.225502e-16, 
    5.227847e-16, 5.233923e-16, 5.239028e-16, 5.228586e-16, 5.240308e-16, 
    5.196259e-16, 5.219364e-16, 5.183163e-16, 5.194071e-16, 5.201652e-16, 
    5.19833e-16, 5.215584e-16, 5.219646e-16, 5.236139e-16, 5.227617e-16, 
    5.278275e-16, 5.255888e-16, 5.317917e-16, 5.300614e-16, 5.183283e-16, 
    5.188817e-16, 5.208052e-16, 5.198904e-16, 5.225057e-16, 5.231485e-16, 
    5.23671e-16, 5.243382e-16, 5.244104e-16, 5.248055e-16, 5.241579e-16, 
    5.247801e-16, 5.224246e-16, 5.234778e-16, 5.205858e-16, 5.212901e-16, 
    5.209662e-16, 5.206107e-16, 5.217077e-16, 5.22875e-16, 5.229003e-16, 
    5.232743e-16, 5.243267e-16, 5.225163e-16, 5.281153e-16, 5.246597e-16, 
    5.194847e-16, 5.205488e-16, 5.207012e-16, 5.202891e-16, 5.23084e-16, 
    5.22072e-16, 5.24796e-16, 5.240604e-16, 5.252655e-16, 5.246668e-16, 
    5.245787e-16, 5.238094e-16, 5.2333e-16, 5.221183e-16, 5.211316e-16, 
    5.20349e-16, 5.20531e-16, 5.213907e-16, 5.229464e-16, 5.244167e-16, 
    5.240948e-16, 5.251739e-16, 5.223162e-16, 5.235151e-16, 5.230517e-16, 
    5.242597e-16, 5.216117e-16, 5.238656e-16, 5.210348e-16, 5.212834e-16, 
    5.220519e-16, 5.235961e-16, 5.239381e-16, 5.243024e-16, 5.240777e-16, 
    5.22986e-16, 5.228072e-16, 5.220333e-16, 5.218193e-16, 5.212293e-16, 
    5.207405e-16, 5.21187e-16, 5.216557e-16, 5.229866e-16, 5.241845e-16, 
    5.254894e-16, 5.258087e-16, 5.273302e-16, 5.260912e-16, 5.281344e-16, 
    5.263967e-16, 5.294037e-16, 5.239968e-16, 5.263463e-16, 5.22087e-16, 
    5.225466e-16, 5.233772e-16, 5.252809e-16, 5.24254e-16, 5.254551e-16, 
    5.228003e-16, 5.214201e-16, 5.210633e-16, 5.203964e-16, 5.210785e-16, 
    5.210231e-16, 5.216754e-16, 5.214658e-16, 5.230308e-16, 5.221905e-16, 
    5.245763e-16, 5.254458e-16, 5.278982e-16, 5.29399e-16, 5.309253e-16, 
    5.315984e-16, 5.318032e-16, 5.318887e-16 ;

 CWDC_TO_LITR3C =
  1.62733e-16, 1.631745e-16, 1.630888e-16, 1.634446e-16, 1.632473e-16, 
    1.634802e-16, 1.628226e-16, 1.63192e-16, 1.629562e-16, 1.627728e-16, 
    1.641341e-16, 1.634605e-16, 1.648332e-16, 1.644044e-16, 1.65481e-16, 
    1.647664e-16, 1.656249e-16, 1.654605e-16, 1.659555e-16, 1.658137e-16, 
    1.664458e-16, 1.660209e-16, 1.667733e-16, 1.663445e-16, 1.664115e-16, 
    1.660068e-16, 1.635962e-16, 1.640503e-16, 1.635693e-16, 1.636341e-16, 
    1.63605e-16, 1.632513e-16, 1.630729e-16, 1.626993e-16, 1.627672e-16, 
    1.630416e-16, 1.636632e-16, 1.634524e-16, 1.639838e-16, 1.639718e-16, 
    1.645625e-16, 1.642963e-16, 1.65288e-16, 1.650064e-16, 1.658197e-16, 
    1.656153e-16, 1.6581e-16, 1.65751e-16, 1.658108e-16, 1.65511e-16, 
    1.656395e-16, 1.653756e-16, 1.643461e-16, 1.646489e-16, 1.637451e-16, 
    1.632006e-16, 1.628388e-16, 1.625818e-16, 1.626181e-16, 1.626874e-16, 
    1.630432e-16, 1.633776e-16, 1.636322e-16, 1.638024e-16, 1.639701e-16, 
    1.644768e-16, 1.647451e-16, 1.653448e-16, 1.652368e-16, 1.654199e-16, 
    1.655949e-16, 1.658885e-16, 1.658402e-16, 1.659694e-16, 1.654152e-16, 
    1.657836e-16, 1.651752e-16, 1.653417e-16, 1.640152e-16, 1.635093e-16, 
    1.632937e-16, 1.631052e-16, 1.62646e-16, 1.629632e-16, 1.628382e-16, 
    1.631356e-16, 1.633244e-16, 1.632311e-16, 1.638071e-16, 1.635832e-16, 
    1.647609e-16, 1.642541e-16, 1.655745e-16, 1.65259e-16, 1.656501e-16, 
    1.654506e-16, 1.657924e-16, 1.654848e-16, 1.660176e-16, 1.661334e-16, 
    1.660542e-16, 1.663585e-16, 1.654677e-16, 1.6581e-16, 1.632284e-16, 
    1.632436e-16, 1.633146e-16, 1.630025e-16, 1.629835e-16, 1.626974e-16, 
    1.62952e-16, 1.630603e-16, 1.633354e-16, 1.634979e-16, 1.636524e-16, 
    1.639919e-16, 1.643706e-16, 1.648997e-16, 1.652794e-16, 1.655338e-16, 
    1.653779e-16, 1.655155e-16, 1.653616e-16, 1.652895e-16, 1.6609e-16, 
    1.656407e-16, 1.663147e-16, 1.662775e-16, 1.659725e-16, 1.662817e-16, 
    1.632543e-16, 1.631667e-16, 1.628622e-16, 1.631005e-16, 1.626662e-16, 
    1.629093e-16, 1.63049e-16, 1.635878e-16, 1.637062e-16, 1.638158e-16, 
    1.640323e-16, 1.643099e-16, 1.647965e-16, 1.652194e-16, 1.656051e-16, 
    1.655769e-16, 1.655868e-16, 1.656729e-16, 1.654596e-16, 1.657079e-16, 
    1.657496e-16, 1.656407e-16, 1.662725e-16, 1.660921e-16, 1.662767e-16, 
    1.661592e-16, 1.631952e-16, 1.633427e-16, 1.63263e-16, 1.634128e-16, 
    1.633072e-16, 1.637763e-16, 1.639168e-16, 1.645738e-16, 1.643044e-16, 
    1.647332e-16, 1.64348e-16, 1.644163e-16, 1.64747e-16, 1.643689e-16, 
    1.65196e-16, 1.646353e-16, 1.656763e-16, 1.651168e-16, 1.657113e-16, 
    1.656035e-16, 1.65782e-16, 1.659418e-16, 1.661428e-16, 1.665132e-16, 
    1.664275e-16, 1.667372e-16, 1.635624e-16, 1.637535e-16, 1.637367e-16, 
    1.639366e-16, 1.640844e-16, 1.644045e-16, 1.649174e-16, 1.647247e-16, 
    1.650786e-16, 1.651495e-16, 1.646119e-16, 1.64942e-16, 1.638813e-16, 
    1.640528e-16, 1.639508e-16, 1.635775e-16, 1.64769e-16, 1.641579e-16, 
    1.652857e-16, 1.649552e-16, 1.65919e-16, 1.654399e-16, 1.663803e-16, 
    1.667814e-16, 1.671589e-16, 1.675991e-16, 1.638578e-16, 1.63728e-16, 
    1.639604e-16, 1.642816e-16, 1.645796e-16, 1.649753e-16, 1.650158e-16, 
    1.650899e-16, 1.652818e-16, 1.65443e-16, 1.651132e-16, 1.654834e-16, 
    1.640924e-16, 1.64822e-16, 1.636788e-16, 1.640233e-16, 1.642627e-16, 
    1.641578e-16, 1.647026e-16, 1.648309e-16, 1.653518e-16, 1.650827e-16, 
    1.666824e-16, 1.659754e-16, 1.679342e-16, 1.673878e-16, 1.636826e-16, 
    1.638574e-16, 1.644648e-16, 1.641759e-16, 1.650018e-16, 1.652048e-16, 
    1.653698e-16, 1.655805e-16, 1.656033e-16, 1.657281e-16, 1.655236e-16, 
    1.6572e-16, 1.649762e-16, 1.653088e-16, 1.643955e-16, 1.646179e-16, 
    1.645157e-16, 1.644034e-16, 1.647498e-16, 1.651184e-16, 1.651264e-16, 
    1.652445e-16, 1.655769e-16, 1.650051e-16, 1.667732e-16, 1.65682e-16, 
    1.640478e-16, 1.643838e-16, 1.64432e-16, 1.643018e-16, 1.651844e-16, 
    1.648648e-16, 1.65725e-16, 1.654928e-16, 1.658733e-16, 1.656843e-16, 
    1.656564e-16, 1.654135e-16, 1.652621e-16, 1.648795e-16, 1.645679e-16, 
    1.643207e-16, 1.643782e-16, 1.646497e-16, 1.65141e-16, 1.656053e-16, 
    1.655036e-16, 1.658444e-16, 1.64942e-16, 1.653205e-16, 1.651742e-16, 
    1.655557e-16, 1.647195e-16, 1.654313e-16, 1.645373e-16, 1.646158e-16, 
    1.648585e-16, 1.653461e-16, 1.654541e-16, 1.655692e-16, 1.654982e-16, 
    1.651535e-16, 1.65097e-16, 1.648526e-16, 1.64785e-16, 1.645987e-16, 
    1.644444e-16, 1.645854e-16, 1.647334e-16, 1.651537e-16, 1.65532e-16, 
    1.65944e-16, 1.660449e-16, 1.665253e-16, 1.661341e-16, 1.667793e-16, 
    1.662305e-16, 1.671801e-16, 1.654727e-16, 1.662146e-16, 1.648696e-16, 
    1.650147e-16, 1.65277e-16, 1.658782e-16, 1.655539e-16, 1.659332e-16, 
    1.650948e-16, 1.64659e-16, 1.645463e-16, 1.643357e-16, 1.645511e-16, 
    1.645336e-16, 1.647396e-16, 1.646734e-16, 1.651676e-16, 1.649023e-16, 
    1.656557e-16, 1.659302e-16, 1.667047e-16, 1.671786e-16, 1.676606e-16, 
    1.678732e-16, 1.679378e-16, 1.679649e-16 ;

 CWDC_vr =
  5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110343e-05, 5.110344e-05, 5.110342e-05, 5.110343e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110343e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  1.030642e-18, 1.033439e-18, 1.032896e-18, 1.035149e-18, 1.0339e-18, 
    1.035375e-18, 1.03121e-18, 1.033549e-18, 1.032056e-18, 1.030895e-18, 
    1.039516e-18, 1.03525e-18, 1.043944e-18, 1.041228e-18, 1.048046e-18, 
    1.043521e-18, 1.048958e-18, 1.047917e-18, 1.051051e-18, 1.050154e-18, 
    1.054157e-18, 1.051465e-18, 1.056231e-18, 1.053515e-18, 1.05394e-18, 
    1.051376e-18, 1.03611e-18, 1.038985e-18, 1.035939e-18, 1.036349e-18, 
    1.036165e-18, 1.033925e-18, 1.032795e-18, 1.030429e-18, 1.030859e-18, 
    1.032597e-18, 1.036534e-18, 1.035198e-18, 1.038564e-18, 1.038488e-18, 
    1.042229e-18, 1.040543e-18, 1.046824e-18, 1.045041e-18, 1.050191e-18, 
    1.048897e-18, 1.05013e-18, 1.049756e-18, 1.050135e-18, 1.048236e-18, 
    1.04905e-18, 1.047379e-18, 1.040859e-18, 1.042776e-18, 1.037052e-18, 
    1.033604e-18, 1.031312e-18, 1.029685e-18, 1.029915e-18, 1.030353e-18, 
    1.032607e-18, 1.034725e-18, 1.036337e-18, 1.037415e-18, 1.038477e-18, 
    1.041687e-18, 1.043385e-18, 1.047184e-18, 1.0465e-18, 1.047659e-18, 
    1.048768e-18, 1.050627e-18, 1.050321e-18, 1.05114e-18, 1.047629e-18, 
    1.049963e-18, 1.046109e-18, 1.047164e-18, 1.038763e-18, 1.035559e-18, 
    1.034193e-18, 1.033e-18, 1.030092e-18, 1.0321e-18, 1.031309e-18, 
    1.033192e-18, 1.034388e-18, 1.033797e-18, 1.037445e-18, 1.036027e-18, 
    1.043486e-18, 1.040276e-18, 1.048639e-18, 1.04664e-18, 1.049118e-18, 
    1.047854e-18, 1.050019e-18, 1.04807e-18, 1.051445e-18, 1.052178e-18, 
    1.051677e-18, 1.053604e-18, 1.047962e-18, 1.05013e-18, 1.03378e-18, 
    1.033876e-18, 1.034326e-18, 1.032349e-18, 1.032229e-18, 1.030417e-18, 
    1.032029e-18, 1.032715e-18, 1.034457e-18, 1.035487e-18, 1.036465e-18, 
    1.038615e-18, 1.041014e-18, 1.044365e-18, 1.04677e-18, 1.04838e-18, 
    1.047393e-18, 1.048265e-18, 1.04729e-18, 1.046833e-18, 1.051903e-18, 
    1.049057e-18, 1.053327e-18, 1.053091e-18, 1.051159e-18, 1.053117e-18, 
    1.033944e-18, 1.033389e-18, 1.031461e-18, 1.03297e-18, 1.03022e-18, 
    1.031759e-18, 1.032644e-18, 1.036056e-18, 1.036806e-18, 1.0375e-18, 
    1.038871e-18, 1.040629e-18, 1.043711e-18, 1.046389e-18, 1.048833e-18, 
    1.048654e-18, 1.048717e-18, 1.049262e-18, 1.047911e-18, 1.049484e-18, 
    1.049747e-18, 1.049057e-18, 1.053059e-18, 1.051916e-18, 1.053086e-18, 
    1.052342e-18, 1.03357e-18, 1.034504e-18, 1.033999e-18, 1.034948e-18, 
    1.034279e-18, 1.03725e-18, 1.03814e-18, 1.042301e-18, 1.040595e-18, 
    1.04331e-18, 1.040871e-18, 1.041303e-18, 1.043398e-18, 1.041003e-18, 
    1.046241e-18, 1.04269e-18, 1.049283e-18, 1.04574e-18, 1.049505e-18, 
    1.048822e-18, 1.049953e-18, 1.050965e-18, 1.052238e-18, 1.054584e-18, 
    1.054041e-18, 1.056002e-18, 1.035895e-18, 1.037105e-18, 1.036999e-18, 
    1.038265e-18, 1.039201e-18, 1.041229e-18, 1.044477e-18, 1.043256e-18, 
    1.045498e-18, 1.045947e-18, 1.042542e-18, 1.044633e-18, 1.037915e-18, 
    1.039001e-18, 1.038355e-18, 1.03599e-18, 1.043537e-18, 1.039666e-18, 
    1.046809e-18, 1.044716e-18, 1.05082e-18, 1.047786e-18, 1.053742e-18, 
    1.056282e-18, 1.058673e-18, 1.061461e-18, 1.037766e-18, 1.036944e-18, 
    1.038416e-18, 1.04045e-18, 1.042337e-18, 1.044844e-18, 1.0451e-18, 
    1.045569e-18, 1.046785e-18, 1.047806e-18, 1.045717e-18, 1.048062e-18, 
    1.039252e-18, 1.043873e-18, 1.036633e-18, 1.038814e-18, 1.04033e-18, 
    1.039666e-18, 1.043117e-18, 1.043929e-18, 1.047228e-18, 1.045524e-18, 
    1.055655e-18, 1.051178e-18, 1.063584e-18, 1.060123e-18, 1.036657e-18, 
    1.037763e-18, 1.04161e-18, 1.039781e-18, 1.045011e-18, 1.046297e-18, 
    1.047342e-18, 1.048676e-18, 1.048821e-18, 1.049611e-18, 1.048316e-18, 
    1.04956e-18, 1.044849e-18, 1.046956e-18, 1.041172e-18, 1.04258e-18, 
    1.041933e-18, 1.041221e-18, 1.043415e-18, 1.04575e-18, 1.045801e-18, 
    1.046549e-18, 1.048653e-18, 1.045032e-18, 1.056231e-18, 1.049319e-18, 
    1.038969e-18, 1.041098e-18, 1.041403e-18, 1.040578e-18, 1.046168e-18, 
    1.044144e-18, 1.049592e-18, 1.048121e-18, 1.050531e-18, 1.049334e-18, 
    1.049157e-18, 1.047619e-18, 1.04666e-18, 1.044237e-18, 1.042263e-18, 
    1.040698e-18, 1.041062e-18, 1.042781e-18, 1.045893e-18, 1.048833e-18, 
    1.04819e-18, 1.050348e-18, 1.044632e-18, 1.04703e-18, 1.046103e-18, 
    1.048519e-18, 1.043224e-18, 1.047731e-18, 1.04207e-18, 1.042567e-18, 
    1.044104e-18, 1.047192e-18, 1.047876e-18, 1.048605e-18, 1.048155e-18, 
    1.045972e-18, 1.045614e-18, 1.044067e-18, 1.043639e-18, 1.042459e-18, 
    1.041481e-18, 1.042374e-18, 1.043311e-18, 1.045973e-18, 1.048369e-18, 
    1.050979e-18, 1.051617e-18, 1.05466e-18, 1.052182e-18, 1.056269e-18, 
    1.052793e-18, 1.058807e-18, 1.047994e-18, 1.052693e-18, 1.044174e-18, 
    1.045093e-18, 1.046754e-18, 1.050562e-18, 1.048508e-18, 1.05091e-18, 
    1.045601e-18, 1.04284e-18, 1.042127e-18, 1.040793e-18, 1.042157e-18, 
    1.042046e-18, 1.043351e-18, 1.042932e-18, 1.046062e-18, 1.044381e-18, 
    1.049153e-18, 1.050892e-18, 1.055796e-18, 1.058798e-18, 1.061851e-18, 
    1.063197e-18, 1.063606e-18, 1.063778e-18 ;

 CWDN_TO_LITR3N =
  3.254659e-19, 3.263491e-19, 3.261775e-19, 3.268892e-19, 3.264946e-19, 
    3.269604e-19, 3.256452e-19, 3.26384e-19, 3.259125e-19, 3.255456e-19, 
    3.282682e-19, 3.26921e-19, 3.296664e-19, 3.288087e-19, 3.309619e-19, 
    3.295329e-19, 3.312499e-19, 3.30921e-19, 3.319109e-19, 3.316275e-19, 
    3.328917e-19, 3.320417e-19, 3.335466e-19, 3.326889e-19, 3.32823e-19, 
    3.320136e-19, 3.271925e-19, 3.281005e-19, 3.271386e-19, 3.272682e-19, 
    3.272101e-19, 3.265026e-19, 3.261457e-19, 3.253986e-19, 3.255343e-19, 
    3.260832e-19, 3.273264e-19, 3.269048e-19, 3.279676e-19, 3.279436e-19, 
    3.29125e-19, 3.285926e-19, 3.30576e-19, 3.300128e-19, 3.316393e-19, 
    3.312305e-19, 3.316201e-19, 3.31502e-19, 3.316216e-19, 3.31022e-19, 
    3.31279e-19, 3.307512e-19, 3.286923e-19, 3.292978e-19, 3.274902e-19, 
    3.264011e-19, 3.256776e-19, 3.251636e-19, 3.252362e-19, 3.253747e-19, 
    3.260864e-19, 3.267552e-19, 3.272644e-19, 3.276048e-19, 3.279401e-19, 
    3.289536e-19, 3.294901e-19, 3.306897e-19, 3.304736e-19, 3.308398e-19, 
    3.311899e-19, 3.317769e-19, 3.316804e-19, 3.319389e-19, 3.308303e-19, 
    3.315672e-19, 3.303504e-19, 3.306833e-19, 3.280304e-19, 3.270186e-19, 
    3.265874e-19, 3.262105e-19, 3.252921e-19, 3.259264e-19, 3.256764e-19, 
    3.262712e-19, 3.266488e-19, 3.264621e-19, 3.276141e-19, 3.271664e-19, 
    3.295219e-19, 3.285082e-19, 3.311491e-19, 3.305179e-19, 3.313003e-19, 
    3.309012e-19, 3.315848e-19, 3.309696e-19, 3.320351e-19, 3.322668e-19, 
    3.321085e-19, 3.327169e-19, 3.309355e-19, 3.3162e-19, 3.264568e-19, 
    3.264873e-19, 3.266292e-19, 3.260051e-19, 3.259669e-19, 3.253948e-19, 
    3.25904e-19, 3.261207e-19, 3.266708e-19, 3.269958e-19, 3.273048e-19, 
    3.279837e-19, 3.287411e-19, 3.297993e-19, 3.305588e-19, 3.310675e-19, 
    3.307557e-19, 3.31031e-19, 3.307232e-19, 3.30579e-19, 3.3218e-19, 
    3.312813e-19, 3.326294e-19, 3.325549e-19, 3.31945e-19, 3.325633e-19, 
    3.265087e-19, 3.263334e-19, 3.257244e-19, 3.262011e-19, 3.253325e-19, 
    3.258187e-19, 3.26098e-19, 3.271756e-19, 3.274123e-19, 3.276316e-19, 
    3.280646e-19, 3.286198e-19, 3.295929e-19, 3.304388e-19, 3.312103e-19, 
    3.311538e-19, 3.311737e-19, 3.313458e-19, 3.309192e-19, 3.314159e-19, 
    3.314991e-19, 3.312813e-19, 3.32545e-19, 3.321842e-19, 3.325534e-19, 
    3.323185e-19, 3.263904e-19, 3.266853e-19, 3.26526e-19, 3.268255e-19, 
    3.266144e-19, 3.275525e-19, 3.278336e-19, 3.291477e-19, 3.286088e-19, 
    3.294665e-19, 3.286961e-19, 3.288326e-19, 3.294941e-19, 3.287378e-19, 
    3.30392e-19, 3.292705e-19, 3.313525e-19, 3.302336e-19, 3.314226e-19, 
    3.312069e-19, 3.31564e-19, 3.318836e-19, 3.322856e-19, 3.330265e-19, 
    3.32855e-19, 3.334744e-19, 3.271248e-19, 3.275069e-19, 3.274734e-19, 
    3.278733e-19, 3.281687e-19, 3.288091e-19, 3.298349e-19, 3.294493e-19, 
    3.301571e-19, 3.302991e-19, 3.292238e-19, 3.29884e-19, 3.277627e-19, 
    3.281056e-19, 3.279016e-19, 3.271549e-19, 3.295379e-19, 3.283157e-19, 
    3.305714e-19, 3.299104e-19, 3.31838e-19, 3.308798e-19, 3.327606e-19, 
    3.335628e-19, 3.343178e-19, 3.351982e-19, 3.277155e-19, 3.27456e-19, 
    3.279208e-19, 3.285632e-19, 3.291592e-19, 3.299507e-19, 3.300317e-19, 
    3.301798e-19, 3.305636e-19, 3.30886e-19, 3.302265e-19, 3.309668e-19, 
    3.281848e-19, 3.29644e-19, 3.273577e-19, 3.280466e-19, 3.285254e-19, 
    3.283156e-19, 3.294053e-19, 3.296619e-19, 3.307035e-19, 3.301653e-19, 
    3.333647e-19, 3.319508e-19, 3.358685e-19, 3.347756e-19, 3.273653e-19, 
    3.277147e-19, 3.289296e-19, 3.283518e-19, 3.300036e-19, 3.304095e-19, 
    3.307396e-19, 3.31161e-19, 3.312066e-19, 3.314561e-19, 3.310471e-19, 
    3.314401e-19, 3.299523e-19, 3.306176e-19, 3.28791e-19, 3.292359e-19, 
    3.290313e-19, 3.288068e-19, 3.294996e-19, 3.302368e-19, 3.302528e-19, 
    3.30489e-19, 3.311537e-19, 3.300103e-19, 3.335465e-19, 3.31364e-19, 
    3.280956e-19, 3.287677e-19, 3.288639e-19, 3.286037e-19, 3.303688e-19, 
    3.297297e-19, 3.314501e-19, 3.309855e-19, 3.317466e-19, 3.313685e-19, 
    3.313128e-19, 3.30827e-19, 3.305242e-19, 3.297589e-19, 3.291358e-19, 
    3.286414e-19, 3.287564e-19, 3.292994e-19, 3.302819e-19, 3.312106e-19, 
    3.310072e-19, 3.316888e-19, 3.298839e-19, 3.306411e-19, 3.303484e-19, 
    3.311114e-19, 3.29439e-19, 3.308625e-19, 3.290747e-19, 3.292316e-19, 
    3.29717e-19, 3.306922e-19, 3.309083e-19, 3.311383e-19, 3.309964e-19, 
    3.303069e-19, 3.30194e-19, 3.297052e-19, 3.295701e-19, 3.291975e-19, 
    3.288887e-19, 3.291707e-19, 3.294668e-19, 3.303073e-19, 3.310639e-19, 
    3.318881e-19, 3.320897e-19, 3.330506e-19, 3.322681e-19, 3.335586e-19, 
    3.324611e-19, 3.343603e-19, 3.309453e-19, 3.324293e-19, 3.297391e-19, 
    3.300295e-19, 3.30554e-19, 3.317564e-19, 3.311078e-19, 3.318664e-19, 
    3.301896e-19, 3.293179e-19, 3.290926e-19, 3.286715e-19, 3.291022e-19, 
    3.290672e-19, 3.294792e-19, 3.293468e-19, 3.303352e-19, 3.298045e-19, 
    3.313114e-19, 3.318605e-19, 3.334094e-19, 3.343572e-19, 3.353213e-19, 
    3.357463e-19, 3.358757e-19, 3.359297e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.194416e-08, 6.221921e-08, 6.216575e-08, 6.238761e-08, 6.226454e-08, 
    6.240981e-08, 6.199993e-08, 6.223013e-08, 6.208317e-08, 6.196893e-08, 
    6.281821e-08, 6.239751e-08, 6.325536e-08, 6.298698e-08, 6.366125e-08, 
    6.321359e-08, 6.375153e-08, 6.364835e-08, 6.395895e-08, 6.386996e-08, 
    6.426725e-08, 6.400002e-08, 6.447324e-08, 6.420344e-08, 6.424563e-08, 
    6.39912e-08, 6.248218e-08, 6.276583e-08, 6.246538e-08, 6.250582e-08, 
    6.248767e-08, 6.226708e-08, 6.215591e-08, 6.192315e-08, 6.19654e-08, 
    6.213637e-08, 6.2524e-08, 6.239242e-08, 6.272409e-08, 6.27166e-08, 
    6.308589e-08, 6.291938e-08, 6.354018e-08, 6.336372e-08, 6.387368e-08, 
    6.374542e-08, 6.386765e-08, 6.383059e-08, 6.386814e-08, 6.368003e-08, 
    6.376062e-08, 6.359511e-08, 6.295056e-08, 6.313996e-08, 6.25751e-08, 
    6.223551e-08, 6.201002e-08, 6.185e-08, 6.187263e-08, 6.191575e-08, 
    6.213737e-08, 6.234576e-08, 6.250459e-08, 6.261083e-08, 6.271553e-08, 
    6.303241e-08, 6.320018e-08, 6.357585e-08, 6.350807e-08, 6.362291e-08, 
    6.373266e-08, 6.39169e-08, 6.388658e-08, 6.396775e-08, 6.361989e-08, 
    6.385107e-08, 6.346945e-08, 6.357381e-08, 6.274394e-08, 6.242792e-08, 
    6.229357e-08, 6.217602e-08, 6.189002e-08, 6.208752e-08, 6.200966e-08, 
    6.219491e-08, 6.231262e-08, 6.22544e-08, 6.261374e-08, 6.247403e-08, 
    6.321012e-08, 6.289304e-08, 6.371985e-08, 6.352198e-08, 6.376729e-08, 
    6.364211e-08, 6.38566e-08, 6.366356e-08, 6.399797e-08, 6.407078e-08, 
    6.402102e-08, 6.421219e-08, 6.365286e-08, 6.386765e-08, 6.225277e-08, 
    6.226226e-08, 6.23065e-08, 6.211204e-08, 6.210015e-08, 6.192198e-08, 
    6.208052e-08, 6.214803e-08, 6.231944e-08, 6.242083e-08, 6.251722e-08, 
    6.272915e-08, 6.296587e-08, 6.329692e-08, 6.353481e-08, 6.369427e-08, 
    6.359649e-08, 6.368282e-08, 6.358631e-08, 6.354109e-08, 6.40435e-08, 
    6.376137e-08, 6.41847e-08, 6.416128e-08, 6.396969e-08, 6.416391e-08, 
    6.226892e-08, 6.221429e-08, 6.202459e-08, 6.217304e-08, 6.190258e-08, 
    6.205396e-08, 6.214101e-08, 6.247694e-08, 6.255076e-08, 6.26192e-08, 
    6.27544e-08, 6.29279e-08, 6.32323e-08, 6.349719e-08, 6.373904e-08, 
    6.372132e-08, 6.372756e-08, 6.378159e-08, 6.364776e-08, 6.380356e-08, 
    6.38297e-08, 6.376134e-08, 6.415814e-08, 6.404477e-08, 6.416078e-08, 
    6.408697e-08, 6.223205e-08, 6.232399e-08, 6.227431e-08, 6.236773e-08, 
    6.230191e-08, 6.259458e-08, 6.268234e-08, 6.309303e-08, 6.292449e-08, 
    6.319274e-08, 6.295173e-08, 6.299444e-08, 6.320148e-08, 6.296477e-08, 
    6.348257e-08, 6.313149e-08, 6.378369e-08, 6.343302e-08, 6.380566e-08, 
    6.3738e-08, 6.385004e-08, 6.395038e-08, 6.407663e-08, 6.430958e-08, 
    6.425564e-08, 6.445048e-08, 6.246106e-08, 6.258032e-08, 6.256982e-08, 
    6.269464e-08, 6.278695e-08, 6.298706e-08, 6.330801e-08, 6.318732e-08, 
    6.340892e-08, 6.345341e-08, 6.311675e-08, 6.332343e-08, 6.266014e-08, 
    6.276728e-08, 6.27035e-08, 6.247047e-08, 6.321512e-08, 6.283292e-08, 
    6.353874e-08, 6.333165e-08, 6.393607e-08, 6.363545e-08, 6.422594e-08, 
    6.447839e-08, 6.471606e-08, 6.499378e-08, 6.264541e-08, 6.256438e-08, 
    6.270949e-08, 6.291025e-08, 6.309657e-08, 6.334428e-08, 6.336963e-08, 
    6.341604e-08, 6.353626e-08, 6.363734e-08, 6.34307e-08, 6.366268e-08, 
    6.279212e-08, 6.32483e-08, 6.253374e-08, 6.274887e-08, 6.289842e-08, 
    6.283283e-08, 6.317353e-08, 6.325383e-08, 6.358018e-08, 6.341148e-08, 
    6.441608e-08, 6.397156e-08, 6.52053e-08, 6.486045e-08, 6.253607e-08, 
    6.264514e-08, 6.302479e-08, 6.284415e-08, 6.336082e-08, 6.348802e-08, 
    6.359143e-08, 6.372361e-08, 6.373789e-08, 6.381621e-08, 6.368786e-08, 
    6.381114e-08, 6.334481e-08, 6.355319e-08, 6.298141e-08, 6.312055e-08, 
    6.305654e-08, 6.298632e-08, 6.320305e-08, 6.343395e-08, 6.34389e-08, 
    6.351294e-08, 6.372157e-08, 6.336292e-08, 6.447343e-08, 6.378752e-08, 
    6.276409e-08, 6.297419e-08, 6.300422e-08, 6.292283e-08, 6.347526e-08, 
    6.327508e-08, 6.38143e-08, 6.366856e-08, 6.390736e-08, 6.37887e-08, 
    6.377123e-08, 6.361883e-08, 6.352395e-08, 6.328425e-08, 6.308925e-08, 
    6.293464e-08, 6.297059e-08, 6.314043e-08, 6.344808e-08, 6.373917e-08, 
    6.367541e-08, 6.388921e-08, 6.332336e-08, 6.356061e-08, 6.34689e-08, 
    6.370803e-08, 6.318411e-08, 6.36302e-08, 6.307009e-08, 6.31192e-08, 
    6.327111e-08, 6.357669e-08, 6.364433e-08, 6.371651e-08, 6.367197e-08, 
    6.34559e-08, 6.34205e-08, 6.326741e-08, 6.322514e-08, 6.310851e-08, 
    6.301195e-08, 6.310017e-08, 6.319282e-08, 6.345599e-08, 6.369318e-08, 
    6.39518e-08, 6.401511e-08, 6.431729e-08, 6.407128e-08, 6.447725e-08, 
    6.413207e-08, 6.472964e-08, 6.365608e-08, 6.412193e-08, 6.327802e-08, 
    6.336893e-08, 6.353335e-08, 6.391052e-08, 6.370691e-08, 6.394504e-08, 
    6.341912e-08, 6.314629e-08, 6.307572e-08, 6.294403e-08, 6.307872e-08, 
    6.306777e-08, 6.319667e-08, 6.315525e-08, 6.346473e-08, 6.329849e-08, 
    6.377079e-08, 6.394317e-08, 6.443005e-08, 6.472857e-08, 6.503251e-08, 
    6.51667e-08, 6.520754e-08, 6.522462e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -1.419495e-14, -1.451915e-14, -1.121135e-14, -9.590271e-15, -1.28268e-14, 
    -5.888992e-15, -1.194167e-14, -1.625317e-14, -3.191106e-15, 
    -1.195784e-14, -1.217117e-14, -1.755472e-14, -1.890472e-14, 
    -8.739503e-15, -3.984805e-15, -6.550426e-15, -1.864371e-14, 
    -1.515054e-14, -1.008338e-14, -4.607991e-15, -8.087831e-15, 
    -1.124913e-14, -1.39672e-14, -1.183647e-14, -1.200807e-14, -1.006721e-14, 
    -1.055797e-14, -1.596014e-14, -1.265971e-14, -1.12871e-14, -9.839363e-15, 
    -1.163318e-14, -9.350558e-15, -1.667478e-14, -1.315719e-14, 
    -1.821757e-14, -1.245493e-14, -1.733935e-14, -6.148343e-15, 
    -1.601207e-14, -9.883712e-15, -1.547859e-14, -8.636446e-15, 
    -1.406236e-14, -1.037998e-14, -1.246067e-14, -1.925942e-14, 
    -7.858807e-15, -1.185932e-14, -7.302578e-15, -9.236505e-15, 
    -1.429329e-14, -1.300217e-14, -1.091151e-14, -1.083409e-14, -3.78757e-15, 
    -1.05121e-14, -1.546679e-14, -2.20615e-14, -1.818588e-14, -9.202684e-15, 
    -1.054834e-14, -1.31546e-14, -1.574289e-14, -1.722188e-14, -1.60629e-14, 
    -1.084803e-14, -1.004326e-14, -1.205331e-14, -1.673657e-14, 
    -1.426597e-14, -1.905935e-14, -1.260102e-14, -1.255685e-14, 
    -6.499333e-15, -1.489051e-14, -9.051874e-15, -1.375698e-14, -1.2214e-14, 
    -1.065473e-14, -1.484765e-14, -1.122333e-14, -1.018246e-14, 
    -1.627617e-14, -1.215594e-14, -1.64944e-14, -1.821267e-14, -1.29102e-14, 
    -9.318617e-15, -2.32524e-14, -9.518551e-15, -1.132769e-14, -1.776684e-14, 
    -1.130577e-14, -1.09023e-14, -1.923679e-14, -2.051789e-14, -6.36654e-15, 
    -8.63215e-15, -4.778035e-15, -7.543826e-15, -1.405478e-14, -1.028909e-14, 
    -1.070292e-14, -9.201198e-15, -1.293708e-14, -1.130389e-14, 
    -1.228531e-14, -1.281276e-14, -1.824778e-14, -1.570136e-14, 
    -1.365862e-14, -1.059289e-14, -9.934957e-15, -1.000067e-14, 
    -1.143888e-14, -1.289164e-14, -1.318386e-14, -1.884495e-14, 
    -1.152108e-14, -1.035161e-14, -1.55635e-14, -1.685e-14, -7.396141e-15, 
    -1.390752e-14, -1.143001e-14, -6.932783e-15, -1.006153e-14, 
    -9.604219e-15, -1.021666e-14, -1.336932e-14, -9.692001e-15, -6.35128e-15, 
    -1.490622e-14, -1.122516e-14, -8.279674e-15, -1.493594e-14, 
    -1.763833e-14, -1.566707e-14, -1.82333e-14, -5.354761e-15, -1.294359e-14, 
    -8.646805e-15, -1.685454e-14, -5.639077e-15, -1.96688e-14, -8.74875e-15, 
    -1.207986e-14, -1.655243e-14, -1.244858e-14, -1.09932e-14, -9.840365e-15, 
    -1.689168e-14, -5.80261e-15, -1.739497e-14, -1.440284e-14, -1.427338e-14, 
    -8.77181e-15, -1.273943e-14, -1.5646e-14, -1.554895e-14, -7.847979e-15, 
    -1.176285e-14, -1.695744e-14, -7.024256e-16, -1.632961e-14, -1.14702e-14, 
    -7.164469e-15, -1.399706e-14, -8.343297e-15, -1.413539e-14, 
    -1.335789e-14, -9.016026e-15, -1.552982e-14, -1.1403e-14, -1.110526e-14, 
    -1.614274e-14, -7.961818e-15, -1.038804e-14, -1.494277e-14, 
    -8.678329e-15, -1.845092e-14, -1.54658e-14, -1.373531e-14, -8.373727e-15, 
    -2.30511e-14, -9.420744e-15, -1.635837e-14, -1.709434e-14, -2.244141e-14, 
    -1.44e-14, -1.299672e-14, -1.604615e-14, -1.143153e-14, -1.164588e-14, 
    -1.049017e-14, -1.203487e-14, -1.563069e-14, -1.518873e-14, 
    -1.352164e-14, -1.209272e-14, -9.012979e-15, -1.234928e-14, 
    -1.253892e-14, -1.420086e-14, -1.591435e-14, -1.566496e-14, 
    -9.423579e-15, -6.792402e-15, -8.072148e-15, -1.506171e-14, 
    -9.597033e-15, -1.204596e-14, -1.850462e-14, -6.180524e-15, 
    -1.267146e-14, -8.919134e-15, -1.933254e-14, -8.830816e-15, -1.51399e-14, 
    -1.34623e-14, -1.837181e-14, -1.243792e-14, -1.242513e-14, -2.045697e-14, 
    -1.000274e-14, -1.81999e-14, -1.086713e-14, -1.224568e-14, -1.022684e-14, 
    -1.752262e-14, -1.822031e-14, -9.553336e-15, -1.055409e-14, 
    -7.810791e-15, -1.438148e-14, -1.559365e-14, -1.700984e-14, -1.14453e-14, 
    -1.508718e-14, -1.438936e-14, -8.344583e-15, -1.072115e-14, 
    -1.444159e-14, -1.791237e-14, -1.505492e-14, -1.08931e-14, -1.457316e-14, 
    -1.486123e-14, -2.356738e-14, -4.027646e-15, -1.856453e-14, 
    -1.461754e-14, -1.991871e-14, -1.751098e-14, -1.277513e-14, 7.596263e-16, 
    -1.36055e-14, -1.375714e-14, -1.471978e-14, -8.01967e-15, -1.243213e-14, 
    -1.166638e-14, -1.22232e-14, -9.2486e-15, -1.377619e-14, -1.173762e-14, 
    -1.487328e-14, -1.481856e-14, -1.254566e-14, -4.339086e-15, 
    -8.307764e-15, -1.739225e-14, -1.358075e-14, -7.143966e-15, 
    -8.123886e-15, -2.040752e-14, -1.529945e-14, -1.37709e-14, -4.950842e-15, 
    -6.988017e-15, -1.19513e-14, -7.933475e-15, -2.135104e-14, -8.162951e-15, 
    -1.269508e-14, -1.916429e-14, -8.573668e-15, -1.728463e-14, -1.25932e-14, 
    -1.215914e-14, -1.599073e-14, -1.621218e-14, -6.553629e-15, 
    -1.587046e-14, -1.388182e-14, -1.153041e-14, -8.159237e-15, 
    -1.406266e-14, -1.658995e-14, -1.85469e-14, -1.118485e-14, -7.451176e-15, 
    -1.576737e-14, -1.5625e-14, -1.015265e-14, -1.303549e-14, -1.351418e-14, 
    -1.442166e-14, -1.035459e-14, -1.223443e-14, -1.156078e-14, -1.52318e-14, 
    -6.594184e-15, -1.284913e-14, -1.094856e-14, -1.383914e-14, 
    -1.726626e-14, -1.32938e-14, -1.561598e-14, -1.465295e-14, -9.352454e-15, 
    -1.760876e-14, -7.285926e-15, -1.202879e-14, -1.074784e-14, 
    -1.627313e-14, -8.036201e-15, -1.567813e-14, -1.345799e-14, 
    -1.087248e-14, -1.232543e-14, -1.024796e-14, -1.382399e-14, 
    -1.707666e-14, -9.060046e-15, -1.57753e-14, -1.536633e-14 ;

 ERRSOI =
  -3.4123e-10, -4.076417e-10, -4.755323e-10, -2.960974e-10, -3.576276e-10, 
    -3.840394e-10, -3.544538e-10, -1.188584e-10, -5.175866e-10, 
    -3.419213e-10, -3.963501e-10, -2.048557e-10, -4.608771e-10, -2.15177e-10, 
    -2.644217e-10, -2.293828e-10, -5.84996e-10, -1.957638e-10, -4.510394e-10, 
    -2.796608e-10, -3.041318e-10, -6.067933e-10, -1.683169e-10, 
    -3.361474e-10, -2.998922e-10, -3.982757e-10, -2.984606e-10, 
    -2.037765e-10, -3.738456e-10, -1.342628e-10, -1.569963e-10, 
    -2.327115e-10, -3.395266e-10, -5.473351e-10, -3.523465e-10, 
    -3.654134e-10, -3.791566e-10, -3.469084e-10, -3.506816e-10, 
    -3.204837e-10, -1.153566e-10, -1.409764e-10, -4.583232e-10, 
    -1.502647e-10, -2.533883e-10, -3.781498e-10, -2.456916e-10, 
    -4.297599e-10, -4.137463e-10, -5.096787e-10, -1.975519e-10, 
    -3.002295e-10, -3.181704e-10, -2.194954e-10, -1.507183e-10, 
    -2.377053e-10, -2.431126e-10, -3.348355e-11, -4.278954e-10, 
    -3.924745e-10, -1.663656e-10, -3.089359e-10, -2.225424e-10, 
    -3.463053e-10, -2.364165e-10, -2.620652e-10, -3.744322e-10, 
    -1.581697e-10, -3.375616e-10, -4.183007e-10, -3.354927e-10, 
    -2.341891e-10, -1.874846e-10, -4.157185e-10, -2.377144e-10, 
    -3.806817e-10, -3.62767e-10, -2.866717e-10, -2.062141e-10, -2.24318e-10, 
    -2.190118e-10, -2.812643e-10, -1.82988e-10, -3.213221e-10, -3.882221e-10, 
    -1.217018e-10, -3.668522e-10, -2.331218e-10, -4.208275e-10, 
    -1.129466e-10, -3.416843e-10, -2.464727e-10, -2.931841e-10, 
    -3.776812e-10, -4.982373e-11, -3.720114e-10, -3.23976e-10, -2.39775e-10, 
    -3.368873e-10, -2.994864e-10, -3.292467e-10, -2.436278e-10, 
    -3.585194e-10, -2.713791e-10, -2.659364e-10, -2.27185e-10, -4.387243e-10, 
    -1.036837e-10, -1.998666e-10, -1.333116e-10, -3.226048e-10, 
    -3.268787e-10, -2.909511e-10, -3.558779e-10, -1.95474e-10, -1.241162e-10, 
    -2.567317e-10, -2.744167e-10, -1.510723e-10, -3.710074e-10, 
    -2.150464e-10, -4.163451e-10, -3.503036e-10, -4.686824e-10, -5.0715e-10, 
    -3.407763e-10, -3.415822e-10, -3.04726e-10, -9.236691e-11, -3.020147e-10, 
    -2.335744e-11, -1.759231e-10, -2.650237e-10, -2.550631e-10, 
    -3.541462e-10, -3.229953e-10, -3.901028e-10, -2.877353e-10, 
    -3.430213e-10, -2.098476e-10, -1.949422e-10, -1.964785e-10, 
    -1.230237e-10, -1.488941e-10, -3.253005e-10, -5.056351e-10, 
    -2.321282e-10, -3.467535e-10, -4.108079e-10, -3.411657e-10, 
    -3.939886e-10, -2.936403e-10, -3.381014e-10, -1.798155e-10, -2.2539e-10, 
    -2.611746e-10, -4.278366e-10, -1.954794e-10, -1.662182e-10, 
    -3.188924e-10, -2.178966e-10, -3.26766e-10, -3.596194e-10, -2.523292e-10, 
    -3.99143e-10, -2.15491e-10, -2.479587e-10, -3.197033e-10, -2.011142e-10, 
    -4.193844e-10, -3.115712e-10, -1.912034e-10, -3.480848e-10, 
    -3.576597e-10, -2.608102e-10, -3.006188e-10, -4.134814e-10, 
    -2.763731e-10, -8.050539e-11, -4.104347e-10, -2.515745e-10, 
    -2.834615e-10, -2.575271e-10, -2.715115e-10, -2.206139e-10, 
    -4.564935e-10, -2.177934e-10, -1.890834e-10, -3.681742e-10, 
    -2.539482e-10, -2.368183e-10, -3.707912e-10, -1.747709e-10, 
    -3.278985e-10, -3.306138e-10, -2.071457e-10, -3.68895e-10, -4.678916e-10, 
    -7.03987e-11, -1.65193e-10, -2.242371e-10, -2.850104e-10, -4.607109e-10, 
    -3.377044e-10, -2.965344e-10, -2.616618e-10, 3.776629e-11, -2.751932e-10, 
    -2.56812e-10, -2.249154e-10, -3.525382e-10, -1.461216e-10, -1.221925e-10, 
    -1.826798e-10, -4.184328e-10, -1.475437e-10, -1.424878e-10, 
    -3.388989e-10, -1.210823e-10, -1.830505e-10, -2.53381e-10, -4.777888e-10, 
    -3.130119e-10, -1.483143e-10, -2.46615e-10, -1.139801e-10, -1.999283e-10, 
    -2.427038e-10, -2.047044e-10, -3.006662e-10, -3.808888e-10, 
    -4.394859e-10, -3.389861e-10, -3.731885e-10, -1.603574e-10, 
    -4.454178e-10, -2.716375e-10, -5.548202e-10, -3.202428e-10, 
    -3.383325e-11, -2.741923e-10, -4.505622e-10, -4.429324e-10, 
    -2.683238e-10, -4.72741e-10, -4.494027e-10, -3.110102e-10, -3.914225e-10, 
    -2.347426e-10, -1.775878e-10, -2.329805e-10, -2.949769e-10, 
    -2.743707e-10, -2.062315e-10, -4.247224e-10, -3.676296e-10, 
    -3.163731e-10, -1.938576e-10, -3.666382e-10, -3.974516e-10, 
    -1.608962e-10, -3.464289e-10, -4.95552e-10, -2.23686e-10, -1.956021e-10, 
    -2.289153e-10, -2.812572e-10, -3.010655e-10, -2.704527e-10, 
    -2.354366e-10, -4.357321e-10, -4.462044e-10, -1.781727e-10, -1.92792e-10, 
    -1.982855e-10, -4.932645e-10, -2.673648e-10, -6.486505e-11, 
    -3.052736e-10, -3.383263e-10, -2.859513e-10, -4.573296e-10, 
    -3.164858e-10, -3.003424e-10, -3.149373e-10, -2.29505e-10, -2.542437e-10, 
    -3.700196e-10, -3.874606e-10, -2.23054e-10, -1.438262e-10, -1.711525e-10, 
    -5.308117e-10, -3.266881e-10, -5.51153e-10, -2.116898e-10, -2.912782e-10, 
    -3.212373e-10, -3.774093e-10, -2.26027e-10, -4.491376e-10, -2.32757e-10, 
    -2.672713e-10, -4.450538e-10, -2.812452e-10, -2.564129e-10, 
    -4.006419e-10, -3.268354e-10, -3.694379e-10, -3.950484e-10, 
    -3.417375e-10, -2.733884e-10, -4.150711e-10, -2.877947e-10, 
    -2.410909e-10, -2.13893e-10, -2.282598e-10, -3.34989e-10, -2.992751e-10, 
    -3.42883e-10, -3.241379e-10, -3.216006e-10, -3.19163e-10, -2.300111e-10, 
    -2.406084e-10, -1.271493e-10, -2.294818e-10, -6.831901e-11, 
    -4.278676e-10, -3.164463e-10, -3.56646e-10, -8.995685e-11, -4.438751e-10, 
    -1.449762e-10, -2.493135e-10, -4.053142e-10, -4.463571e-10, -2.46636e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  5.789056e-16, 5.727179e-16, 5.739225e-16, 5.689207e-16, 5.716972e-16, 
    5.684196e-16, 5.77653e-16, 5.724715e-16, 5.75781e-16, 5.783499e-16, 
    5.591791e-16, 5.686974e-16, 5.492518e-16, 5.553543e-16, 5.39994e-16, 
    5.502021e-16, 5.379303e-16, 5.402902e-16, 5.331827e-16, 5.352212e-16, 
    5.261039e-16, 5.322413e-16, 5.213654e-16, 5.275717e-16, 5.266014e-16, 
    5.324433e-16, 5.667863e-16, 5.603661e-16, 5.671659e-16, 5.662518e-16, 
    5.666622e-16, 5.716395e-16, 5.741426e-16, 5.793785e-16, 5.784291e-16, 
    5.745834e-16, 5.658406e-16, 5.688131e-16, 5.613157e-16, 5.614853e-16, 
    5.531077e-16, 5.56889e-16, 5.427608e-16, 5.467857e-16, 5.351362e-16, 
    5.380714e-16, 5.352739e-16, 5.361227e-16, 5.352629e-16, 5.395662e-16, 
    5.377234e-16, 5.415068e-16, 5.561811e-16, 5.518782e-16, 5.646859e-16, 
    5.723488e-16, 5.774259e-16, 5.810203e-16, 5.805125e-16, 5.79544e-16, 
    5.745609e-16, 5.698658e-16, 5.662805e-16, 5.638787e-16, 5.615097e-16, 
    5.543203e-16, 5.505078e-16, 5.419455e-16, 5.434941e-16, 5.408708e-16, 
    5.383632e-16, 5.341457e-16, 5.348405e-16, 5.329803e-16, 5.409408e-16, 
    5.35653e-16, 5.443754e-16, 5.41993e-16, 5.608616e-16, 5.680118e-16, 
    5.710406e-16, 5.736909e-16, 5.80122e-16, 5.756827e-16, 5.774337e-16, 
    5.732662e-16, 5.706133e-16, 5.71926e-16, 5.638129e-16, 5.669707e-16, 
    5.502816e-16, 5.574859e-16, 5.386558e-16, 5.431764e-16, 5.375711e-16, 
    5.404333e-16, 5.355266e-16, 5.399431e-16, 5.322879e-16, 5.306172e-16, 
    5.317589e-16, 5.273712e-16, 5.401875e-16, 5.352736e-16, 5.719626e-16, 
    5.717485e-16, 5.707514e-16, 5.751308e-16, 5.753985e-16, 5.794043e-16, 
    5.758407e-16, 5.74321e-16, 5.704597e-16, 5.681718e-16, 5.659949e-16, 
    5.612006e-16, 5.558331e-16, 5.483063e-16, 5.428836e-16, 5.392412e-16, 
    5.414756e-16, 5.39503e-16, 5.417079e-16, 5.427407e-16, 5.312431e-16, 
    5.37706e-16, 5.280028e-16, 5.285409e-16, 5.329359e-16, 5.284803e-16, 
    5.715983e-16, 5.728297e-16, 5.770984e-16, 5.737585e-16, 5.798401e-16, 
    5.764376e-16, 5.744785e-16, 5.66904e-16, 5.65237e-16, 5.636889e-16, 
    5.606291e-16, 5.566956e-16, 5.497776e-16, 5.437414e-16, 5.382174e-16, 
    5.386227e-16, 5.3848e-16, 5.372439e-16, 5.403041e-16, 5.367411e-16, 
    5.361423e-16, 5.377072e-16, 5.286129e-16, 5.312148e-16, 5.285523e-16, 
    5.302469e-16, 5.724296e-16, 5.703569e-16, 5.714771e-16, 5.6937e-16, 
    5.708544e-16, 5.642448e-16, 5.622591e-16, 5.529444e-16, 5.567729e-16, 
    5.506776e-16, 5.561548e-16, 5.55185e-16, 5.50477e-16, 5.558594e-16, 
    5.44074e-16, 5.520697e-16, 5.371958e-16, 5.452033e-16, 5.36693e-16, 
    5.382413e-16, 5.356776e-16, 5.333786e-16, 5.304838e-16, 5.251319e-16, 
    5.263725e-16, 5.218904e-16, 5.672636e-16, 5.64568e-16, 5.648061e-16, 
    5.619822e-16, 5.598913e-16, 5.553532e-16, 5.480542e-16, 5.508021e-16, 
    5.457556e-16, 5.447409e-16, 5.52407e-16, 5.477026e-16, 5.627624e-16, 
    5.603357e-16, 5.617814e-16, 5.670507e-16, 5.501682e-16, 5.588484e-16, 
    5.427937e-16, 5.475161e-16, 5.337065e-16, 5.405841e-16, 5.27055e-16, 
    5.212454e-16, 5.15768e-16, 5.093474e-16, 5.63096e-16, 5.649293e-16, 
    5.616463e-16, 5.570948e-16, 5.528652e-16, 5.472282e-16, 5.46651e-16, 
    5.45593e-16, 5.428508e-16, 5.405422e-16, 5.452577e-16, 5.399632e-16, 
    5.597711e-16, 5.494134e-16, 5.656213e-16, 5.607525e-16, 5.573637e-16, 
    5.588516e-16, 5.511161e-16, 5.492885e-16, 5.418469e-16, 5.456973e-16, 
    5.2268e-16, 5.328918e-16, 5.044496e-16, 5.124314e-16, 5.655692e-16, 
    5.631026e-16, 5.544953e-16, 5.585951e-16, 5.468518e-16, 5.439513e-16, 
    5.415913e-16, 5.385697e-16, 5.382438e-16, 5.364514e-16, 5.393877e-16, 
    5.365677e-16, 5.472162e-16, 5.424639e-16, 5.554817e-16, 5.5232e-16, 
    5.537753e-16, 5.5537e-16, 5.504444e-16, 5.451833e-16, 5.450719e-16, 
    5.43382e-16, 5.386114e-16, 5.468041e-16, 5.213567e-16, 5.371038e-16, 
    5.604098e-16, 5.556435e-16, 5.549632e-16, 5.568111e-16, 5.442422e-16, 
    5.488045e-16, 5.364953e-16, 5.398289e-16, 5.343646e-16, 5.370814e-16, 
    5.374808e-16, 5.409651e-16, 5.431314e-16, 5.485953e-16, 5.530315e-16, 
    5.565433e-16, 5.557273e-16, 5.518679e-16, 5.448614e-16, 5.382137e-16, 
    5.396714e-16, 5.347803e-16, 5.477053e-16, 5.422941e-16, 5.443867e-16, 
    5.389263e-16, 5.508748e-16, 5.407007e-16, 5.534675e-16, 5.523513e-16, 
    5.488949e-16, 5.419258e-16, 5.403827e-16, 5.387319e-16, 5.397509e-16, 
    5.446834e-16, 5.45491e-16, 5.489793e-16, 5.49941e-16, 5.525944e-16, 
    5.547884e-16, 5.527837e-16, 5.506762e-16, 5.446818e-16, 5.392654e-16, 
    5.333457e-16, 5.318951e-16, 5.249522e-16, 5.306041e-16, 5.212685e-16, 
    5.292055e-16, 5.154503e-16, 5.401113e-16, 5.294408e-16, 5.487379e-16, 
    5.466672e-16, 5.429157e-16, 5.342902e-16, 5.38952e-16, 5.334997e-16, 
    5.455227e-16, 5.51734e-16, 5.533396e-16, 5.563298e-16, 5.532712e-16, 
    5.535201e-16, 5.505897e-16, 5.515319e-16, 5.444825e-16, 5.482719e-16, 
    5.374905e-16, 5.33543e-16, 5.223601e-16, 5.154776e-16, 5.084532e-16, 
    5.053452e-16, 5.043984e-16, 5.040025e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGR =
  -383.7672, -384.821, -384.6164, -385.4658, -384.9948, -385.5508, -383.9812, 
    -384.8626, -384.3001, -383.8625, -387.1216, -385.5038, -388.8035, 
    -387.7688, -390.355, -388.6348, -390.7001, -390.3063, -391.4929, 
    -391.153, -392.6688, -391.6497, -393.4552, -392.4258, -392.5866, 
    -391.616, -385.8282, -386.9211, -385.7639, -385.9185, -385.8492, 
    -385.0044, -384.5781, -383.6871, -383.849, -384.5036, -385.9881, 
    -385.4846, -386.7631, -386.7345, -388.1472, -387.5103, -389.8929, 
    -389.2185, -391.1672, -390.6772, -391.1441, -391.0026, -391.1459, 
    -390.4272, -390.7351, -390.1029, -387.6295, -388.3539, -386.1839, 
    -384.8827, -384.0197, -383.4067, -383.4934, -383.6585, -384.5074, 
    -385.306, -385.9142, -386.3296, -386.7303, -387.9416, -388.5838, 
    -390.0289, -389.7703, -390.2088, -390.6284, -391.3321, -391.2164, 
    -391.5262, -390.1976, -391.0805, -389.6228, -390.0215, -386.8372, 
    -385.6206, -385.1052, -384.6556, -383.56, -384.3165, -384.0182, 
    -384.7282, -385.179, -384.9562, -386.3407, -385.7971, -388.6218, 
    -387.4092, -390.5795, -389.8234, -390.7608, -390.2826, -391.1017, 
    -390.3645, -391.6417, -391.9195, -391.7296, -392.4596, -390.3236, 
    -391.1439, -384.9498, -384.9861, -385.1556, -384.4105, -384.365, 
    -383.6825, -384.29, -384.5484, -385.2053, -385.5934, -385.9624, 
    -386.7823, -387.6878, -388.9627, -389.8724, -390.4819, -390.1083, 
    -390.4381, -390.0693, -389.8966, -391.8153, -390.7379, -392.3546, 
    -392.2653, -391.5335, -392.2754, -385.0117, -384.8026, -384.0756, 
    -384.6445, -383.6082, -384.1881, -384.5213, -385.8078, -386.0909, 
    -386.3615, -386.879, -387.5429, -388.7157, -389.7284, -390.653, 
    -390.5853, -390.6091, -390.8153, -390.3041, -390.8993, -390.999, 
    -390.738, -392.2533, -391.8205, -392.2634, -391.9817, -384.8706, 
    -385.2226, -385.0323, -385.39, -385.1379, -386.2668, -386.6026, -388.174, 
    -387.5297, -388.5556, -387.6341, -387.7973, -388.5882, -387.6841, 
    -389.6722, -388.3209, -390.8234, -389.4824, -390.9073, -390.649, 
    -391.0769, -391.46, -391.9421, -392.8309, -392.6252, -393.3687, 
    -385.7475, -386.2038, -386.164, -386.6503, -387.0035, -387.7693, 
    -389.0054, -388.5353, -389.3914, -389.5613, -388.2655, -389.0641, 
    -386.518, -386.9277, -386.6841, -385.7833, -388.6411, -387.179, 
    -389.8873, -389.0958, -391.4053, -390.2566, -392.5119, -393.4744, 
    -394.3817, -395.4394, -386.4618, -386.1431, -386.7072, -387.4749, 
    -388.1881, -389.144, -389.2411, -389.4184, -389.8781, -390.2643, 
    -389.4741, -390.3612, -387.022, -388.7769, -386.0255, -386.8572, 
    -387.4298, -387.179, -388.4826, -388.7984, -390.0455, -389.4012, 
    -393.2365, -391.5403, -396.2457, -394.9315, -386.0347, -386.4609, 
    -387.9133, -387.2224, -389.2075, -389.6935, -390.089, -390.5937, 
    -390.6485, -390.9475, -390.4574, -390.9283, -389.146, -389.9427, 
    -387.7478, -388.2798, -388.0352, -387.7666, -388.5955, -389.4865, 
    -389.5059, -389.7886, -390.584, -389.2155, -393.4542, -390.8362, 
    -386.9162, -387.7194, -387.8349, -387.5237, -389.6448, -388.8795, 
    -390.9403, -390.3836, -391.2958, -390.8425, -390.7758, -390.1936, 
    -389.8309, -388.9145, -388.16, -387.5689, -387.7064, -388.3557, 
    -389.5406, -390.6531, -390.4094, -391.2265, -389.0642, -389.9708, 
    -389.6202, -390.5343, -388.5229, -390.2352, -388.087, -388.2748, 
    -388.8643, -390.0318, -390.291, -390.5666, -390.3967, -389.5705, 
    -389.4354, -388.8503, -388.6797, -388.234, -387.8646, -388.2019, 
    -388.556, -389.5711, -390.4774, -391.4653, -391.7073, -392.8594, 
    -391.9207, -393.4686, -392.1514, -394.4318, -390.3349, -392.1139, 
    -388.8909, -389.2385, -389.8663, -391.3071, -390.5301, -391.4391, 
    -389.4302, -388.3778, -388.1085, -387.6047, -388.12, -388.0782, 
    -388.5711, -388.4128, -389.6046, -388.9691, -390.774, -391.4321, 
    -393.2906, -394.4287, -395.5877, -396.0989, -396.2545, -396.3195 ;

 FGR12 =
  -49.04824, -49.12321, -49.10867, -49.16917, -49.13564, -49.17525, 
    -49.06347, -49.12615, -49.08615, -49.05504, -49.28682, -49.17192, 
    -49.40692, -49.33339, -49.51856, -49.39547, -49.54348, -49.51513, 
    -49.6008, -49.57624, -49.68585, -49.61216, -49.74296, -49.6683, 
    -49.67991, -49.60971, -49.1951, -49.27247, -49.19049, -49.20152, 
    -49.19658, -49.13629, -49.10587, -49.04258, -49.05408, -49.10061, 
    -49.20647, -49.17057, -49.26134, -49.2593, -49.36053, -49.31487, 
    -49.48533, -49.43683, -49.57726, -49.54188, -49.57559, -49.56538, 
    -49.57571, -49.52385, -49.54605, -49.50047, -49.32339, -49.37532, 
    -49.22048, -49.12756, -49.0662, -49.02266, -49.0288, -49.04052, 
    -49.10089, -49.15781, -49.20124, -49.23031, -49.25901, -49.34568, 
    -49.39182, -49.49509, -49.47652, -49.50807, -49.53837, -49.58915, 
    -49.58082, -49.60319, -49.50731, -49.57096, -49.46592, -49.4946, 
    -49.26646, -49.18027, -49.14341, -49.11145, -49.03354, -49.08729, 
    -49.06609, -49.11663, -49.14876, -49.13289, -49.23111, -49.19288, 
    -49.39452, -49.30759, -49.53481, -49.48034, -49.5479, -49.51344, 
    -49.57251, -49.51934, -49.61155, -49.63163, -49.61791, -49.67076, 
    -49.51639, -49.57555, -49.13243, -49.13501, -49.14709, -49.09398, 
    -49.09074, -49.04225, -49.08543, -49.10381, -49.15065, -49.17833, 
    -49.20469, -49.26269, -49.32756, -49.41838, -49.48386, -49.52779, 
    -49.50088, -49.52464, -49.49806, -49.48563, -49.62408, -49.54625, 
    -49.66316, -49.6567, -49.60373, -49.65742, -49.13683, -49.12194, 
    -49.07018, -49.11068, -49.03698, -49.07816, -49.10187, -49.19359, 
    -49.21388, -49.23258, -49.26963, -49.31719, -49.40067, -49.47346, 
    -49.54014, -49.53525, -49.53698, -49.55185, -49.51498, -49.5579, 
    -49.56509, -49.54627, -49.65582, -49.6245, -49.65656, -49.63617, 
    -49.12679, -49.15187, -49.13831, -49.1638, -49.14583, -49.22576, 
    -49.24979, -49.36239, -49.31625, -49.3898, -49.32374, -49.33543, 
    -49.39206, -49.32734, -49.46938, -49.37293, -49.55241, -49.45571, 
    -49.55848, -49.53985, -49.57075, -49.5984, -49.6333, -49.69765, 
    -49.68277, -49.73671, -49.18934, -49.2219, -49.21909, -49.25325, 
    -49.27853, -49.33344, -49.42147, -49.3884, -49.44925, -49.46146, 
    -49.36904, -49.42569, -49.24378, -49.27306, -49.25566, -49.19188, 
    -49.39592, -49.29108, -49.48493, -49.428, -49.59444, -49.51152, 
    -49.67456, -49.74431, -49.81041, -49.88744, -49.23976, -49.21761, 
    -49.25735, -49.31227, -49.36347, -49.43144, -49.43845, -49.45119, 
    -49.48429, -49.51211, -49.45517, -49.51908, -49.27975, -49.40503, 
    -49.20919, -49.26799, -49.30906, -49.2911, -49.38462, -49.40664, 
    -49.49631, -49.44997, -49.72702, -49.60418, -49.94641, -49.85041, 
    -49.20986, -49.23972, -49.34374, -49.29422, -49.43603, -49.47098, 
    -49.49948, -49.53584, -49.53981, -49.56138, -49.52604, -49.56, -49.4316, 
    -49.48892, -49.33191, -49.37004, -49.35252, -49.33326, -49.39273, 
    -49.45603, -49.4575, -49.47781, -49.53495, -49.43663, -49.74271, 
    -49.55322, -49.27231, -49.32979, -49.33814, -49.31583, -49.46747, 
    -49.41245, -49.56086, -49.52072, -49.58655, -49.55382, -49.54899, 
    -49.50702, -49.48087, -49.41496, -49.36145, -49.31908, -49.32895, 
    -49.37548, -49.45995, -49.54011, -49.52254, -49.58154, -49.42575, 
    -49.49093, -49.4657, -49.53157, -49.38751, -49.50982, -49.35625, 
    -49.36971, -49.41137, -49.49527, -49.51404, -49.53387, -49.52164, 
    -49.46212, -49.4524, -49.41037, -49.39874, -49.36679, -49.3403, 
    -49.36447, -49.38986, -49.46217, -49.52745, -49.59877, -49.61632, 
    -49.69962, -49.63166, -49.74376, -49.64825, -49.81389, -49.51711, 
    -49.64559, -49.4133, -49.43826, -49.48339, -49.58728, -49.53127, 
    -49.59684, -49.45203, -49.37705, -49.35778, -49.32164, -49.3586, 
    -49.35561, -49.39097, -49.37961, -49.46458, -49.41891, -49.54885, 
    -49.59636, -49.73103, -49.81376, -49.89835, -49.93571, -49.94709, 
    -49.95186 ;

 FGR_R =
  -383.7672, -384.821, -384.6164, -385.4658, -384.9948, -385.5508, -383.9812, 
    -384.8626, -384.3001, -383.8625, -387.1216, -385.5038, -388.8035, 
    -387.7688, -390.355, -388.6348, -390.7001, -390.3063, -391.4929, 
    -391.153, -392.6688, -391.6497, -393.4552, -392.4258, -392.5866, 
    -391.616, -385.8282, -386.9211, -385.7639, -385.9185, -385.8492, 
    -385.0044, -384.5781, -383.6871, -383.849, -384.5036, -385.9881, 
    -385.4846, -386.7631, -386.7345, -388.1472, -387.5103, -389.8929, 
    -389.2185, -391.1672, -390.6772, -391.1441, -391.0026, -391.1459, 
    -390.4272, -390.7351, -390.1029, -387.6295, -388.3539, -386.1839, 
    -384.8827, -384.0197, -383.4067, -383.4934, -383.6585, -384.5074, 
    -385.306, -385.9142, -386.3296, -386.7303, -387.9416, -388.5838, 
    -390.0289, -389.7703, -390.2088, -390.6284, -391.3321, -391.2164, 
    -391.5262, -390.1976, -391.0805, -389.6228, -390.0215, -386.8372, 
    -385.6206, -385.1052, -384.6556, -383.56, -384.3165, -384.0182, 
    -384.7282, -385.179, -384.9562, -386.3407, -385.7971, -388.6218, 
    -387.4092, -390.5795, -389.8234, -390.7608, -390.2826, -391.1017, 
    -390.3645, -391.6417, -391.9195, -391.7296, -392.4596, -390.3236, 
    -391.1439, -384.9498, -384.9861, -385.1556, -384.4105, -384.365, 
    -383.6825, -384.29, -384.5484, -385.2053, -385.5934, -385.9624, 
    -386.7823, -387.6878, -388.9627, -389.8724, -390.4819, -390.1083, 
    -390.4381, -390.0693, -389.8966, -391.8153, -390.7379, -392.3546, 
    -392.2653, -391.5335, -392.2754, -385.0117, -384.8026, -384.0756, 
    -384.6445, -383.6082, -384.1881, -384.5213, -385.8078, -386.0909, 
    -386.3615, -386.879, -387.5429, -388.7157, -389.7284, -390.653, 
    -390.5853, -390.6091, -390.8153, -390.3041, -390.8993, -390.999, 
    -390.738, -392.2533, -391.8205, -392.2634, -391.9817, -384.8706, 
    -385.2226, -385.0323, -385.39, -385.1379, -386.2668, -386.6026, -388.174, 
    -387.5297, -388.5556, -387.6341, -387.7973, -388.5882, -387.6841, 
    -389.6722, -388.3209, -390.8234, -389.4824, -390.9073, -390.649, 
    -391.0769, -391.46, -391.9421, -392.8309, -392.6252, -393.3687, 
    -385.7475, -386.2038, -386.164, -386.6503, -387.0035, -387.7693, 
    -389.0054, -388.5353, -389.3914, -389.5613, -388.2655, -389.0641, 
    -386.518, -386.9277, -386.6841, -385.7833, -388.6411, -387.179, 
    -389.8873, -389.0958, -391.4053, -390.2566, -392.5119, -393.4744, 
    -394.3817, -395.4394, -386.4618, -386.1431, -386.7072, -387.4749, 
    -388.1881, -389.144, -389.2411, -389.4184, -389.8781, -390.2643, 
    -389.4741, -390.3612, -387.022, -388.7769, -386.0255, -386.8572, 
    -387.4298, -387.179, -388.4826, -388.7984, -390.0455, -389.4012, 
    -393.2365, -391.5403, -396.2457, -394.9315, -386.0347, -386.4609, 
    -387.9133, -387.2224, -389.2075, -389.6935, -390.089, -390.5937, 
    -390.6485, -390.9475, -390.4574, -390.9283, -389.146, -389.9427, 
    -387.7478, -388.2798, -388.0352, -387.7666, -388.5955, -389.4865, 
    -389.5059, -389.7886, -390.584, -389.2155, -393.4542, -390.8362, 
    -386.9162, -387.7194, -387.8349, -387.5237, -389.6448, -388.8795, 
    -390.9403, -390.3836, -391.2958, -390.8425, -390.7758, -390.1936, 
    -389.8309, -388.9145, -388.16, -387.5689, -387.7064, -388.3557, 
    -389.5406, -390.6531, -390.4094, -391.2265, -389.0642, -389.9708, 
    -389.6202, -390.5343, -388.5229, -390.2352, -388.087, -388.2748, 
    -388.8643, -390.0318, -390.291, -390.5666, -390.3967, -389.5705, 
    -389.4354, -388.8503, -388.6797, -388.234, -387.8646, -388.2019, 
    -388.556, -389.5711, -390.4774, -391.4653, -391.7073, -392.8594, 
    -391.9207, -393.4686, -392.1514, -394.4318, -390.3349, -392.1139, 
    -388.8909, -389.2385, -389.8663, -391.3071, -390.5301, -391.4391, 
    -389.4302, -388.3778, -388.1085, -387.6047, -388.12, -388.0782, 
    -388.5711, -388.4128, -389.6046, -388.9691, -390.774, -391.4321, 
    -393.2906, -394.4287, -395.5877, -396.0989, -396.2545, -396.3195 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  47.7017, 47.77869, 47.76374, 47.82581, 47.7914, 47.83202, 47.71733, 
    47.78173, 47.74063, 47.70866, 47.94583, 47.82858, 48.06783, 47.99315, 
    48.18122, 48.05642, 48.20644, 48.17767, 48.26439, 48.23956, 48.35033, 
    48.27586, 48.40782, 48.33258, 48.34433, 48.27339, 47.8523, 47.93118, 
    47.84759, 47.85889, 47.85383, 47.79209, 47.76094, 47.69585, 47.70768, 
    47.7555, 47.86397, 47.82719, 47.91967, 47.91758, 48.0208, 47.97426, 
    48.14745, 48.09818, 48.24059, 48.20478, 48.2389, 48.22856, 48.23904, 
    48.18651, 48.20901, 48.1628, 47.98297, 48.0359, 47.87828, 47.78319, 
    47.72015, 47.67537, 47.6817, 47.69376, 47.75578, 47.81413, 47.85858, 
    47.88799, 47.91727, 48.00576, 48.0527, 48.15739, 48.13849, 48.17054, 
    48.20121, 48.25264, 48.24419, 48.26683, 48.16973, 48.23425, 48.12772, 
    48.15686, 47.92505, 47.83712, 47.79945, 47.76661, 47.68656, 47.74183, 
    47.72004, 47.77192, 47.80486, 47.78857, 47.8888, 47.85003, 48.05548, 
    47.96687, 48.19764, 48.14238, 48.21089, 48.17594, 48.2358, 48.18193, 
    48.27527, 48.29557, 48.2817, 48.33506, 48.17894, 48.23888, 47.78811, 
    47.79076, 47.80315, 47.7487, 47.74537, 47.69551, 47.73989, 47.75878, 
    47.80678, 47.83514, 47.8621, 47.92107, 47.98722, 48.07947, 48.14596, 
    48.1905, 48.1632, 48.18731, 48.16035, 48.14773, 48.28795, 48.20921, 
    48.32738, 48.32085, 48.26736, 48.32159, 47.79263, 47.77735, 47.72424, 
    47.7658, 47.69009, 47.73245, 47.75679, 47.8508, 47.87149, 47.89031, 
    47.92813, 47.97664, 48.06142, 48.13543, 48.20301, 48.19806, 48.1998, 
    48.21487, 48.17751, 48.22101, 48.22829, 48.20922, 48.31998, 48.28834, 
    48.32071, 48.30012, 47.78232, 47.80804, 47.79414, 47.82027, 47.80185, 
    47.88339, 47.90792, 48.02275, 47.97568, 48.05064, 47.98331, 47.99523, 
    48.05301, 47.98696, 48.13132, 48.03348, 48.21546, 48.11744, 48.2216, 
    48.20271, 48.23399, 48.26199, 48.29723, 48.36219, 48.34716, 48.4015, 
    47.8464, 47.87973, 47.87683, 47.91142, 47.93723, 47.99319, 48.08259, 
    48.04917, 48.1108, 48.12322, 48.02945, 48.08688, 47.90175, 47.93168, 
    47.91389, 47.84901, 48.05688, 47.95004, 48.14705, 48.0892, 48.25799, 
    48.17403, 48.33887, 48.40921, 48.47555, 48.55286, 47.89765, 47.87531, 
    47.91558, 47.97167, 48.02379, 48.09272, 48.09983, 48.11278, 48.14638, 
    48.1746, 48.11684, 48.18168, 47.93856, 48.06589, 47.86671, 47.92653, 
    47.96838, 47.95005, 48.04532, 48.06747, 48.15861, 48.11152, 48.39182, 
    48.26785, 48.61182, 48.51573, 47.86739, 47.89759, 48.00371, 47.95322, 
    48.09736, 48.13288, 48.16179, 48.19867, 48.20268, 48.22453, 48.18871, 
    48.22313, 48.09287, 48.1511, 47.99162, 48.03049, 48.01262, 47.99299, 
    48.05357, 48.11774, 48.11918, 48.13983, 48.19793, 48.09795, 48.40771, 
    48.21637, 47.93085, 47.98953, 47.99798, 47.97524, 48.12932, 48.07339, 
    48.22401, 48.18332, 48.24999, 48.21686, 48.21198, 48.16943, 48.14293, 
    48.07595, 48.02174, 47.97855, 47.98859, 48.03604, 48.1217, 48.20301, 
    48.1852, 48.24493, 48.08689, 48.15314, 48.12752, 48.19434, 48.04826, 
    48.17245, 48.01641, 48.03013, 48.07228, 48.1576, 48.17656, 48.19669, 
    48.18428, 48.12389, 48.11402, 48.07127, 48.05972, 48.02715, 48.00016, 
    48.02481, 48.05068, 48.12394, 48.19017, 48.26237, 48.28006, 48.36425, 
    48.29565, 48.40877, 48.31248, 48.47919, 48.17974, 48.30976, 48.07423, 
    48.09963, 48.14551, 48.2508, 48.19402, 48.26046, 48.11364, 48.03765, 
    48.01798, 47.98116, 48.01882, 48.01576, 48.05179, 48.04021, 48.12638, 
    48.07995, 48.21185, 48.25994, 48.39579, 48.47898, 48.56372, 48.60109, 
    48.61246, 48.61722 ;

 FIRA_R =
  47.7017, 47.77869, 47.76374, 47.82581, 47.7914, 47.83202, 47.71733, 
    47.78173, 47.74063, 47.70866, 47.94583, 47.82858, 48.06783, 47.99315, 
    48.18122, 48.05642, 48.20644, 48.17767, 48.26439, 48.23956, 48.35033, 
    48.27586, 48.40782, 48.33258, 48.34433, 48.27339, 47.8523, 47.93118, 
    47.84759, 47.85889, 47.85383, 47.79209, 47.76094, 47.69585, 47.70768, 
    47.7555, 47.86397, 47.82719, 47.91967, 47.91758, 48.0208, 47.97426, 
    48.14745, 48.09818, 48.24059, 48.20478, 48.2389, 48.22856, 48.23904, 
    48.18651, 48.20901, 48.1628, 47.98297, 48.0359, 47.87828, 47.78319, 
    47.72015, 47.67537, 47.6817, 47.69376, 47.75578, 47.81413, 47.85858, 
    47.88799, 47.91727, 48.00576, 48.0527, 48.15739, 48.13849, 48.17054, 
    48.20121, 48.25264, 48.24419, 48.26683, 48.16973, 48.23425, 48.12772, 
    48.15686, 47.92505, 47.83712, 47.79945, 47.76661, 47.68656, 47.74183, 
    47.72004, 47.77192, 47.80486, 47.78857, 47.8888, 47.85003, 48.05548, 
    47.96687, 48.19764, 48.14238, 48.21089, 48.17594, 48.2358, 48.18193, 
    48.27527, 48.29557, 48.2817, 48.33506, 48.17894, 48.23888, 47.78811, 
    47.79076, 47.80315, 47.7487, 47.74537, 47.69551, 47.73989, 47.75878, 
    47.80678, 47.83514, 47.8621, 47.92107, 47.98722, 48.07947, 48.14596, 
    48.1905, 48.1632, 48.18731, 48.16035, 48.14773, 48.28795, 48.20921, 
    48.32738, 48.32085, 48.26736, 48.32159, 47.79263, 47.77735, 47.72424, 
    47.7658, 47.69009, 47.73245, 47.75679, 47.8508, 47.87149, 47.89031, 
    47.92813, 47.97664, 48.06142, 48.13543, 48.20301, 48.19806, 48.1998, 
    48.21487, 48.17751, 48.22101, 48.22829, 48.20922, 48.31998, 48.28834, 
    48.32071, 48.30012, 47.78232, 47.80804, 47.79414, 47.82027, 47.80185, 
    47.88339, 47.90792, 48.02275, 47.97568, 48.05064, 47.98331, 47.99523, 
    48.05301, 47.98696, 48.13132, 48.03348, 48.21546, 48.11744, 48.2216, 
    48.20271, 48.23399, 48.26199, 48.29723, 48.36219, 48.34716, 48.4015, 
    47.8464, 47.87973, 47.87683, 47.91142, 47.93723, 47.99319, 48.08259, 
    48.04917, 48.1108, 48.12322, 48.02945, 48.08688, 47.90175, 47.93168, 
    47.91389, 47.84901, 48.05688, 47.95004, 48.14705, 48.0892, 48.25799, 
    48.17403, 48.33887, 48.40921, 48.47555, 48.55286, 47.89765, 47.87531, 
    47.91558, 47.97167, 48.02379, 48.09272, 48.09983, 48.11278, 48.14638, 
    48.1746, 48.11684, 48.18168, 47.93856, 48.06589, 47.86671, 47.92653, 
    47.96838, 47.95005, 48.04532, 48.06747, 48.15861, 48.11152, 48.39182, 
    48.26785, 48.61182, 48.51573, 47.86739, 47.89759, 48.00371, 47.95322, 
    48.09736, 48.13288, 48.16179, 48.19867, 48.20268, 48.22453, 48.18871, 
    48.22313, 48.09287, 48.1511, 47.99162, 48.03049, 48.01262, 47.99299, 
    48.05357, 48.11774, 48.11918, 48.13983, 48.19793, 48.09795, 48.40771, 
    48.21637, 47.93085, 47.98953, 47.99798, 47.97524, 48.12932, 48.07339, 
    48.22401, 48.18332, 48.24999, 48.21686, 48.21198, 48.16943, 48.14293, 
    48.07595, 48.02174, 47.97855, 47.98859, 48.03604, 48.1217, 48.20301, 
    48.1852, 48.24493, 48.08689, 48.15314, 48.12752, 48.19434, 48.04826, 
    48.17245, 48.01641, 48.03013, 48.07228, 48.1576, 48.17656, 48.19669, 
    48.18428, 48.12389, 48.11402, 48.07127, 48.05972, 48.02715, 48.00016, 
    48.02481, 48.05068, 48.12394, 48.19017, 48.26237, 48.28006, 48.36425, 
    48.29565, 48.40877, 48.31248, 48.47919, 48.17974, 48.30976, 48.07423, 
    48.09963, 48.14551, 48.2508, 48.19402, 48.26046, 48.11364, 48.03765, 
    48.01798, 47.98116, 48.01882, 48.01576, 48.05179, 48.04021, 48.12638, 
    48.07995, 48.21185, 48.25994, 48.39579, 48.47898, 48.56372, 48.60109, 
    48.61246, 48.61722 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  262.0479, 262.1248, 262.1099, 262.1719, 262.1375, 262.1782, 262.0635, 
    262.1279, 262.0868, 262.0548, 262.292, 262.1747, 262.414, 262.3393, 
    262.5274, 262.4026, 262.5526, 262.5238, 262.6105, 262.5857, 262.6965, 
    262.622, 262.754, 262.6787, 262.6905, 262.6195, 262.1985, 262.2773, 
    262.1937, 262.205, 262.2, 262.1382, 262.1071, 262.042, 262.0538, 
    262.1017, 262.2101, 262.1733, 262.2658, 262.2637, 262.3669, 262.3204, 
    262.4936, 262.4443, 262.5867, 262.5509, 262.5851, 262.5747, 262.5852, 
    262.5327, 262.5551, 262.5089, 262.3291, 262.382, 262.2244, 262.1293, 
    262.0663, 262.0215, 262.0278, 262.0399, 262.1019, 262.1603, 262.2047, 
    262.2341, 262.2634, 262.3519, 262.3988, 262.5035, 262.4846, 262.5167, 
    262.5474, 262.5988, 262.5903, 262.613, 262.5159, 262.5804, 262.4739, 
    262.503, 262.2712, 262.1833, 262.1456, 262.1128, 262.0327, 262.088, 
    262.0662, 262.1181, 262.151, 262.1347, 262.235, 262.1962, 262.4016, 
    262.313, 262.5438, 262.4885, 262.557, 262.5221, 262.5819, 262.5281, 
    262.6214, 262.6417, 262.6278, 262.6812, 262.5251, 262.585, 262.1342, 
    262.1369, 262.1493, 262.0948, 262.0915, 262.0417, 262.086, 262.1049, 
    262.1529, 262.1813, 262.2083, 262.2672, 262.3334, 262.4256, 262.4921, 
    262.5367, 262.5093, 262.5334, 262.5065, 262.4939, 262.6341, 262.5554, 
    262.6735, 262.667, 262.6135, 262.6677, 262.1388, 262.1235, 262.0704, 
    262.1119, 262.0362, 262.0786, 262.1029, 262.1969, 262.2177, 262.2365, 
    262.2743, 262.3228, 262.4076, 262.4816, 262.5492, 262.5442, 262.5459, 
    262.561, 262.5237, 262.5671, 262.5744, 262.5554, 262.6661, 262.6345, 
    262.6669, 262.6463, 262.1285, 262.1542, 262.1403, 262.1664, 262.148, 
    262.2295, 262.2541, 262.3689, 262.3218, 262.3968, 262.3295, 262.3414, 
    262.3991, 262.3331, 262.4774, 262.3796, 262.5616, 262.4636, 262.5677, 
    262.5489, 262.5801, 262.6081, 262.6434, 262.7083, 262.6933, 262.7477, 
    262.1925, 262.2259, 262.223, 262.2576, 262.2834, 262.3393, 262.4287, 
    262.3953, 262.4569, 262.4694, 262.3756, 262.433, 262.2479, 262.2778, 
    262.26, 262.1952, 262.403, 262.2962, 262.4932, 262.4353, 262.6041, 
    262.5202, 262.685, 262.7554, 262.8217, 262.899, 262.2438, 262.2215, 
    262.2617, 262.3178, 262.3699, 262.4389, 262.446, 262.4589, 262.4925, 
    262.5208, 262.463, 262.5278, 262.2847, 262.412, 262.2129, 262.2727, 
    262.3145, 262.2962, 262.3915, 262.4136, 262.5048, 262.4577, 262.738, 
    262.614, 262.9579, 262.8619, 262.2135, 262.2437, 262.3499, 262.2994, 
    262.4435, 262.479, 262.5079, 262.5448, 262.5488, 262.5707, 262.5349, 
    262.5693, 262.439, 262.4973, 262.3378, 262.3766, 262.3588, 262.3391, 
    262.3997, 262.4639, 262.4653, 262.486, 262.5441, 262.4441, 262.7538, 
    262.5625, 262.277, 262.3357, 262.3441, 262.3214, 262.4755, 262.4195, 
    262.5702, 262.5295, 262.5961, 262.563, 262.5581, 262.5156, 262.4891, 
    262.4221, 262.3679, 262.3247, 262.3347, 262.3822, 262.4678, 262.5492, 
    262.5313, 262.5911, 262.433, 262.4993, 262.4737, 262.5405, 262.3944, 
    262.5186, 262.3625, 262.3763, 262.4184, 262.5038, 262.5227, 262.5428, 
    262.5304, 262.47, 262.4602, 262.4174, 262.4059, 262.3733, 262.3463, 
    262.3709, 262.3968, 262.4701, 262.5363, 262.6085, 262.6262, 262.7104, 
    262.6418, 262.7549, 262.6586, 262.8253, 262.5259, 262.6559, 262.4204, 
    262.4458, 262.4916, 262.597, 262.5402, 262.6066, 262.4598, 262.3838, 
    262.3641, 262.3273, 262.365, 262.3619, 262.3979, 262.3864, 262.4725, 
    262.4261, 262.558, 262.6061, 262.7419, 262.8251, 262.9099, 262.9472, 
    262.9586, 262.9633 ;

 FIRE_R =
  262.0479, 262.1248, 262.1099, 262.1719, 262.1375, 262.1782, 262.0635, 
    262.1279, 262.0868, 262.0548, 262.292, 262.1747, 262.414, 262.3393, 
    262.5274, 262.4026, 262.5526, 262.5238, 262.6105, 262.5857, 262.6965, 
    262.622, 262.754, 262.6787, 262.6905, 262.6195, 262.1985, 262.2773, 
    262.1937, 262.205, 262.2, 262.1382, 262.1071, 262.042, 262.0538, 
    262.1017, 262.2101, 262.1733, 262.2658, 262.2637, 262.3669, 262.3204, 
    262.4936, 262.4443, 262.5867, 262.5509, 262.5851, 262.5747, 262.5852, 
    262.5327, 262.5551, 262.5089, 262.3291, 262.382, 262.2244, 262.1293, 
    262.0663, 262.0215, 262.0278, 262.0399, 262.1019, 262.1603, 262.2047, 
    262.2341, 262.2634, 262.3519, 262.3988, 262.5035, 262.4846, 262.5167, 
    262.5474, 262.5988, 262.5903, 262.613, 262.5159, 262.5804, 262.4739, 
    262.503, 262.2712, 262.1833, 262.1456, 262.1128, 262.0327, 262.088, 
    262.0662, 262.1181, 262.151, 262.1347, 262.235, 262.1962, 262.4016, 
    262.313, 262.5438, 262.4885, 262.557, 262.5221, 262.5819, 262.5281, 
    262.6214, 262.6417, 262.6278, 262.6812, 262.5251, 262.585, 262.1342, 
    262.1369, 262.1493, 262.0948, 262.0915, 262.0417, 262.086, 262.1049, 
    262.1529, 262.1813, 262.2083, 262.2672, 262.3334, 262.4256, 262.4921, 
    262.5367, 262.5093, 262.5334, 262.5065, 262.4939, 262.6341, 262.5554, 
    262.6735, 262.667, 262.6135, 262.6677, 262.1388, 262.1235, 262.0704, 
    262.1119, 262.0362, 262.0786, 262.1029, 262.1969, 262.2177, 262.2365, 
    262.2743, 262.3228, 262.4076, 262.4816, 262.5492, 262.5442, 262.5459, 
    262.561, 262.5237, 262.5671, 262.5744, 262.5554, 262.6661, 262.6345, 
    262.6669, 262.6463, 262.1285, 262.1542, 262.1403, 262.1664, 262.148, 
    262.2295, 262.2541, 262.3689, 262.3218, 262.3968, 262.3295, 262.3414, 
    262.3991, 262.3331, 262.4774, 262.3796, 262.5616, 262.4636, 262.5677, 
    262.5489, 262.5801, 262.6081, 262.6434, 262.7083, 262.6933, 262.7477, 
    262.1925, 262.2259, 262.223, 262.2576, 262.2834, 262.3393, 262.4287, 
    262.3953, 262.4569, 262.4694, 262.3756, 262.433, 262.2479, 262.2778, 
    262.26, 262.1952, 262.403, 262.2962, 262.4932, 262.4353, 262.6041, 
    262.5202, 262.685, 262.7554, 262.8217, 262.899, 262.2438, 262.2215, 
    262.2617, 262.3178, 262.3699, 262.4389, 262.446, 262.4589, 262.4925, 
    262.5208, 262.463, 262.5278, 262.2847, 262.412, 262.2129, 262.2727, 
    262.3145, 262.2962, 262.3915, 262.4136, 262.5048, 262.4577, 262.738, 
    262.614, 262.9579, 262.8619, 262.2135, 262.2437, 262.3499, 262.2994, 
    262.4435, 262.479, 262.5079, 262.5448, 262.5488, 262.5707, 262.5349, 
    262.5693, 262.439, 262.4973, 262.3378, 262.3766, 262.3588, 262.3391, 
    262.3997, 262.4639, 262.4653, 262.486, 262.5441, 262.4441, 262.7538, 
    262.5625, 262.277, 262.3357, 262.3441, 262.3214, 262.4755, 262.4195, 
    262.5702, 262.5295, 262.5961, 262.563, 262.5581, 262.5156, 262.4891, 
    262.4221, 262.3679, 262.3247, 262.3347, 262.3822, 262.4678, 262.5492, 
    262.5313, 262.5911, 262.433, 262.4993, 262.4737, 262.5405, 262.3944, 
    262.5186, 262.3625, 262.3763, 262.4184, 262.5038, 262.5227, 262.5428, 
    262.5304, 262.47, 262.4602, 262.4174, 262.4059, 262.3733, 262.3463, 
    262.3709, 262.3968, 262.4701, 262.5363, 262.6085, 262.6262, 262.7104, 
    262.6418, 262.7549, 262.6586, 262.8253, 262.5259, 262.6559, 262.4204, 
    262.4458, 262.4916, 262.597, 262.5402, 262.6066, 262.4598, 262.3838, 
    262.3641, 262.3273, 262.365, 262.3619, 262.3979, 262.3864, 262.4725, 
    262.4261, 262.558, 262.6061, 262.7419, 262.8251, 262.9099, 262.9472, 
    262.9586, 262.9633 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  336.1178, 337.0946, 336.9049, 337.6923, 337.2557, 337.7711, 336.3161, 
    337.1332, 336.6118, 336.2061, 339.2281, 337.7275, 340.788, 339.8279, 
    342.226, 340.6307, 342.5459, 342.1809, 343.2808, 342.9658, 344.3708, 
    343.4261, 345.0997, 344.1455, 344.2946, 343.3949, 338.0282, 339.0422, 
    337.9686, 338.1119, 338.0477, 337.2646, 336.8694, 336.0435, 336.1936, 
    336.8004, 338.1764, 337.7097, 338.8958, 338.8692, 340.1787, 339.5883, 
    341.7977, 341.1726, 342.9789, 342.5247, 342.9575, 342.8263, 342.9592, 
    342.293, 342.5784, 341.9924, 339.6988, 340.3702, 338.3579, 337.1518, 
    336.3519, 335.7837, 335.864, 336.017, 336.804, 337.5441, 338.1079, 
    338.4939, 338.8654, 339.9881, 340.5833, 341.9238, 341.6841, 342.0905, 
    342.4795, 343.1318, 343.0245, 343.3117, 342.0802, 342.8986, 341.5474, 
    341.9169, 338.9645, 337.8357, 337.3581, 336.9413, 335.9257, 336.627, 
    336.3505, 337.0086, 337.4265, 337.2199, 338.5042, 337.9994, 340.6186, 
    339.4946, 342.4342, 341.7333, 342.6022, 342.159, 342.9182, 342.2349, 
    343.4188, 343.6762, 343.5002, 344.1768, 342.197, 342.9573, 337.214, 
    337.2477, 337.4048, 336.7141, 336.6719, 336.0393, 336.6024, 336.8419, 
    337.4508, 337.8105, 338.1526, 338.9135, 339.7528, 340.9355, 341.7787, 
    342.3437, 341.9974, 342.3031, 341.9613, 341.8011, 343.5796, 342.581, 
    344.0796, 343.9967, 343.3185, 344.0061, 337.2714, 337.0775, 336.4037, 
    336.931, 335.9704, 336.5079, 336.8168, 338.0093, 338.2718, 338.5234, 
    339.0032, 339.6185, 340.7065, 341.6453, 342.5022, 342.4395, 342.4616, 
    342.6528, 342.1789, 342.7306, 342.823, 342.5811, 343.9856, 343.5845, 
    343.995, 343.7338, 337.1406, 337.4668, 337.2905, 337.622, 337.3883, 
    338.4357, 338.7469, 340.2035, 339.6063, 340.5572, 339.7031, 339.8544, 
    340.5875, 339.7494, 341.5932, 340.3397, 342.6602, 341.4172, 342.738, 
    342.4985, 342.8952, 343.2503, 343.6972, 344.521, 344.3304, 345.0195, 
    337.9534, 338.3763, 338.3394, 338.7912, 339.1186, 339.8284, 340.9751, 
    340.5384, 341.3328, 341.4904, 340.2883, 341.0295, 338.6686, 339.0483, 
    338.8225, 337.9865, 340.6364, 339.2812, 341.7926, 341.0589, 343.1996, 
    342.1349, 344.2253, 345.1175, 345.9584, 346.9388, 338.6165, 338.3201, 
    338.844, 339.5555, 340.2166, 341.1036, 341.1936, 341.3579, 341.784, 
    342.142, 341.4096, 342.2318, 339.1357, 340.7632, 338.2111, 338.9829, 
    339.5137, 339.2813, 340.4896, 340.7832, 341.9392, 341.3419, 344.897, 
    343.3248, 347.6862, 346.468, 338.2196, 338.6156, 339.9619, 339.3215, 
    341.1624, 341.6129, 341.9795, 342.4473, 342.4981, 342.7753, 342.321, 
    342.7575, 341.1055, 341.8439, 339.8085, 340.3016, 340.0749, 339.8259, 
    340.5942, 341.421, 341.4391, 341.7011, 342.4384, 341.1698, 345.0988, 
    342.6721, 339.0376, 339.7822, 339.8892, 339.6007, 341.5677, 340.8584, 
    342.7686, 342.2526, 343.0981, 342.678, 342.6161, 342.0765, 341.7403, 
    340.8908, 340.1906, 339.6426, 339.7701, 340.372, 341.4712, 342.5024, 
    342.2765, 343.0339, 341.0296, 341.8699, 341.545, 342.3923, 340.5269, 
    342.1151, 340.1229, 340.297, 340.8443, 341.9265, 342.1667, 342.4222, 
    342.2647, 341.4989, 341.3737, 340.8314, 340.6723, 340.2591, 339.9167, 
    340.2294, 340.5576, 341.4995, 342.3395, 343.2552, 343.4795, 344.5474, 
    343.6773, 345.1122, 343.8912, 346.0049, 342.2074, 343.8564, 340.869, 
    341.1911, 341.7731, 343.1086, 342.3883, 343.231, 341.3688, 340.3925, 
    340.1428, 339.6758, 340.1535, 340.1147, 340.5716, 340.4248, 341.5305, 
    340.9415, 342.6144, 343.2245, 344.9471, 346.002, 347.0763, 347.5501, 
    347.6943, 347.7546 ;

 FSH_G =
  342.8148, 343.7922, 343.6024, 344.3902, 343.9534, 344.4691, 343.0132, 
    343.8308, 343.3091, 342.9032, 345.9269, 344.4254, 347.4878, 346.5272, 
    348.9267, 347.3304, 349.2468, 348.8816, 349.9821, 349.6669, 351.0728, 
    350.1276, 351.8022, 350.8474, 350.9966, 350.0963, 344.7264, 345.7409, 
    344.6667, 344.8101, 344.7459, 343.9622, 343.5669, 342.7405, 342.8906, 
    343.4978, 344.8746, 344.4077, 345.5944, 345.5679, 346.8781, 346.2874, 
    348.4981, 347.8727, 349.6801, 349.2256, 349.6586, 349.5274, 349.6603, 
    348.9938, 349.2793, 348.6929, 346.3979, 347.0698, 345.0562, 343.8495, 
    343.049, 342.4805, 342.5608, 342.714, 343.5014, 344.242, 344.8061, 
    345.1923, 345.564, 346.6874, 347.2831, 348.6243, 348.3844, 348.7912, 
    349.1804, 349.833, 349.7257, 350.0131, 348.7808, 349.5997, 348.2477, 
    348.6174, 345.6631, 344.5338, 344.0558, 343.6388, 342.6226, 343.3243, 
    343.0477, 343.7061, 344.1242, 343.9175, 345.2026, 344.6975, 347.3183, 
    346.1937, 349.135, 348.4337, 349.3031, 348.8596, 349.6193, 348.9356, 
    350.1202, 350.3778, 350.2017, 350.8788, 348.8976, 349.6584, 343.9117, 
    343.9454, 344.1026, 343.4114, 343.3692, 342.7363, 343.2997, 343.5394, 
    344.1486, 344.5086, 344.8508, 345.6122, 346.452, 347.6354, 348.4791, 
    349.0444, 348.6979, 349.0038, 348.6618, 348.5016, 350.2812, 349.2819, 
    350.7814, 350.6985, 350.0198, 350.7079, 343.9691, 343.7751, 343.1009, 
    343.6285, 342.6674, 343.2051, 343.5142, 344.7075, 344.9701, 345.2219, 
    345.7019, 346.3177, 347.4063, 348.3456, 349.2031, 349.1403, 349.1624, 
    349.3537, 348.8795, 349.4316, 349.524, 349.282, 350.6874, 350.286, 
    350.6967, 350.4355, 343.8382, 344.1647, 343.9882, 344.3199, 344.0861, 
    345.1341, 345.4455, 346.903, 346.3054, 347.2569, 346.4023, 346.5536, 
    347.2871, 346.4486, 348.2935, 347.0392, 349.3611, 348.1174, 349.439, 
    349.1994, 349.5963, 349.9516, 350.3988, 351.2231, 351.0323, 351.7219, 
    344.6515, 345.0747, 345.0378, 345.4898, 345.8174, 346.5276, 347.675, 
    347.2381, 348.033, 348.1906, 346.9878, 347.7295, 345.3671, 345.7471, 
    345.5211, 344.6847, 347.3362, 345.9801, 348.493, 347.7589, 349.9009, 
    348.8355, 350.9272, 351.8199, 352.6614, 353.6424, 345.315, 345.0185, 
    345.5426, 346.2546, 346.916, 347.8036, 347.8937, 348.0581, 348.4844, 
    348.8427, 348.1097, 348.9325, 345.8345, 347.463, 344.9094, 345.6817, 
    346.2128, 345.9802, 347.1893, 347.483, 348.6397, 348.0421, 351.5993, 
    350.0261, 354.3902, 353.1713, 344.9179, 345.3141, 346.6612, 346.0204, 
    347.8624, 348.3132, 348.68, 349.1481, 349.1989, 349.4763, 349.0217, 
    349.4585, 347.8055, 348.5443, 346.5077, 347.0011, 346.7743, 346.5251, 
    347.2939, 348.1212, 348.1393, 348.4015, 349.1392, 347.8699, 351.8011, 
    349.3731, 345.7364, 346.4814, 346.5885, 346.2998, 348.268, 347.5582, 
    349.4696, 348.9533, 349.7994, 349.3789, 349.317, 348.7771, 348.4407, 
    347.5907, 346.89, 346.3417, 346.4693, 347.0715, 348.1714, 349.2033, 
    348.9772, 349.7351, 347.7296, 348.5704, 348.2453, 349.0931, 347.2266, 
    348.8157, 346.8224, 346.9965, 347.5442, 348.627, 348.8674, 349.123, 
    348.9654, 348.1992, 348.0739, 347.5312, 347.372, 346.9586, 346.6161, 
    346.9289, 347.2573, 348.1997, 349.0403, 349.9565, 350.181, 351.2495, 
    350.3789, 351.8146, 350.5928, 352.7079, 348.9081, 350.558, 347.5688, 
    347.8912, 348.4735, 349.8098, 349.0891, 349.9323, 348.069, 347.092, 
    346.8423, 346.375, 346.8529, 346.8141, 347.2713, 347.1244, 348.2307, 
    347.6414, 349.3153, 349.9258, 351.6494, 352.705, 353.78, 354.2541, 
    354.3984, 354.4587 ;

 FSH_NODYNLNDUSE =
  336.1178, 337.0946, 336.9049, 337.6923, 337.2557, 337.7711, 336.3161, 
    337.1332, 336.6118, 336.2061, 339.2281, 337.7275, 340.788, 339.8279, 
    342.226, 340.6307, 342.5459, 342.1809, 343.2808, 342.9658, 344.3708, 
    343.4261, 345.0997, 344.1455, 344.2946, 343.3949, 338.0282, 339.0422, 
    337.9686, 338.1119, 338.0477, 337.2646, 336.8694, 336.0435, 336.1936, 
    336.8004, 338.1764, 337.7097, 338.8958, 338.8692, 340.1787, 339.5883, 
    341.7977, 341.1726, 342.9789, 342.5247, 342.9575, 342.8263, 342.9592, 
    342.293, 342.5784, 341.9924, 339.6988, 340.3702, 338.3579, 337.1518, 
    336.3519, 335.7837, 335.864, 336.017, 336.804, 337.5441, 338.1079, 
    338.4939, 338.8654, 339.9881, 340.5833, 341.9238, 341.6841, 342.0905, 
    342.4795, 343.1318, 343.0245, 343.3117, 342.0802, 342.8986, 341.5474, 
    341.9169, 338.9645, 337.8357, 337.3581, 336.9413, 335.9257, 336.627, 
    336.3505, 337.0086, 337.4265, 337.2199, 338.5042, 337.9994, 340.6186, 
    339.4946, 342.4342, 341.7333, 342.6022, 342.159, 342.9182, 342.2349, 
    343.4188, 343.6762, 343.5002, 344.1768, 342.197, 342.9573, 337.214, 
    337.2477, 337.4048, 336.7141, 336.6719, 336.0393, 336.6024, 336.8419, 
    337.4508, 337.8105, 338.1526, 338.9135, 339.7528, 340.9355, 341.7787, 
    342.3437, 341.9974, 342.3031, 341.9613, 341.8011, 343.5796, 342.581, 
    344.0796, 343.9967, 343.3185, 344.0061, 337.2714, 337.0775, 336.4037, 
    336.931, 335.9704, 336.5079, 336.8168, 338.0093, 338.2718, 338.5234, 
    339.0032, 339.6185, 340.7065, 341.6453, 342.5022, 342.4395, 342.4616, 
    342.6528, 342.1789, 342.7306, 342.823, 342.5811, 343.9856, 343.5845, 
    343.995, 343.7338, 337.1406, 337.4668, 337.2905, 337.622, 337.3883, 
    338.4357, 338.7469, 340.2035, 339.6063, 340.5572, 339.7031, 339.8544, 
    340.5875, 339.7494, 341.5932, 340.3397, 342.6602, 341.4172, 342.738, 
    342.4985, 342.8952, 343.2503, 343.6972, 344.521, 344.3304, 345.0195, 
    337.9534, 338.3763, 338.3394, 338.7912, 339.1186, 339.8284, 340.9751, 
    340.5384, 341.3328, 341.4904, 340.2883, 341.0295, 338.6686, 339.0483, 
    338.8225, 337.9865, 340.6364, 339.2812, 341.7926, 341.0589, 343.1996, 
    342.1349, 344.2253, 345.1175, 345.9584, 346.9388, 338.6165, 338.3201, 
    338.844, 339.5555, 340.2166, 341.1036, 341.1936, 341.3579, 341.784, 
    342.142, 341.4096, 342.2318, 339.1357, 340.7632, 338.2111, 338.9829, 
    339.5137, 339.2813, 340.4896, 340.7832, 341.9392, 341.3419, 344.897, 
    343.3248, 347.6862, 346.468, 338.2196, 338.6156, 339.9619, 339.3215, 
    341.1624, 341.6129, 341.9795, 342.4473, 342.4981, 342.7753, 342.321, 
    342.7575, 341.1055, 341.8439, 339.8085, 340.3016, 340.0749, 339.8259, 
    340.5942, 341.421, 341.4391, 341.7011, 342.4384, 341.1698, 345.0988, 
    342.6721, 339.0376, 339.7822, 339.8892, 339.6007, 341.5677, 340.8584, 
    342.7686, 342.2526, 343.0981, 342.678, 342.6161, 342.0765, 341.7403, 
    340.8908, 340.1906, 339.6426, 339.7701, 340.372, 341.4712, 342.5024, 
    342.2765, 343.0339, 341.0296, 341.8699, 341.545, 342.3923, 340.5269, 
    342.1151, 340.1229, 340.297, 340.8443, 341.9265, 342.1667, 342.4222, 
    342.2647, 341.4989, 341.3737, 340.8314, 340.6723, 340.2591, 339.9167, 
    340.2294, 340.5576, 341.4995, 342.3395, 343.2552, 343.4795, 344.5474, 
    343.6773, 345.1122, 343.8912, 346.0049, 342.2074, 343.8564, 340.869, 
    341.1911, 341.7731, 343.1086, 342.3883, 343.231, 341.3688, 340.3925, 
    340.1428, 339.6758, 340.1535, 340.1147, 340.5716, 340.4248, 341.5305, 
    340.9415, 342.6144, 343.2245, 344.9471, 346.002, 347.0763, 347.5501, 
    347.6943, 347.7546 ;

 FSH_R =
  336.1178, 337.0946, 336.9049, 337.6923, 337.2557, 337.7711, 336.3161, 
    337.1332, 336.6118, 336.2061, 339.2281, 337.7275, 340.788, 339.8279, 
    342.226, 340.6307, 342.5459, 342.1809, 343.2808, 342.9658, 344.3708, 
    343.4261, 345.0997, 344.1455, 344.2946, 343.3949, 338.0282, 339.0422, 
    337.9686, 338.1119, 338.0477, 337.2646, 336.8694, 336.0435, 336.1936, 
    336.8004, 338.1764, 337.7097, 338.8958, 338.8692, 340.1787, 339.5883, 
    341.7977, 341.1726, 342.9789, 342.5247, 342.9575, 342.8263, 342.9592, 
    342.293, 342.5784, 341.9924, 339.6988, 340.3702, 338.3579, 337.1518, 
    336.3519, 335.7837, 335.864, 336.017, 336.804, 337.5441, 338.1079, 
    338.4939, 338.8654, 339.9881, 340.5833, 341.9238, 341.6841, 342.0905, 
    342.4795, 343.1318, 343.0245, 343.3117, 342.0802, 342.8986, 341.5474, 
    341.9169, 338.9645, 337.8357, 337.3581, 336.9413, 335.9257, 336.627, 
    336.3505, 337.0086, 337.4265, 337.2199, 338.5042, 337.9994, 340.6186, 
    339.4946, 342.4342, 341.7333, 342.6022, 342.159, 342.9182, 342.2349, 
    343.4188, 343.6762, 343.5002, 344.1768, 342.197, 342.9573, 337.214, 
    337.2477, 337.4048, 336.7141, 336.6719, 336.0393, 336.6024, 336.8419, 
    337.4508, 337.8105, 338.1526, 338.9135, 339.7528, 340.9355, 341.7787, 
    342.3437, 341.9974, 342.3031, 341.9613, 341.8011, 343.5796, 342.581, 
    344.0796, 343.9967, 343.3185, 344.0061, 337.2714, 337.0775, 336.4037, 
    336.931, 335.9704, 336.5079, 336.8168, 338.0093, 338.2718, 338.5234, 
    339.0032, 339.6185, 340.7065, 341.6453, 342.5022, 342.4395, 342.4616, 
    342.6528, 342.1789, 342.7306, 342.823, 342.5811, 343.9856, 343.5845, 
    343.995, 343.7338, 337.1406, 337.4668, 337.2905, 337.622, 337.3883, 
    338.4357, 338.7469, 340.2035, 339.6063, 340.5572, 339.7031, 339.8544, 
    340.5875, 339.7494, 341.5932, 340.3397, 342.6602, 341.4172, 342.738, 
    342.4985, 342.8952, 343.2503, 343.6972, 344.521, 344.3304, 345.0195, 
    337.9534, 338.3763, 338.3394, 338.7912, 339.1186, 339.8284, 340.9751, 
    340.5384, 341.3328, 341.4904, 340.2883, 341.0295, 338.6686, 339.0483, 
    338.8225, 337.9865, 340.6364, 339.2812, 341.7926, 341.0589, 343.1996, 
    342.1349, 344.2253, 345.1175, 345.9584, 346.9388, 338.6165, 338.3201, 
    338.844, 339.5555, 340.2166, 341.1036, 341.1936, 341.3579, 341.784, 
    342.142, 341.4096, 342.2318, 339.1357, 340.7632, 338.2111, 338.9829, 
    339.5137, 339.2813, 340.4896, 340.7832, 341.9392, 341.3419, 344.897, 
    343.3248, 347.6862, 346.468, 338.2196, 338.6156, 339.9619, 339.3215, 
    341.1624, 341.6129, 341.9795, 342.4473, 342.4981, 342.7753, 342.321, 
    342.7575, 341.1055, 341.8439, 339.8085, 340.3016, 340.0749, 339.8259, 
    340.5942, 341.421, 341.4391, 341.7011, 342.4384, 341.1698, 345.0988, 
    342.6721, 339.0376, 339.7822, 339.8892, 339.6007, 341.5677, 340.8584, 
    342.7686, 342.2526, 343.0981, 342.678, 342.6161, 342.0765, 341.7403, 
    340.8908, 340.1906, 339.6426, 339.7701, 340.372, 341.4712, 342.5024, 
    342.2765, 343.0339, 341.0296, 341.8699, 341.545, 342.3923, 340.5269, 
    342.1151, 340.1229, 340.297, 340.8443, 341.9265, 342.1667, 342.4222, 
    342.2647, 341.4989, 341.3737, 340.8314, 340.6723, 340.2591, 339.9167, 
    340.2294, 340.5576, 341.4995, 342.3395, 343.2552, 343.4795, 344.5474, 
    343.6773, 345.1122, 343.8912, 346.0049, 342.2074, 343.8564, 340.869, 
    341.1911, 341.7731, 343.1086, 342.3883, 343.231, 341.3688, 340.3925, 
    340.1428, 339.6758, 340.1535, 340.1147, 340.5716, 340.4248, 341.5305, 
    340.9415, 342.6144, 343.2245, 344.9471, 346.002, 347.0763, 347.5501, 
    347.6943, 347.7546 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.697002, -6.697589, -6.697478, -6.697947, -6.69769, -6.697994, -6.697126, 
    -6.697608, -6.697303, -6.697061, -6.698845, -6.697969, -6.699804, 
    -6.699235, -6.700679, -6.699708, -6.700878, -6.700662, -6.701337, 
    -6.701145, -6.701988, -6.701427, -6.702444, -6.701859, -6.701947, 
    -6.701406, -6.698155, -6.698733, -6.698118, -6.698201, -6.698166, 
    -6.697692, -6.697446, -6.696964, -6.697054, -6.697412, -6.698239, 
    -6.697965, -6.698677, -6.698661, -6.699449, -6.699093, -6.700428, 
    -6.700051, -6.701153, -6.700873, -6.701138, -6.701059, -6.701139, 
    -6.70073, -6.700904, -6.700549, -6.699157, -6.699562, -6.698351, 
    -6.69761, -6.697145, -6.696807, -6.696855, -6.696944, -6.697413, 
    -6.697865, -6.698206, -6.698433, -6.698658, -6.699314, -6.699685, 
    -6.7005, -6.700361, -6.700603, -6.700846, -6.701243, -6.70118, -6.701352, 
    -6.700603, -6.701097, -6.700281, -6.700502, -6.698684, -6.69804, 
    -6.697736, -6.697498, -6.696891, -6.697308, -6.697143, -6.697544, 
    -6.697793, -6.697671, -6.69844, -6.698139, -6.699707, -6.699031, 
    -6.700818, -6.70039, -6.700922, -6.700652, -6.701111, -6.700698, 
    -6.70142, -6.701573, -6.701468, -6.701885, -6.700675, -6.701134, 
    -6.697666, -6.697686, -6.697782, -6.69736, -6.697336, -6.69696, 
    -6.697298, -6.697439, -6.697811, -6.698025, -6.69823, -6.698684, 
    -6.699185, -6.699899, -6.700418, -6.700765, -6.700554, -6.70074, 
    -6.700531, -6.700435, -6.701513, -6.700904, -6.701825, -6.701775, 
    -6.701355, -6.701781, -6.697701, -6.697586, -6.697177, -6.697497, 
    -6.69692, -6.697238, -6.697419, -6.698137, -6.698304, -6.698448, 
    -6.69874, -6.699111, -6.699761, -6.700333, -6.700862, -6.700824, 
    -6.700837, -6.700952, -6.700663, -6.700999, -6.701052, -6.700908, 
    -6.701768, -6.701523, -6.701774, -6.701615, -6.697624, -6.697818, 
    -6.697713, -6.697909, -6.697768, -6.698388, -6.698574, -6.699455, 
    -6.699101, -6.699674, -6.699162, -6.699251, -6.699677, -6.699193, 
    -6.700294, -6.699533, -6.700956, -6.70018, -6.701004, -6.70086, 
    -6.701102, -6.701315, -6.701591, -6.70209, -6.701976, -6.7024, -6.698112, 
    -6.698361, -6.698346, -6.698612, -6.698807, -6.69924, -6.699927, 
    -6.69967, -6.700149, -6.700243, -6.69952, -6.699957, -6.698534, 
    -6.698756, -6.698628, -6.698128, -6.69972, -6.698897, -6.700425, 
    -6.699979, -6.701284, -6.700627, -6.701911, -6.702445, -6.70298, 
    -6.70357, -6.698505, -6.698334, -6.698646, -6.699064, -6.699472, 
    -6.700005, -6.700064, -6.700161, -6.700424, -6.700642, -6.700186, 
    -6.700696, -6.698794, -6.699795, -6.698264, -6.698715, -6.699042, 
    -6.698905, -6.699643, -6.699815, -6.700511, -6.700155, -6.702307, 
    -6.701351, -6.704042, -6.703283, -6.698273, -6.698508, -6.699314, 
    -6.698931, -6.700045, -6.700316, -6.700543, -6.700823, -6.700858, 
    -6.701025, -6.700751, -6.701016, -6.700006, -6.700459, -6.699229, 
    -6.699524, -6.69939, -6.69924, -6.699705, -6.700191, -6.700213, 
    -6.700367, -6.700783, -6.700049, -6.702411, -6.700931, -6.698762, 
    -6.699199, -6.699275, -6.699103, -6.700289, -6.699857, -6.701022, 
    -6.700709, -6.701225, -6.700968, -6.700929, -6.700602, -6.700395, 
    -6.699875, -6.699455, -6.699129, -6.699206, -6.699564, -6.700224, 
    -6.700856, -6.700716, -6.701186, -6.699964, -6.700469, -6.70027, 
    -6.700792, -6.699661, -6.700591, -6.69942, -6.699524, -6.699849, 
    -6.700497, -6.700656, -6.700808, -6.700716, -6.700243, -6.70017, 
    -6.699843, -6.699748, -6.699502, -6.699295, -6.699482, -6.699677, 
    -6.700247, -6.700757, -6.701317, -6.701459, -6.702088, -6.70156, 
    -6.702417, -6.701666, -6.702979, -6.700662, -6.701666, -6.699867, 
    -6.700063, -6.700406, -6.701217, -6.70079, -6.701295, -6.700168, 
    -6.699572, -6.699431, -6.699147, -6.699438, -6.699414, -6.699692, 
    -6.699604, -6.700266, -6.699911, -6.700925, -6.701294, -6.702351, 
    -6.702995, -6.70367, -6.703963, -6.704053, -6.70409 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_NIT =
  2.302195e-14, 2.322149e-14, 2.318263e-14, 2.334409e-14, 2.325445e-14, 
    2.336027e-14, 2.306232e-14, 2.322941e-14, 2.312267e-14, 2.303986e-14, 
    2.36591e-14, 2.335129e-14, 2.398116e-14, 2.378316e-14, 2.42822e-14, 
    2.395028e-14, 2.434942e-14, 2.42726e-14, 2.450423e-14, 2.443775e-14, 
    2.473528e-14, 2.453494e-14, 2.489029e-14, 2.468736e-14, 2.471904e-14, 
    2.452833e-14, 2.341309e-14, 2.362068e-14, 2.340081e-14, 2.343035e-14, 
    2.341709e-14, 2.325628e-14, 2.317546e-14, 2.300672e-14, 2.30373e-14, 
    2.316126e-14, 2.344361e-14, 2.334757e-14, 2.359004e-14, 2.358455e-14, 
    2.385602e-14, 2.373341e-14, 2.419218e-14, 2.406132e-14, 2.444052e-14, 
    2.434485e-14, 2.443601e-14, 2.440835e-14, 2.443637e-14, 2.429615e-14, 
    2.435616e-14, 2.423297e-14, 2.375638e-14, 2.389593e-14, 2.348098e-14, 
    2.323332e-14, 2.306962e-14, 2.295383e-14, 2.297017e-14, 2.300136e-14, 
    2.316199e-14, 2.331356e-14, 2.342942e-14, 2.350709e-14, 2.358375e-14, 
    2.38166e-14, 2.394036e-14, 2.421868e-14, 2.416833e-14, 2.425366e-14, 
    2.433534e-14, 2.447279e-14, 2.445014e-14, 2.451079e-14, 2.42514e-14, 
    2.442362e-14, 2.413965e-14, 2.421714e-14, 2.360461e-14, 2.337347e-14, 
    2.327556e-14, 2.319007e-14, 2.298275e-14, 2.312581e-14, 2.306935e-14, 
    2.320378e-14, 2.328941e-14, 2.324703e-14, 2.350921e-14, 2.340709e-14, 
    2.394769e-14, 2.371404e-14, 2.432581e-14, 2.417866e-14, 2.436114e-14, 
    2.426793e-14, 2.442775e-14, 2.428389e-14, 2.453338e-14, 2.458789e-14, 
    2.455063e-14, 2.469391e-14, 2.427591e-14, 2.443598e-14, 2.324586e-14, 
    2.325277e-14, 2.328496e-14, 2.31436e-14, 2.313497e-14, 2.300586e-14, 
    2.312072e-14, 2.316972e-14, 2.329438e-14, 2.336827e-14, 2.343863e-14, 
    2.359373e-14, 2.37676e-14, 2.401186e-14, 2.418818e-14, 2.430674e-14, 
    2.4234e-14, 2.429821e-14, 2.422643e-14, 2.419282e-14, 2.456745e-14, 
    2.435671e-14, 2.467327e-14, 2.46557e-14, 2.451221e-14, 2.465767e-14, 
    2.325762e-14, 2.321787e-14, 2.308017e-14, 2.318789e-14, 2.299182e-14, 
    2.310145e-14, 2.316462e-14, 2.340921e-14, 2.346314e-14, 2.35132e-14, 
    2.361224e-14, 2.373966e-14, 2.396407e-14, 2.416025e-14, 2.434009e-14, 
    2.432688e-14, 2.433153e-14, 2.437178e-14, 2.427212e-14, 2.438816e-14, 
    2.440766e-14, 2.435668e-14, 2.465334e-14, 2.456839e-14, 2.465531e-14, 
    2.459998e-14, 2.323078e-14, 2.329769e-14, 2.326152e-14, 2.332955e-14, 
    2.32816e-14, 2.349519e-14, 2.355943e-14, 2.386126e-14, 2.373714e-14, 
    2.393485e-14, 2.375718e-14, 2.378861e-14, 2.394129e-14, 2.376676e-14, 
    2.414939e-14, 2.388961e-14, 2.437334e-14, 2.411263e-14, 2.438973e-14, 
    2.433929e-14, 2.442282e-14, 2.449777e-14, 2.459224e-14, 2.476705e-14, 
    2.472651e-14, 2.487308e-14, 2.339763e-14, 2.348476e-14, 2.347708e-14, 
    2.356844e-14, 2.363612e-14, 2.378319e-14, 2.402007e-14, 2.393084e-14, 
    2.409478e-14, 2.412776e-14, 2.387874e-14, 2.403146e-14, 2.354314e-14, 
    2.362167e-14, 2.35749e-14, 2.340445e-14, 2.395135e-14, 2.366983e-14, 
    2.419106e-14, 2.403752e-14, 2.448707e-14, 2.426294e-14, 2.47042e-14, 
    2.489412e-14, 2.507359e-14, 2.528417e-14, 2.353239e-14, 2.34731e-14, 
    2.357931e-14, 2.372668e-14, 2.386387e-14, 2.40469e-14, 2.406567e-14, 
    2.410005e-14, 2.418924e-14, 2.426437e-14, 2.411092e-14, 2.428321e-14, 
    2.363988e-14, 2.397587e-14, 2.345066e-14, 2.360815e-14, 2.371794e-14, 
    2.366975e-14, 2.392062e-14, 2.397994e-14, 2.422184e-14, 2.409663e-14, 
    2.484716e-14, 2.451359e-14, 2.544515e-14, 2.518295e-14, 2.345239e-14, 
    2.353217e-14, 2.381097e-14, 2.36781e-14, 2.405914e-14, 2.415343e-14, 
    2.423022e-14, 2.432858e-14, 2.433921e-14, 2.43976e-14, 2.430195e-14, 
    2.439381e-14, 2.404726e-14, 2.42018e-14, 2.377899e-14, 2.388152e-14, 
    2.383432e-14, 2.37826e-14, 2.394241e-14, 2.411329e-14, 2.411696e-14, 
    2.417189e-14, 2.432702e-14, 2.406064e-14, 2.489035e-14, 2.437616e-14, 
    2.361934e-14, 2.377371e-14, 2.379581e-14, 2.373591e-14, 2.414396e-14, 
    2.399568e-14, 2.439617e-14, 2.428758e-14, 2.446563e-14, 2.437707e-14, 
    2.436405e-14, 2.425058e-14, 2.418007e-14, 2.400244e-14, 2.385842e-14, 
    2.374456e-14, 2.377101e-14, 2.389618e-14, 2.412376e-14, 2.434013e-14, 
    2.429264e-14, 2.445204e-14, 2.403135e-14, 2.420727e-14, 2.413919e-14, 
    2.431692e-14, 2.392846e-14, 2.425906e-14, 2.384433e-14, 2.388054e-14, 
    2.399274e-14, 2.421926e-14, 2.426955e-14, 2.432328e-14, 2.429011e-14, 
    2.412958e-14, 2.410333e-14, 2.398999e-14, 2.395873e-14, 2.387263e-14, 
    2.380145e-14, 2.386647e-14, 2.393484e-14, 2.412962e-14, 2.430587e-14, 
    2.44988e-14, 2.454615e-14, 2.477281e-14, 2.45882e-14, 2.489322e-14, 
    2.463374e-14, 2.508384e-14, 2.42783e-14, 2.46262e-14, 2.399785e-14, 
    2.406513e-14, 2.418706e-14, 2.446798e-14, 2.431612e-14, 2.449378e-14, 
    2.41023e-14, 2.39005e-14, 2.384844e-14, 2.375147e-14, 2.385066e-14, 
    2.384258e-14, 2.393768e-14, 2.39071e-14, 2.41361e-14, 2.401295e-14, 
    2.436368e-14, 2.449234e-14, 2.485766e-14, 2.508303e-14, 2.531357e-14, 
    2.54157e-14, 2.544683e-14, 2.545985e-14 ;

 F_NIT =
  3.836991e-11, 3.870249e-11, 3.863771e-11, 3.890682e-11, 3.875741e-11, 
    3.893379e-11, 3.84372e-11, 3.871568e-11, 3.853778e-11, 3.839976e-11, 
    3.943183e-11, 3.891881e-11, 3.996859e-11, 3.96386e-11, 4.047033e-11, 
    3.991713e-11, 4.058237e-11, 4.045433e-11, 4.084039e-11, 4.072958e-11, 
    4.122547e-11, 4.089157e-11, 4.148381e-11, 4.11456e-11, 4.11984e-11, 
    4.088055e-11, 3.902182e-11, 3.93678e-11, 3.900135e-11, 3.905058e-11, 
    3.902848e-11, 3.876047e-11, 3.862577e-11, 3.834453e-11, 3.83955e-11, 
    3.860211e-11, 3.907269e-11, 3.891261e-11, 3.931673e-11, 3.930758e-11, 
    3.976003e-11, 3.955569e-11, 4.032031e-11, 4.010219e-11, 4.07342e-11, 
    4.057475e-11, 4.072669e-11, 4.068058e-11, 4.072728e-11, 4.049358e-11, 
    4.05936e-11, 4.038829e-11, 3.959397e-11, 3.982656e-11, 3.913497e-11, 
    3.872221e-11, 3.844937e-11, 3.825638e-11, 3.828362e-11, 3.83356e-11, 
    3.860331e-11, 3.885593e-11, 3.904903e-11, 3.917848e-11, 3.930626e-11, 
    3.969433e-11, 3.99006e-11, 4.036447e-11, 4.028056e-11, 4.042277e-11, 
    4.05589e-11, 4.078798e-11, 4.075023e-11, 4.085132e-11, 4.0419e-11, 
    4.070604e-11, 4.023275e-11, 4.03619e-11, 3.934102e-11, 3.895579e-11, 
    3.87926e-11, 3.865011e-11, 3.830458e-11, 3.854301e-11, 3.844892e-11, 
    3.867296e-11, 3.881568e-11, 3.874506e-11, 3.918202e-11, 3.901182e-11, 
    3.991283e-11, 3.952339e-11, 4.054301e-11, 4.029776e-11, 4.06019e-11, 
    4.044656e-11, 4.071292e-11, 4.047315e-11, 4.088897e-11, 4.097982e-11, 
    4.091772e-11, 4.115652e-11, 4.045985e-11, 4.072663e-11, 3.874311e-11, 
    3.875462e-11, 3.880827e-11, 3.857267e-11, 3.855828e-11, 3.83431e-11, 
    3.853453e-11, 3.86162e-11, 3.882396e-11, 3.894711e-11, 3.906438e-11, 
    3.932289e-11, 3.961266e-11, 4.001976e-11, 4.031363e-11, 4.051124e-11, 
    4.039e-11, 4.049702e-11, 4.037739e-11, 4.032137e-11, 4.094575e-11, 
    4.059452e-11, 4.112212e-11, 4.109283e-11, 4.085369e-11, 4.109611e-11, 
    3.876269e-11, 3.869646e-11, 3.846694e-11, 3.864649e-11, 3.831969e-11, 
    3.850242e-11, 3.86077e-11, 3.901535e-11, 3.910524e-11, 3.918867e-11, 
    3.935373e-11, 3.95661e-11, 3.994012e-11, 4.026708e-11, 4.056681e-11, 
    4.05448e-11, 4.055255e-11, 4.061964e-11, 4.045353e-11, 4.064693e-11, 
    4.067944e-11, 4.059447e-11, 4.108889e-11, 4.094731e-11, 4.109219e-11, 
    4.099997e-11, 3.871797e-11, 3.882948e-11, 3.87692e-11, 3.888259e-11, 
    3.880267e-11, 3.915865e-11, 3.926571e-11, 3.976877e-11, 3.956191e-11, 
    3.989141e-11, 3.959531e-11, 3.964768e-11, 3.990215e-11, 3.961127e-11, 
    4.024899e-11, 3.981602e-11, 4.062224e-11, 4.018771e-11, 4.064955e-11, 
    4.056547e-11, 4.070471e-11, 4.082962e-11, 4.098706e-11, 4.127841e-11, 
    4.121084e-11, 4.145513e-11, 3.899605e-11, 3.914126e-11, 3.912847e-11, 
    3.928073e-11, 3.939353e-11, 3.963864e-11, 4.003344e-11, 3.988473e-11, 
    4.015796e-11, 4.021293e-11, 3.97979e-11, 4.005244e-11, 3.923857e-11, 
    3.936944e-11, 3.929149e-11, 3.900742e-11, 3.991892e-11, 3.944972e-11, 
    4.031843e-11, 4.006253e-11, 4.081178e-11, 4.043823e-11, 4.117367e-11, 
    4.149019e-11, 4.178932e-11, 4.214028e-11, 3.922064e-11, 3.912182e-11, 
    3.929885e-11, 3.954447e-11, 3.977312e-11, 4.007817e-11, 4.010945e-11, 
    4.016675e-11, 4.03154e-11, 4.044062e-11, 4.018486e-11, 4.047202e-11, 
    3.939981e-11, 3.995978e-11, 3.908443e-11, 3.934691e-11, 3.952991e-11, 
    3.944959e-11, 3.98677e-11, 3.996657e-11, 4.036973e-11, 4.016106e-11, 
    4.141193e-11, 4.085599e-11, 4.240858e-11, 4.197158e-11, 3.908732e-11, 
    3.922029e-11, 3.968494e-11, 3.94635e-11, 4.009857e-11, 4.025572e-11, 
    4.038371e-11, 4.054763e-11, 4.056535e-11, 4.066266e-11, 4.050325e-11, 
    4.065635e-11, 4.007877e-11, 4.033633e-11, 3.963165e-11, 3.980254e-11, 
    3.972387e-11, 3.963766e-11, 3.990402e-11, 4.018882e-11, 4.019493e-11, 
    4.028648e-11, 4.054504e-11, 4.010107e-11, 4.148392e-11, 4.062693e-11, 
    3.936556e-11, 3.962284e-11, 3.965968e-11, 3.955986e-11, 4.023993e-11, 
    3.99928e-11, 4.066029e-11, 4.047931e-11, 4.077605e-11, 4.062845e-11, 
    4.060674e-11, 4.041764e-11, 4.030012e-11, 4.000407e-11, 3.976404e-11, 
    3.957427e-11, 3.961835e-11, 3.982696e-11, 4.020627e-11, 4.056688e-11, 
    4.048774e-11, 4.07534e-11, 4.005225e-11, 4.034545e-11, 4.023198e-11, 
    4.05282e-11, 3.988077e-11, 4.043177e-11, 3.974055e-11, 3.98009e-11, 
    3.998789e-11, 4.036544e-11, 4.044924e-11, 4.05388e-11, 4.048352e-11, 
    4.021596e-11, 4.017222e-11, 3.998331e-11, 3.993122e-11, 3.978771e-11, 
    3.966909e-11, 3.977745e-11, 3.989141e-11, 4.021604e-11, 4.050979e-11, 
    4.083134e-11, 4.091025e-11, 4.128801e-11, 4.098033e-11, 4.148869e-11, 
    4.105623e-11, 4.180639e-11, 4.046384e-11, 4.104367e-11, 3.999642e-11, 
    4.010854e-11, 4.031177e-11, 4.077998e-11, 4.052686e-11, 4.082297e-11, 
    4.01705e-11, 3.983417e-11, 3.974741e-11, 3.958579e-11, 3.97511e-11, 
    3.973764e-11, 3.989614e-11, 3.984516e-11, 4.022683e-11, 4.002158e-11, 
    4.060613e-11, 4.082057e-11, 4.142944e-11, 4.180505e-11, 4.218928e-11, 
    4.23595e-11, 4.241138e-11, 4.243308e-11 ;

 F_NIT_vr =
  2.474889e-10, 2.485921e-10, 2.48377e-10, 2.492673e-10, 2.487732e-10, 
    2.493557e-10, 2.477113e-10, 2.486339e-10, 2.480445e-10, 2.475861e-10, 
    2.509944e-10, 2.493049e-10, 2.527535e-10, 2.516733e-10, 2.543881e-10, 
    2.525845e-10, 2.547519e-10, 2.543357e-10, 2.555885e-10, 2.55229e-10, 
    2.568318e-10, 2.557535e-10, 2.576638e-10, 2.565739e-10, 2.567438e-10, 
    2.557166e-10, 2.49647e-10, 2.507858e-10, 2.495789e-10, 2.497413e-10, 
    2.496682e-10, 2.487821e-10, 2.483357e-10, 2.474024e-10, 2.475714e-10, 
    2.482568e-10, 2.498124e-10, 2.492838e-10, 2.506158e-10, 2.505858e-10, 
    2.520702e-10, 2.514004e-10, 2.538994e-10, 2.531881e-10, 2.552437e-10, 
    2.547259e-10, 2.552188e-10, 2.550689e-10, 2.5522e-10, 2.544613e-10, 
    2.547857e-10, 2.541185e-10, 2.51529e-10, 2.522905e-10, 2.500191e-10, 
    2.486548e-10, 2.477505e-10, 2.471094e-10, 2.471994e-10, 2.473722e-10, 
    2.482603e-10, 2.490963e-10, 2.497339e-10, 2.501603e-10, 2.505807e-10, 
    2.518542e-10, 2.525294e-10, 2.540424e-10, 2.537693e-10, 2.542316e-10, 
    2.546741e-10, 2.554169e-10, 2.552945e-10, 2.556214e-10, 2.542182e-10, 
    2.551503e-10, 2.536114e-10, 2.54032e-10, 2.506964e-10, 2.494275e-10, 
    2.488875e-10, 2.484159e-10, 2.472688e-10, 2.480606e-10, 2.47748e-10, 
    2.484908e-10, 2.489629e-10, 2.48729e-10, 2.501717e-10, 2.4961e-10, 
    2.52569e-10, 2.512934e-10, 2.546229e-10, 2.538248e-10, 2.548134e-10, 
    2.543088e-10, 2.551729e-10, 2.543947e-10, 2.557429e-10, 2.560367e-10, 
    2.558353e-10, 2.566073e-10, 2.543498e-10, 2.552159e-10, 2.487239e-10, 
    2.487621e-10, 2.489393e-10, 2.481585e-10, 2.481107e-10, 2.473961e-10, 
    2.480313e-10, 2.483021e-10, 2.489897e-10, 2.493962e-10, 2.497829e-10, 
    2.506345e-10, 2.515857e-10, 2.529177e-10, 2.538761e-10, 2.545186e-10, 
    2.541243e-10, 2.544719e-10, 2.540827e-10, 2.539001e-10, 2.559258e-10, 
    2.547876e-10, 2.564955e-10, 2.56401e-10, 2.556271e-10, 2.564108e-10, 
    2.487883e-10, 2.485687e-10, 2.478076e-10, 2.484027e-10, 2.473178e-10, 
    2.479246e-10, 2.482732e-10, 2.496211e-10, 2.499175e-10, 2.501924e-10, 
    2.507355e-10, 2.514326e-10, 2.526573e-10, 2.537238e-10, 2.546988e-10, 
    2.54627e-10, 2.54652e-10, 2.548694e-10, 2.543296e-10, 2.549575e-10, 
    2.550624e-10, 2.547869e-10, 2.563875e-10, 2.559299e-10, 2.563979e-10, 
    2.560995e-10, 2.486397e-10, 2.490081e-10, 2.488084e-10, 2.491833e-10, 
    2.489185e-10, 2.500936e-10, 2.504458e-10, 2.520969e-10, 2.514188e-10, 
    2.524981e-10, 2.51528e-10, 2.516997e-10, 2.525319e-10, 2.515797e-10, 
    2.536639e-10, 2.522494e-10, 2.548775e-10, 2.53463e-10, 2.549656e-10, 
    2.546924e-10, 2.551439e-10, 2.555487e-10, 2.560577e-10, 2.569982e-10, 
    2.567798e-10, 2.575671e-10, 2.495582e-10, 2.500365e-10, 2.499945e-10, 
    2.504956e-10, 2.508662e-10, 2.51671e-10, 2.529624e-10, 2.524761e-10, 
    2.533682e-10, 2.535474e-10, 2.521912e-10, 2.530232e-10, 2.503545e-10, 
    2.507845e-10, 2.505283e-10, 2.495916e-10, 2.525855e-10, 2.510473e-10, 
    2.538887e-10, 2.53054e-10, 2.554902e-10, 2.542776e-10, 2.566597e-10, 
    2.576792e-10, 2.586402e-10, 2.597629e-10, 2.502979e-10, 2.49972e-10, 
    2.505547e-10, 2.513615e-10, 2.521108e-10, 2.531081e-10, 2.5321e-10, 
    2.533964e-10, 2.538806e-10, 2.54288e-10, 2.534546e-10, 2.543894e-10, 
    2.508835e-10, 2.527191e-10, 2.498452e-10, 2.507094e-10, 2.513103e-10, 
    2.510467e-10, 2.524172e-10, 2.5274e-10, 2.540541e-10, 2.533746e-10, 
    2.574265e-10, 2.556318e-10, 2.60619e-10, 2.59223e-10, 2.49858e-10, 
    2.502958e-10, 2.518216e-10, 2.510953e-10, 2.53174e-10, 2.536864e-10, 
    2.541027e-10, 2.546355e-10, 2.546926e-10, 2.550084e-10, 2.544904e-10, 
    2.549876e-10, 2.531073e-10, 2.53947e-10, 2.516444e-10, 2.522037e-10, 
    2.519462e-10, 2.516632e-10, 2.52535e-10, 2.534646e-10, 2.534845e-10, 
    2.537822e-10, 2.54622e-10, 2.531775e-10, 2.576565e-10, 2.548871e-10, 
    2.507735e-10, 2.516175e-10, 2.517383e-10, 2.514111e-10, 2.536343e-10, 
    2.52828e-10, 2.550008e-10, 2.544127e-10, 2.553755e-10, 2.548968e-10, 
    2.548258e-10, 2.542114e-10, 2.538283e-10, 2.528627e-10, 2.520771e-10, 
    2.514554e-10, 2.515994e-10, 2.522826e-10, 2.535208e-10, 2.546943e-10, 
    2.544367e-10, 2.552988e-10, 2.530176e-10, 2.539733e-10, 2.536031e-10, 
    2.545672e-10, 2.52462e-10, 2.542581e-10, 2.52003e-10, 2.522001e-10, 
    2.528112e-10, 2.54042e-10, 2.543145e-10, 2.546054e-10, 2.544254e-10, 
    2.535543e-10, 2.534115e-10, 2.527946e-10, 2.526239e-10, 2.521547e-10, 
    2.517656e-10, 2.521205e-10, 2.524927e-10, 2.535527e-10, 2.545082e-10, 
    2.55551e-10, 2.558065e-10, 2.570254e-10, 2.560321e-10, 2.576705e-10, 
    2.56276e-10, 2.586908e-10, 2.543621e-10, 2.562414e-10, 2.528392e-10, 
    2.532049e-10, 2.538668e-10, 2.553872e-10, 2.54566e-10, 2.555263e-10, 
    2.534058e-10, 2.523065e-10, 2.520225e-10, 2.514927e-10, 2.520341e-10, 
    2.5199e-10, 2.525085e-10, 2.523413e-10, 2.535872e-10, 2.529177e-10, 
    2.548203e-10, 2.555156e-10, 2.574813e-10, 2.586874e-10, 2.599174e-10, 
    2.604602e-10, 2.606255e-10, 2.606944e-10,
  1.257274e-10, 1.266888e-10, 1.265017e-10, 1.272786e-10, 1.268475e-10, 
    1.273565e-10, 1.259222e-10, 1.267269e-10, 1.26213e-10, 1.25814e-10, 
    1.287913e-10, 1.273133e-10, 1.303343e-10, 1.293865e-10, 1.317728e-10, 
    1.301866e-10, 1.320936e-10, 1.317272e-10, 1.328317e-10, 1.325149e-10, 
    1.33931e-10, 1.32978e-10, 1.346676e-10, 1.337033e-10, 1.338539e-10, 
    1.329465e-10, 1.276104e-10, 1.286069e-10, 1.275514e-10, 1.276933e-10, 
    1.276297e-10, 1.268563e-10, 1.264671e-10, 1.256542e-10, 1.258017e-10, 
    1.263989e-10, 1.277572e-10, 1.272956e-10, 1.284605e-10, 1.284342e-10, 
    1.297356e-10, 1.291482e-10, 1.313433e-10, 1.30718e-10, 1.325281e-10, 
    1.32072e-10, 1.325067e-10, 1.323748e-10, 1.325084e-10, 1.318396e-10, 
    1.32126e-10, 1.315382e-10, 1.292581e-10, 1.299265e-10, 1.279367e-10, 
    1.267456e-10, 1.259574e-10, 1.253991e-10, 1.25478e-10, 1.256283e-10, 
    1.264024e-10, 1.27132e-10, 1.276891e-10, 1.280623e-10, 1.284304e-10, 
    1.295465e-10, 1.301392e-10, 1.314698e-10, 1.312294e-10, 1.316368e-10, 
    1.320267e-10, 1.326819e-10, 1.32574e-10, 1.32863e-10, 1.316262e-10, 
    1.324476e-10, 1.310926e-10, 1.314626e-10, 1.285298e-10, 1.274201e-10, 
    1.26949e-10, 1.265376e-10, 1.255386e-10, 1.262282e-10, 1.259561e-10, 
    1.266038e-10, 1.270159e-10, 1.26812e-10, 1.280725e-10, 1.275818e-10, 
    1.301744e-10, 1.290552e-10, 1.319811e-10, 1.312788e-10, 1.321497e-10, 
    1.317051e-10, 1.324673e-10, 1.317812e-10, 1.329706e-10, 1.332301e-10, 
    1.330527e-10, 1.337347e-10, 1.317432e-10, 1.325066e-10, 1.268063e-10, 
    1.268395e-10, 1.269945e-10, 1.263139e-10, 1.262723e-10, 1.256501e-10, 
    1.262038e-10, 1.264397e-10, 1.270399e-10, 1.273952e-10, 1.277334e-10, 
    1.284783e-10, 1.29312e-10, 1.304814e-10, 1.313242e-10, 1.318903e-10, 
    1.315431e-10, 1.318496e-10, 1.31507e-10, 1.313466e-10, 1.331328e-10, 
    1.321286e-10, 1.336365e-10, 1.335529e-10, 1.328698e-10, 1.335623e-10, 
    1.268629e-10, 1.266716e-10, 1.260083e-10, 1.265273e-10, 1.255825e-10, 
    1.261109e-10, 1.264151e-10, 1.275919e-10, 1.278512e-10, 1.280916e-10, 
    1.285671e-10, 1.291782e-10, 1.302529e-10, 1.311908e-10, 1.320494e-10, 
    1.319864e-10, 1.320086e-10, 1.322006e-10, 1.317251e-10, 1.322787e-10, 
    1.323716e-10, 1.321286e-10, 1.335417e-10, 1.331374e-10, 1.335511e-10, 
    1.332879e-10, 1.267338e-10, 1.270557e-10, 1.268817e-10, 1.27209e-10, 
    1.269784e-10, 1.28005e-10, 1.283134e-10, 1.297607e-10, 1.291661e-10, 
    1.30113e-10, 1.292622e-10, 1.294128e-10, 1.301436e-10, 1.293082e-10, 
    1.311389e-10, 1.298964e-10, 1.32208e-10, 1.309631e-10, 1.322862e-10, 
    1.320457e-10, 1.32444e-10, 1.328011e-10, 1.33251e-10, 1.340824e-10, 
    1.338897e-10, 1.345862e-10, 1.275363e-10, 1.27955e-10, 1.279182e-10, 
    1.283569e-10, 1.286817e-10, 1.293868e-10, 1.305208e-10, 1.300939e-10, 
    1.308781e-10, 1.310357e-10, 1.298446e-10, 1.305753e-10, 1.282355e-10, 
    1.286123e-10, 1.28388e-10, 1.275693e-10, 1.301921e-10, 1.288434e-10, 
    1.313381e-10, 1.306044e-10, 1.327502e-10, 1.316813e-10, 1.337837e-10, 
    1.346859e-10, 1.355377e-10, 1.36535e-10, 1.281838e-10, 1.278991e-10, 
    1.284091e-10, 1.291159e-10, 1.297733e-10, 1.306491e-10, 1.307389e-10, 
    1.309033e-10, 1.313294e-10, 1.316881e-10, 1.309551e-10, 1.317781e-10, 
    1.286995e-10, 1.303095e-10, 1.277914e-10, 1.285475e-10, 1.290742e-10, 
    1.288432e-10, 1.300452e-10, 1.303291e-10, 1.314851e-10, 1.308871e-10, 
    1.344629e-10, 1.328764e-10, 1.372965e-10, 1.360558e-10, 1.277996e-10, 
    1.281829e-10, 1.295199e-10, 1.288831e-10, 1.307077e-10, 1.311583e-10, 
    1.315252e-10, 1.319944e-10, 1.320452e-10, 1.323236e-10, 1.318675e-10, 
    1.323057e-10, 1.30651e-10, 1.313895e-10, 1.293669e-10, 1.29858e-10, 
    1.296321e-10, 1.293843e-10, 1.301496e-10, 1.309666e-10, 1.309843e-10, 
    1.312467e-10, 1.319867e-10, 1.307152e-10, 1.346678e-10, 1.322212e-10, 
    1.286012e-10, 1.293413e-10, 1.294474e-10, 1.291604e-10, 1.311131e-10, 
    1.304042e-10, 1.323169e-10, 1.31799e-10, 1.32648e-10, 1.322258e-10, 
    1.321638e-10, 1.316224e-10, 1.312857e-10, 1.304367e-10, 1.297474e-10, 
    1.29202e-10, 1.293288e-10, 1.299282e-10, 1.310167e-10, 1.320497e-10, 
    1.318232e-10, 1.325834e-10, 1.305751e-10, 1.314157e-10, 1.310905e-10, 
    1.319391e-10, 1.300826e-10, 1.316623e-10, 1.296799e-10, 1.298533e-10, 
    1.303902e-10, 1.314727e-10, 1.317129e-10, 1.319692e-10, 1.318111e-10, 
    1.310444e-10, 1.309191e-10, 1.303772e-10, 1.302276e-10, 1.298155e-10, 
    1.294747e-10, 1.29786e-10, 1.301133e-10, 1.310448e-10, 1.318863e-10, 
    1.328062e-10, 1.330317e-10, 1.341097e-10, 1.332316e-10, 1.346814e-10, 
    1.33448e-10, 1.35586e-10, 1.317544e-10, 1.334122e-10, 1.304147e-10, 
    1.307364e-10, 1.313189e-10, 1.32659e-10, 1.319351e-10, 1.32782e-10, 
    1.309142e-10, 1.299488e-10, 1.296997e-10, 1.292351e-10, 1.297104e-10, 
    1.296717e-10, 1.30127e-10, 1.299806e-10, 1.310758e-10, 1.304871e-10, 
    1.321621e-10, 1.327753e-10, 1.345131e-10, 1.355824e-10, 1.366745e-10, 
    1.371575e-10, 1.373047e-10, 1.373662e-10,
  1.178461e-10, 1.188978e-10, 1.186931e-10, 1.195437e-10, 1.190715e-10, 
    1.196289e-10, 1.18059e-10, 1.189396e-10, 1.183772e-10, 1.179407e-10, 
    1.212018e-10, 1.195817e-10, 1.228952e-10, 1.218545e-10, 1.244763e-10, 
    1.227329e-10, 1.248291e-10, 1.24426e-10, 1.256414e-10, 1.252927e-10, 
    1.268525e-10, 1.258025e-10, 1.276645e-10, 1.266015e-10, 1.267675e-10, 
    1.257679e-10, 1.199071e-10, 1.209995e-10, 1.198424e-10, 1.199979e-10, 
    1.199282e-10, 1.190812e-10, 1.186553e-10, 1.177659e-10, 1.179272e-10, 
    1.185806e-10, 1.200679e-10, 1.195622e-10, 1.208387e-10, 1.208098e-10, 
    1.222376e-10, 1.21593e-10, 1.240038e-10, 1.233166e-10, 1.253072e-10, 
    1.248053e-10, 1.252836e-10, 1.251385e-10, 1.252855e-10, 1.245497e-10, 
    1.248647e-10, 1.242181e-10, 1.217135e-10, 1.224473e-10, 1.202645e-10, 
    1.189602e-10, 1.180976e-10, 1.17487e-10, 1.175733e-10, 1.177377e-10, 
    1.185844e-10, 1.193831e-10, 1.199932e-10, 1.204021e-10, 1.208056e-10, 
    1.220303e-10, 1.226809e-10, 1.241429e-10, 1.238787e-10, 1.243266e-10, 
    1.247554e-10, 1.254765e-10, 1.253577e-10, 1.256759e-10, 1.243149e-10, 
    1.252186e-10, 1.237282e-10, 1.24135e-10, 1.20915e-10, 1.196985e-10, 
    1.191828e-10, 1.187324e-10, 1.176396e-10, 1.183938e-10, 1.180962e-10, 
    1.188047e-10, 1.192559e-10, 1.190327e-10, 1.204133e-10, 1.198757e-10, 
    1.227195e-10, 1.21491e-10, 1.247053e-10, 1.239329e-10, 1.248908e-10, 
    1.244016e-10, 1.252403e-10, 1.244854e-10, 1.257944e-10, 1.260801e-10, 
    1.258848e-10, 1.26636e-10, 1.244436e-10, 1.252835e-10, 1.190264e-10, 
    1.190628e-10, 1.192324e-10, 1.184876e-10, 1.184421e-10, 1.177615e-10, 
    1.18367e-10, 1.186253e-10, 1.192821e-10, 1.196713e-10, 1.200418e-10, 
    1.208582e-10, 1.217727e-10, 1.230567e-10, 1.239829e-10, 1.246054e-10, 
    1.242235e-10, 1.245606e-10, 1.241838e-10, 1.240074e-10, 1.25973e-10, 
    1.248676e-10, 1.265278e-10, 1.264357e-10, 1.256834e-10, 1.264461e-10, 
    1.190884e-10, 1.18879e-10, 1.181533e-10, 1.187211e-10, 1.176875e-10, 
    1.182655e-10, 1.185984e-10, 1.198869e-10, 1.201709e-10, 1.204344e-10, 
    1.209556e-10, 1.216259e-10, 1.228057e-10, 1.238362e-10, 1.247804e-10, 
    1.247111e-10, 1.247355e-10, 1.249467e-10, 1.244237e-10, 1.250327e-10, 
    1.25135e-10, 1.248675e-10, 1.264234e-10, 1.259781e-10, 1.264338e-10, 
    1.261437e-10, 1.189471e-10, 1.192995e-10, 1.19109e-10, 1.194674e-10, 
    1.192148e-10, 1.203395e-10, 1.206776e-10, 1.222652e-10, 1.216127e-10, 
    1.226521e-10, 1.217181e-10, 1.218834e-10, 1.226859e-10, 1.217685e-10, 
    1.237792e-10, 1.224143e-10, 1.249549e-10, 1.235862e-10, 1.250409e-10, 
    1.247763e-10, 1.252146e-10, 1.256077e-10, 1.261031e-10, 1.270193e-10, 
    1.268069e-10, 1.275748e-10, 1.198259e-10, 1.202846e-10, 1.202443e-10, 
    1.207251e-10, 1.210812e-10, 1.218548e-10, 1.230999e-10, 1.226311e-10, 
    1.234925e-10, 1.236657e-10, 1.223573e-10, 1.231598e-10, 1.205921e-10, 
    1.210053e-10, 1.207592e-10, 1.19862e-10, 1.227389e-10, 1.212587e-10, 
    1.239982e-10, 1.231918e-10, 1.255517e-10, 1.243756e-10, 1.2669e-10, 
    1.276848e-10, 1.286245e-10, 1.297259e-10, 1.205353e-10, 1.202233e-10, 
    1.207824e-10, 1.215576e-10, 1.22279e-10, 1.232409e-10, 1.233395e-10, 
    1.235202e-10, 1.239886e-10, 1.24383e-10, 1.235772e-10, 1.24482e-10, 
    1.21101e-10, 1.228678e-10, 1.201053e-10, 1.209342e-10, 1.215119e-10, 
    1.212584e-10, 1.225776e-10, 1.228894e-10, 1.241598e-10, 1.235024e-10, 
    1.274389e-10, 1.256907e-10, 1.305675e-10, 1.291966e-10, 1.201143e-10, 
    1.205343e-10, 1.220009e-10, 1.213021e-10, 1.233053e-10, 1.238005e-10, 
    1.242038e-10, 1.2472e-10, 1.247758e-10, 1.250822e-10, 1.245803e-10, 
    1.250624e-10, 1.23243e-10, 1.240546e-10, 1.21833e-10, 1.22372e-10, 
    1.221239e-10, 1.21852e-10, 1.226921e-10, 1.235898e-10, 1.236092e-10, 
    1.238976e-10, 1.247118e-10, 1.233134e-10, 1.27665e-10, 1.249697e-10, 
    1.20993e-10, 1.218049e-10, 1.219213e-10, 1.216063e-10, 1.237508e-10, 
    1.229719e-10, 1.250747e-10, 1.245049e-10, 1.254392e-10, 1.249745e-10, 
    1.249062e-10, 1.243107e-10, 1.239406e-10, 1.230075e-10, 1.222506e-10, 
    1.21652e-10, 1.217911e-10, 1.224491e-10, 1.236449e-10, 1.247808e-10, 
    1.245316e-10, 1.253681e-10, 1.231596e-10, 1.240835e-10, 1.23726e-10, 
    1.246591e-10, 1.226186e-10, 1.243549e-10, 1.221764e-10, 1.223668e-10, 
    1.229565e-10, 1.241462e-10, 1.244103e-10, 1.246923e-10, 1.245182e-10, 
    1.236753e-10, 1.235375e-10, 1.229421e-10, 1.227779e-10, 1.223254e-10, 
    1.219512e-10, 1.22293e-10, 1.226524e-10, 1.236757e-10, 1.246011e-10, 
    1.256133e-10, 1.258616e-10, 1.270495e-10, 1.26082e-10, 1.276801e-10, 
    1.263206e-10, 1.286781e-10, 1.244561e-10, 1.26281e-10, 1.229833e-10, 
    1.233368e-10, 1.239771e-10, 1.254514e-10, 1.246547e-10, 1.255868e-10, 
    1.235321e-10, 1.224718e-10, 1.221982e-10, 1.216883e-10, 1.222099e-10, 
    1.221674e-10, 1.226674e-10, 1.225066e-10, 1.237098e-10, 1.230629e-10, 
    1.249045e-10, 1.255794e-10, 1.274941e-10, 1.28674e-10, 1.298799e-10, 
    1.304138e-10, 1.305765e-10, 1.306445e-10,
  1.203267e-10, 1.214804e-10, 1.212557e-10, 1.221892e-10, 1.21671e-10, 
    1.222829e-10, 1.205602e-10, 1.215262e-10, 1.209091e-10, 1.204304e-10, 
    1.24011e-10, 1.22231e-10, 1.258737e-10, 1.247286e-10, 1.276151e-10, 
    1.256952e-10, 1.28004e-10, 1.275596e-10, 1.288996e-10, 1.28515e-10, 
    1.302364e-10, 1.290773e-10, 1.311333e-10, 1.299592e-10, 1.301425e-10, 
    1.290392e-10, 1.225883e-10, 1.237887e-10, 1.225173e-10, 1.226881e-10, 
    1.226114e-10, 1.216816e-10, 1.212144e-10, 1.202388e-10, 1.204156e-10, 
    1.211323e-10, 1.227649e-10, 1.222095e-10, 1.236117e-10, 1.2358e-10, 
    1.2515e-10, 1.244409e-10, 1.270945e-10, 1.263375e-10, 1.285311e-10, 
    1.279777e-10, 1.285051e-10, 1.28345e-10, 1.285071e-10, 1.27696e-10, 
    1.280432e-10, 1.273306e-10, 1.245735e-10, 1.253807e-10, 1.229809e-10, 
    1.215489e-10, 1.206025e-10, 1.19933e-10, 1.200276e-10, 1.202078e-10, 
    1.211365e-10, 1.220129e-10, 1.226829e-10, 1.23132e-10, 1.235754e-10, 
    1.24922e-10, 1.256378e-10, 1.272478e-10, 1.269565e-10, 1.274502e-10, 
    1.279227e-10, 1.287178e-10, 1.285868e-10, 1.289377e-10, 1.274372e-10, 
    1.284335e-10, 1.267908e-10, 1.27239e-10, 1.236959e-10, 1.223593e-10, 
    1.217932e-10, 1.212988e-10, 1.201003e-10, 1.209273e-10, 1.20601e-10, 
    1.213782e-10, 1.218733e-10, 1.216283e-10, 1.231443e-10, 1.225538e-10, 
    1.256803e-10, 1.243289e-10, 1.278675e-10, 1.270163e-10, 1.28072e-10, 
    1.275328e-10, 1.284573e-10, 1.276251e-10, 1.290685e-10, 1.293838e-10, 
    1.291683e-10, 1.299972e-10, 1.27579e-10, 1.28505e-10, 1.216214e-10, 
    1.216614e-10, 1.218475e-10, 1.210302e-10, 1.209803e-10, 1.202339e-10, 
    1.20898e-10, 1.211813e-10, 1.21902e-10, 1.223293e-10, 1.227362e-10, 
    1.236332e-10, 1.246387e-10, 1.260515e-10, 1.270714e-10, 1.277573e-10, 
    1.273365e-10, 1.27708e-10, 1.272927e-10, 1.270984e-10, 1.292656e-10, 
    1.280464e-10, 1.298778e-10, 1.297762e-10, 1.289461e-10, 1.297876e-10, 
    1.216894e-10, 1.214597e-10, 1.206635e-10, 1.212863e-10, 1.201528e-10, 
    1.207866e-10, 1.211518e-10, 1.225661e-10, 1.22878e-10, 1.231674e-10, 
    1.237402e-10, 1.244771e-10, 1.257751e-10, 1.269099e-10, 1.279502e-10, 
    1.278738e-10, 1.279007e-10, 1.281336e-10, 1.275571e-10, 1.282284e-10, 
    1.283412e-10, 1.280463e-10, 1.297626e-10, 1.292711e-10, 1.29774e-10, 
    1.294539e-10, 1.215343e-10, 1.219212e-10, 1.217121e-10, 1.221055e-10, 
    1.218282e-10, 1.230633e-10, 1.234348e-10, 1.251804e-10, 1.244626e-10, 
    1.256061e-10, 1.245785e-10, 1.247603e-10, 1.256434e-10, 1.24634e-10, 
    1.268471e-10, 1.253445e-10, 1.281427e-10, 1.266346e-10, 1.282375e-10, 
    1.279457e-10, 1.28429e-10, 1.288626e-10, 1.294091e-10, 1.304205e-10, 
    1.30186e-10, 1.31034e-10, 1.224991e-10, 1.230029e-10, 1.229586e-10, 
    1.234869e-10, 1.238783e-10, 1.247289e-10, 1.26099e-10, 1.255829e-10, 
    1.265312e-10, 1.267219e-10, 1.252816e-10, 1.26165e-10, 1.233408e-10, 
    1.237949e-10, 1.235244e-10, 1.225388e-10, 1.257017e-10, 1.240735e-10, 
    1.270883e-10, 1.262001e-10, 1.288007e-10, 1.275041e-10, 1.30057e-10, 
    1.311558e-10, 1.321942e-10, 1.334127e-10, 1.232784e-10, 1.229356e-10, 
    1.235498e-10, 1.244021e-10, 1.251955e-10, 1.262542e-10, 1.263628e-10, 
    1.265617e-10, 1.270776e-10, 1.275122e-10, 1.266246e-10, 1.276213e-10, 
    1.239003e-10, 1.258435e-10, 1.22806e-10, 1.237168e-10, 1.243518e-10, 
    1.240731e-10, 1.25524e-10, 1.258672e-10, 1.272664e-10, 1.265421e-10, 
    1.308841e-10, 1.289542e-10, 1.343442e-10, 1.328271e-10, 1.228159e-10, 
    1.232772e-10, 1.248896e-10, 1.241212e-10, 1.263251e-10, 1.268705e-10, 
    1.273147e-10, 1.278837e-10, 1.279452e-10, 1.28283e-10, 1.277297e-10, 
    1.282611e-10, 1.262565e-10, 1.271504e-10, 1.247048e-10, 1.252979e-10, 
    1.250249e-10, 1.247257e-10, 1.256501e-10, 1.266385e-10, 1.266597e-10, 
    1.269775e-10, 1.27875e-10, 1.263341e-10, 1.311341e-10, 1.281593e-10, 
    1.237813e-10, 1.246741e-10, 1.24802e-10, 1.244556e-10, 1.268157e-10, 
    1.25958e-10, 1.282747e-10, 1.276466e-10, 1.286766e-10, 1.281643e-10, 
    1.28089e-10, 1.274326e-10, 1.270248e-10, 1.259973e-10, 1.251643e-10, 
    1.245058e-10, 1.246588e-10, 1.253827e-10, 1.266991e-10, 1.279507e-10, 
    1.276761e-10, 1.285982e-10, 1.261646e-10, 1.271823e-10, 1.267885e-10, 
    1.278166e-10, 1.255692e-10, 1.274816e-10, 1.250826e-10, 1.252921e-10, 
    1.25941e-10, 1.272514e-10, 1.275423e-10, 1.278531e-10, 1.276613e-10, 
    1.267327e-10, 1.265808e-10, 1.259252e-10, 1.257445e-10, 1.252465e-10, 
    1.248349e-10, 1.252109e-10, 1.256064e-10, 1.26733e-10, 1.277526e-10, 
    1.288687e-10, 1.291427e-10, 1.304541e-10, 1.29386e-10, 1.311508e-10, 
    1.296495e-10, 1.322537e-10, 1.275929e-10, 1.296056e-10, 1.259706e-10, 
    1.263598e-10, 1.270652e-10, 1.286903e-10, 1.278117e-10, 1.288395e-10, 
    1.265749e-10, 1.254077e-10, 1.251066e-10, 1.245458e-10, 1.251194e-10, 
    1.250727e-10, 1.256228e-10, 1.254459e-10, 1.267705e-10, 1.260582e-10, 
    1.280871e-10, 1.288314e-10, 1.30945e-10, 1.32249e-10, 1.33583e-10, 
    1.34174e-10, 1.343541e-10, 1.344295e-10,
  1.309803e-10, 1.322135e-10, 1.319732e-10, 1.329718e-10, 1.324173e-10, 
    1.33072e-10, 1.312297e-10, 1.322626e-10, 1.316027e-10, 1.31091e-10, 
    1.349223e-10, 1.330165e-10, 1.369187e-10, 1.356909e-10, 1.387876e-10, 
    1.367273e-10, 1.392053e-10, 1.38728e-10, 1.401676e-10, 1.397542e-10, 
    1.416053e-10, 1.403586e-10, 1.425705e-10, 1.41307e-10, 1.415042e-10, 
    1.403176e-10, 1.333987e-10, 1.346842e-10, 1.333228e-10, 1.335056e-10, 
    1.334235e-10, 1.324288e-10, 1.319291e-10, 1.308862e-10, 1.310752e-10, 
    1.318413e-10, 1.335878e-10, 1.329934e-10, 1.344943e-10, 1.344603e-10, 
    1.361426e-10, 1.353826e-10, 1.382286e-10, 1.374161e-10, 1.397715e-10, 
    1.391769e-10, 1.397435e-10, 1.395716e-10, 1.397458e-10, 1.388744e-10, 
    1.392473e-10, 1.38482e-10, 1.355247e-10, 1.3639e-10, 1.33819e-10, 
    1.322869e-10, 1.312749e-10, 1.305596e-10, 1.306606e-10, 1.308532e-10, 
    1.318459e-10, 1.327831e-10, 1.334999e-10, 1.339807e-10, 1.344554e-10, 
    1.358984e-10, 1.366658e-10, 1.383932e-10, 1.380805e-10, 1.386105e-10, 
    1.391179e-10, 1.399722e-10, 1.398314e-10, 1.402086e-10, 1.385965e-10, 
    1.396666e-10, 1.379026e-10, 1.383837e-10, 1.345848e-10, 1.331536e-10, 
    1.325481e-10, 1.320194e-10, 1.307383e-10, 1.316222e-10, 1.312733e-10, 
    1.321042e-10, 1.326337e-10, 1.323717e-10, 1.339939e-10, 1.333618e-10, 
    1.367113e-10, 1.352626e-10, 1.390586e-10, 1.381446e-10, 1.392782e-10, 
    1.386991e-10, 1.396923e-10, 1.387982e-10, 1.403491e-10, 1.406881e-10, 
    1.404564e-10, 1.413478e-10, 1.387488e-10, 1.397435e-10, 1.323644e-10, 
    1.324071e-10, 1.326062e-10, 1.317322e-10, 1.316788e-10, 1.308811e-10, 
    1.315908e-10, 1.318937e-10, 1.326645e-10, 1.331216e-10, 1.335571e-10, 
    1.345173e-10, 1.355946e-10, 1.371094e-10, 1.382038e-10, 1.389402e-10, 
    1.384884e-10, 1.388872e-10, 1.384414e-10, 1.382327e-10, 1.40561e-10, 
    1.392508e-10, 1.412194e-10, 1.411101e-10, 1.402176e-10, 1.411224e-10, 
    1.324371e-10, 1.321913e-10, 1.313402e-10, 1.32006e-10, 1.307944e-10, 
    1.314718e-10, 1.318622e-10, 1.33375e-10, 1.337088e-10, 1.340187e-10, 
    1.34632e-10, 1.354214e-10, 1.368129e-10, 1.380304e-10, 1.391474e-10, 
    1.390654e-10, 1.390943e-10, 1.393445e-10, 1.387252e-10, 1.394463e-10, 
    1.395675e-10, 1.392507e-10, 1.410954e-10, 1.405669e-10, 1.411077e-10, 
    1.407635e-10, 1.322712e-10, 1.32685e-10, 1.324613e-10, 1.328821e-10, 
    1.325856e-10, 1.339072e-10, 1.34305e-10, 1.361753e-10, 1.354059e-10, 
    1.366317e-10, 1.355301e-10, 1.357249e-10, 1.366718e-10, 1.355895e-10, 
    1.379631e-10, 1.363513e-10, 1.393542e-10, 1.377351e-10, 1.39456e-10, 
    1.391426e-10, 1.396618e-10, 1.401278e-10, 1.407153e-10, 1.418033e-10, 
    1.415509e-10, 1.424636e-10, 1.333033e-10, 1.338426e-10, 1.33795e-10, 
    1.343607e-10, 1.347799e-10, 1.356912e-10, 1.371603e-10, 1.366067e-10, 
    1.376239e-10, 1.378287e-10, 1.362837e-10, 1.372311e-10, 1.342042e-10, 
    1.346906e-10, 1.344009e-10, 1.333458e-10, 1.367342e-10, 1.349891e-10, 
    1.382219e-10, 1.372688e-10, 1.400613e-10, 1.386684e-10, 1.414121e-10, 
    1.425948e-10, 1.437131e-10, 1.450267e-10, 1.341375e-10, 1.337704e-10, 
    1.34428e-10, 1.353411e-10, 1.361914e-10, 1.373268e-10, 1.374433e-10, 
    1.376567e-10, 1.382104e-10, 1.38677e-10, 1.377243e-10, 1.387941e-10, 
    1.348036e-10, 1.368863e-10, 1.336318e-10, 1.34607e-10, 1.352872e-10, 
    1.349885e-10, 1.365435e-10, 1.369116e-10, 1.384132e-10, 1.376357e-10, 
    1.423024e-10, 1.402264e-10, 1.460316e-10, 1.443952e-10, 1.336423e-10, 
    1.341362e-10, 1.358635e-10, 1.3504e-10, 1.374028e-10, 1.379881e-10, 
    1.38465e-10, 1.39076e-10, 1.391421e-10, 1.395049e-10, 1.389106e-10, 
    1.394814e-10, 1.373292e-10, 1.382886e-10, 1.356654e-10, 1.363011e-10, 
    1.360084e-10, 1.356878e-10, 1.366788e-10, 1.377392e-10, 1.377619e-10, 
    1.38103e-10, 1.39067e-10, 1.374124e-10, 1.425717e-10, 1.393723e-10, 
    1.34676e-10, 1.356326e-10, 1.357695e-10, 1.353983e-10, 1.379293e-10, 
    1.370091e-10, 1.394961e-10, 1.388213e-10, 1.399279e-10, 1.393774e-10, 
    1.392965e-10, 1.385915e-10, 1.381537e-10, 1.370512e-10, 1.36158e-10, 
    1.354521e-10, 1.35616e-10, 1.363921e-10, 1.378043e-10, 1.39148e-10, 
    1.38853e-10, 1.398436e-10, 1.372307e-10, 1.383228e-10, 1.379001e-10, 
    1.390039e-10, 1.365921e-10, 1.386444e-10, 1.360703e-10, 1.362949e-10, 
    1.369908e-10, 1.383971e-10, 1.387093e-10, 1.390432e-10, 1.388371e-10, 
    1.378402e-10, 1.376773e-10, 1.369739e-10, 1.367801e-10, 1.36246e-10, 
    1.358048e-10, 1.362079e-10, 1.36632e-10, 1.378406e-10, 1.389352e-10, 
    1.401344e-10, 1.404288e-10, 1.418395e-10, 1.406906e-10, 1.425896e-10, 
    1.409742e-10, 1.437775e-10, 1.387639e-10, 1.409268e-10, 1.370226e-10, 
    1.3744e-10, 1.381971e-10, 1.399427e-10, 1.389987e-10, 1.401031e-10, 
    1.376709e-10, 1.364189e-10, 1.360961e-10, 1.354949e-10, 1.361098e-10, 
    1.360597e-10, 1.366495e-10, 1.364598e-10, 1.378808e-10, 1.371165e-10, 
    1.392945e-10, 1.400943e-10, 1.423678e-10, 1.437722e-10, 1.452102e-10, 
    1.458479e-10, 1.460422e-10, 1.461236e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24572.98, 24593.23, 24589.26, 24605.83, 24596.6, 24607.5, 24577.05, 
    24594.04, 24583.16, 24574.78, 24638.73, 24606.57, 24673.14, 24651.87, 
    24705.73, 24669.8, 24713.11, 24704.67, 24730.29, 24722.88, 24756.45, 
    24733.73, 24774.34, 24750.97, 24754.59, 24732.99, 24612.97, 24634.68, 
    24611.7, 24614.77, 24613.39, 24596.79, 24588.53, 24571.45, 24574.53, 
    24587.08, 24616.15, 24606.19, 24631.46, 24630.88, 24659.66, 24646.58, 
    24695.91, 24681.79, 24723.19, 24712.6, 24722.69, 24719.62, 24722.73, 
    24707.25, 24713.85, 24700.35, 24649.02, 24663.94, 24620.05, 24594.44, 
    24577.79, 24566.13, 24567.77, 24570.91, 24587.16, 24602.68, 24614.67, 
    24622.78, 24630.8, 24655.45, 24668.73, 24698.79, 24693.32, 24702.61, 
    24711.56, 24726.78, 24724.26, 24731.03, 24702.36, 24721.32, 24690.22, 
    24698.63, 24633, 24608.87, 24598.77, 24590.02, 24569.04, 24583.48, 
    24577.76, 24591.42, 24600.19, 24595.84, 24623, 24612.36, 24669.53, 
    24644.53, 24710.51, 24694.44, 24714.4, 24704.16, 24721.77, 24705.91, 
    24733.56, 24739.7, 24735.5, 24751.72, 24705.04, 24722.69, 24595.72, 
    24596.43, 24599.74, 24585.29, 24584.41, 24571.36, 24582.96, 24587.95, 
    24600.71, 24608.33, 24615.63, 24631.85, 24650.22, 24676.47, 24695.48, 
    24708.41, 24700.46, 24707.48, 24699.64, 24695.98, 24737.39, 24713.91, 
    24749.37, 24747.37, 24731.19, 24747.6, 24596.93, 24592.86, 24578.86, 
    24589.8, 24569.95, 24581.01, 24587.43, 24612.58, 24618.19, 24623.42, 
    24633.79, 24647.25, 24671.29, 24692.45, 24712.08, 24710.63, 24711.14, 
    24715.58, 24704.62, 24717.39, 24719.55, 24713.91, 24747.1, 24737.5, 
    24747.33, 24741.06, 24594.18, 24601.05, 24597.33, 24604.33, 24599.39, 
    24621.54, 24628.26, 24660.23, 24646.98, 24668.14, 24649.11, 24652.46, 
    24668.84, 24650.13, 24691.28, 24663.27, 24715.75, 24687.32, 24717.56, 
    24711.99, 24721.23, 24729.58, 24740.19, 24760.09, 24755.45, 24772.34, 
    24611.37, 24620.45, 24619.64, 24629.2, 24636.3, 24651.88, 24677.36, 
    24667.7, 24685.39, 24688.94, 24662.1, 24678.6, 24626.56, 24634.79, 
    24629.88, 24612.09, 24669.92, 24639.86, 24695.79, 24679.25, 24728.38, 
    24703.62, 24752.9, 24774.79, 24795.88, 24820.93, 24625.43, 24619.23, 
    24630.34, 24645.87, 24660.51, 24680.25, 24682.26, 24685.96, 24695.59, 
    24703.78, 24687.13, 24705.84, 24636.71, 24672.57, 24616.89, 24633.37, 
    24644.95, 24639.85, 24666.61, 24673.01, 24699.14, 24685.59, 24769.34, 
    24731.35, 24840.21, 24808.91, 24617.07, 24625.41, 24654.85, 24640.73, 
    24681.56, 24691.71, 24700.05, 24710.82, 24711.98, 24718.43, 24707.89, 
    24718.01, 24680.29, 24696.96, 24651.43, 24662.4, 24657.34, 24651.82, 
    24668.96, 24687.39, 24687.78, 24693.72, 24710.66, 24681.73, 24774.37, 
    24716.08, 24634.54, 24650.87, 24653.23, 24646.85, 24690.69, 24674.72, 
    24718.27, 24706.32, 24725.99, 24716.16, 24714.72, 24702.27, 24694.6, 
    24675.45, 24659.93, 24647.77, 24650.59, 24663.98, 24688.52, 24712.09, 
    24706.88, 24724.48, 24678.59, 24697.56, 24690.18, 24709.54, 24667.45, 
    24703.21, 24658.41, 24662.29, 24674.4, 24698.86, 24704.34, 24710.24, 
    24706.6, 24689.14, 24686.31, 24674.1, 24670.72, 24661.45, 24653.83, 
    24660.79, 24668.14, 24689.15, 24708.33, 24729.7, 24735, 24760.77, 
    24739.74, 24774.7, 24744.9, 24797.11, 24705.31, 24744.03, 24674.95, 
    24682.2, 24695.36, 24726.26, 24709.45, 24729.13, 24686.2, 24664.45, 
    24658.86, 24648.51, 24659.1, 24658.23, 24668.45, 24665.15, 24689.85, 
    24676.59, 24714.69, 24728.98, 24770.56, 24797, 24824.43, 24836.67, 
    24840.42, 24841.99 ;

 GC_ICE1 =
  17681.28, 17713.7, 17707.35, 17733.88, 17719.11, 17736.56, 17687.8, 
    17715.01, 17697.59, 17684.17, 17786.54, 17735.07, 17841.57, 17807.56, 
    17893.56, 17836.23, 17905.34, 17891.88, 17932.75, 17920.92, 17974.46, 
    17938.23, 18002.98, 17965.72, 17971.49, 17937.05, 17745.32, 17780.06, 
    17743.28, 17748.2, 17745.99, 17719.41, 17706.19, 17678.83, 17683.76, 
    17703.87, 17750.41, 17734.46, 17774.91, 17773.99, 17820.02, 17799.1, 
    17877.91, 17855.38, 17921.42, 17904.54, 17920.62, 17915.72, 17920.68, 
    17896, 17906.53, 17884.99, 17802.99, 17826.86, 17756.65, 17715.65, 
    17688.99, 17670.31, 17672.95, 17677.96, 17703.99, 17728.84, 17748.04, 
    17761.02, 17773.86, 17813.28, 17834.52, 17882.51, 17873.78, 17888.59, 
    17902.87, 17927.15, 17923.12, 17933.92, 17888.19, 17918.43, 17868.84, 
    17882.24, 17777.37, 17738.74, 17722.59, 17708.57, 17674.97, 17698.1, 
    17688.95, 17710.81, 17724.86, 17717.89, 17761.38, 17744.33, 17835.79, 
    17795.81, 17901.19, 17875.57, 17907.4, 17891.07, 17919.16, 17893.86, 
    17937.96, 17947.74, 17941.05, 17966.91, 17892.47, 17920.62, 17717.7, 
    17718.83, 17724.13, 17700.99, 17699.59, 17678.69, 17697.27, 17705.25, 
    17725.68, 17737.89, 17749.58, 17775.53, 17804.91, 17846.89, 17877.22, 
    17897.85, 17885.17, 17896.36, 17883.85, 17878.02, 17944.07, 17906.63, 
    17963.16, 17959.98, 17934.18, 17960.34, 17719.63, 17713.11, 17690.7, 
    17708.21, 17676.43, 17694.15, 17704.42, 17744.69, 17753.67, 17762.05, 
    17778.64, 17800.16, 17838.61, 17872.39, 17903.7, 17901.38, 17902.2, 
    17909.28, 17891.81, 17912.16, 17915.61, 17906.62, 17959.55, 17944.24, 
    17959.91, 17949.92, 17715.23, 17726.22, 17720.27, 17731.48, 17723.58, 
    17759.04, 17769.79, 17820.93, 17799.73, 17833.57, 17803.14, 17808.49, 
    17834.69, 17804.77, 17870.53, 17825.79, 17909.55, 17864.2, 17912.44, 
    17903.56, 17918.29, 17931.61, 17948.53, 17980.27, 17972.86, 17999.79, 
    17742.76, 17757.29, 17756, 17771.29, 17782.66, 17807.57, 17848.32, 
    17832.87, 17861.12, 17866.79, 17823.92, 17850.29, 17767.07, 17780.23, 
    17772.38, 17743.9, 17836.42, 17788.35, 17877.72, 17851.33, 17929.7, 
    17890.21, 17968.79, 18003.71, 18037.31, 18077.19, 17765.27, 17755.33, 
    17773.12, 17797.96, 17821.37, 17852.92, 17856.13, 17862.03, 17877.4, 
    17890.46, 17863.9, 17893.74, 17783.31, 17840.66, 17751.6, 17777.96, 
    17796.49, 17788.33, 17831.12, 17841.36, 17883.06, 17861.45, 17995.01, 
    17934.44, 18107.83, 18058.07, 17751.88, 17765.23, 17812.31, 17789.74, 
    17855.02, 17871.21, 17884.51, 17901.69, 17903.55, 17913.83, 17897.02, 
    17913.16, 17852.99, 17879.58, 17806.86, 17824.4, 17816.31, 17807.47, 
    17834.88, 17864.31, 17864.94, 17874.41, 17901.44, 17855.28, 18003.02, 
    17910.07, 17779.83, 17805.96, 17809.72, 17799.53, 17869.58, 17844.09, 
    17913.58, 17894.51, 17925.88, 17910.21, 17907.92, 17888.06, 17875.82, 
    17845.26, 17820.44, 17801, 17805.5, 17826.92, 17866.12, 17903.72, 
    17895.4, 17923.47, 17850.28, 17880.54, 17868.77, 17899.65, 17832.47, 
    17889.55, 17818.02, 17824.23, 17843.58, 17882.62, 17891.36, 17900.76, 
    17894.95, 17867.11, 17862.6, 17843.1, 17837.7, 17822.87, 17810.69, 
    17821.82, 17833.58, 17867.12, 17897.71, 17931.8, 17940.26, 17981.34, 
    17947.81, 18003.56, 17956.04, 18039.27, 17892.9, 17954.66, 17844.46, 
    17856.04, 17877.04, 17926.31, 17899.5, 17930.9, 17862.42, 17827.66, 
    17818.73, 17802.18, 17819.11, 17817.73, 17834.06, 17828.79, 17868.24, 
    17847.09, 17907.86, 17930.65, 17996.95, 18039.1, 18082.76, 18102.2, 
    18108.15, 18110.65 ;

 GC_LIQ1 =
  5232.713, 5234.742, 5234.345, 5236.006, 5235.081, 5236.174, 5233.122, 
    5234.824, 5233.733, 5232.895, 5239.315, 5236.081, 5242.794, 5240.642, 
    5246.144, 5242.456, 5246.906, 5246.036, 5248.679, 5247.914, 5251.38, 
    5249.034, 5253.229, 5250.814, 5251.188, 5248.958, 5236.723, 5238.906, 
    5236.595, 5236.903, 5236.764, 5235.1, 5234.272, 5232.56, 5232.869, 
    5234.127, 5237.042, 5236.042, 5238.581, 5238.523, 5241.43, 5240.108, 
    5245.132, 5243.676, 5247.946, 5246.854, 5247.894, 5247.577, 5247.898, 
    5246.302, 5246.982, 5245.589, 5240.354, 5241.863, 5237.432, 5234.864, 
    5233.195, 5232.028, 5232.193, 5232.506, 5234.134, 5235.69, 5236.893, 
    5237.706, 5238.514, 5241.004, 5242.348, 5245.429, 5244.865, 5245.822, 
    5246.746, 5248.317, 5248.056, 5248.755, 5245.797, 5247.752, 5244.546, 
    5245.412, 5238.736, 5236.311, 5235.299, 5234.421, 5232.319, 5233.766, 
    5233.193, 5234.561, 5235.441, 5235.005, 5237.729, 5236.661, 5242.428, 
    5239.9, 5246.637, 5244.981, 5247.039, 5245.983, 5247.8, 5246.163, 
    5249.017, 5249.65, 5249.217, 5250.892, 5246.073, 5247.894, 5234.993, 
    5235.063, 5235.395, 5233.947, 5233.859, 5232.552, 5233.714, 5234.213, 
    5235.492, 5236.257, 5236.989, 5238.62, 5240.475, 5243.131, 5245.087, 
    5246.421, 5245.601, 5246.325, 5245.516, 5245.139, 5249.412, 5246.989, 
    5250.649, 5250.442, 5248.772, 5250.466, 5235.113, 5234.706, 5233.302, 
    5234.399, 5232.41, 5233.519, 5234.161, 5236.683, 5237.246, 5237.771, 
    5238.816, 5240.175, 5242.607, 5244.775, 5246.799, 5246.65, 5246.703, 
    5247.16, 5246.03, 5247.347, 5247.57, 5246.988, 5250.415, 5249.423, 
    5250.438, 5249.791, 5234.838, 5235.526, 5235.154, 5235.855, 5235.361, 
    5237.582, 5238.258, 5241.487, 5240.148, 5242.288, 5240.363, 5240.702, 
    5242.358, 5240.466, 5244.655, 5241.795, 5247.178, 5244.246, 5247.365, 
    5246.791, 5247.744, 5248.605, 5249.701, 5251.757, 5251.277, 5253.023, 
    5236.562, 5237.472, 5237.392, 5238.353, 5239.07, 5240.643, 5243.222, 
    5242.244, 5244.047, 5244.414, 5241.676, 5243.348, 5238.086, 5238.917, 
    5238.421, 5236.633, 5242.468, 5239.429, 5245.12, 5243.415, 5248.482, 
    5245.927, 5251.014, 5253.277, 5255.458, 5258.077, 5237.973, 5237.35, 
    5238.468, 5240.036, 5241.515, 5243.518, 5243.725, 5244.105, 5245.099, 
    5245.943, 5244.227, 5246.156, 5239.111, 5242.737, 5237.116, 5238.774, 
    5239.943, 5239.428, 5242.132, 5242.781, 5245.465, 5244.068, 5252.713, 
    5248.789, 5260.122, 5256.81, 5237.133, 5237.97, 5240.942, 5239.517, 
    5243.653, 5244.699, 5245.559, 5246.669, 5246.79, 5247.455, 5246.368, 
    5247.412, 5243.522, 5245.24, 5240.598, 5241.707, 5241.195, 5240.637, 
    5242.371, 5244.253, 5244.294, 5244.906, 5246.653, 5243.67, 5253.232, 
    5247.212, 5238.892, 5240.542, 5240.779, 5240.135, 5244.594, 5242.954, 
    5247.438, 5246.205, 5248.235, 5247.221, 5247.072, 5245.788, 5244.997, 
    5243.028, 5241.457, 5240.228, 5240.512, 5241.867, 5244.37, 5246.801, 
    5246.263, 5248.079, 5243.347, 5245.302, 5244.542, 5246.538, 5242.218, 
    5245.884, 5241.303, 5241.696, 5242.921, 5245.436, 5246.001, 5246.609, 
    5246.234, 5244.434, 5244.143, 5242.892, 5242.549, 5241.61, 5240.84, 
    5241.543, 5242.288, 5244.435, 5246.413, 5248.618, 5249.165, 5251.827, 
    5249.655, 5253.267, 5250.188, 5255.586, 5246.101, 5250.098, 5242.978, 
    5243.719, 5245.075, 5248.262, 5246.528, 5248.56, 5244.131, 5241.914, 
    5241.348, 5240.302, 5241.372, 5241.285, 5242.319, 5241.985, 5244.507, 
    5243.144, 5247.069, 5248.543, 5252.839, 5255.575, 5258.447, 5259.745, 
    5260.144, 5260.311 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.726522e-09, 8.765269e-09, 8.757737e-09, 8.788989e-09, 8.771654e-09, 
    8.792117e-09, 8.734378e-09, 8.766806e-09, 8.746104e-09, 8.730011e-09, 
    8.849647e-09, 8.790384e-09, 8.911227e-09, 8.873422e-09, 8.968403e-09, 
    8.905344e-09, 8.981121e-09, 8.966587e-09, 9.010338e-09, 8.997804e-09, 
    9.053768e-09, 9.016125e-09, 9.082785e-09, 9.044779e-09, 9.050723e-09, 
    9.014882e-09, 8.802312e-09, 8.842268e-09, 8.799944e-09, 8.805642e-09, 
    8.803085e-09, 8.772011e-09, 8.75635e-09, 8.723562e-09, 8.729515e-09, 
    8.753598e-09, 8.808204e-09, 8.789668e-09, 8.836389e-09, 8.835334e-09, 
    8.887355e-09, 8.863899e-09, 8.951348e-09, 8.926492e-09, 8.998327e-09, 
    8.98026e-09, 8.997478e-09, 8.992258e-09, 8.997546e-09, 8.971049e-09, 
    8.982401e-09, 8.959087e-09, 8.868291e-09, 8.894971e-09, 8.815403e-09, 
    8.767565e-09, 8.7358e-09, 8.713259e-09, 8.716445e-09, 8.72252e-09, 
    8.753739e-09, 8.783095e-09, 8.805468e-09, 8.820435e-09, 8.835182e-09, 
    8.87982e-09, 8.903454e-09, 8.956373e-09, 8.946825e-09, 8.963003e-09, 
    8.978462e-09, 9.004416e-09, 9.000145e-09, 9.011579e-09, 8.962578e-09, 
    8.995142e-09, 8.941385e-09, 8.956087e-09, 8.839184e-09, 8.794669e-09, 
    8.775743e-09, 8.759184e-09, 8.718896e-09, 8.746716e-09, 8.735749e-09, 
    8.761844e-09, 8.778426e-09, 8.770225e-09, 8.820844e-09, 8.801163e-09, 
    8.904855e-09, 8.860187e-09, 8.976659e-09, 8.948785e-09, 8.98334e-09, 
    8.965708e-09, 8.995921e-09, 8.96873e-09, 9.015835e-09, 9.026093e-09, 
    9.019083e-09, 9.046013e-09, 8.967222e-09, 8.997477e-09, 8.769995e-09, 
    8.771332e-09, 8.777564e-09, 8.750172e-09, 8.748496e-09, 8.723398e-09, 
    8.745731e-09, 8.755241e-09, 8.779388e-09, 8.79367e-09, 8.807247e-09, 
    8.837102e-09, 8.870447e-09, 8.917082e-09, 8.950591e-09, 8.973054e-09, 
    8.959281e-09, 8.971441e-09, 8.957847e-09, 8.951476e-09, 9.022249e-09, 
    8.982507e-09, 9.042139e-09, 9.03884e-09, 9.011851e-09, 9.039211e-09, 
    8.772272e-09, 8.764575e-09, 8.737852e-09, 8.758765e-09, 8.720665e-09, 
    8.74199e-09, 8.754252e-09, 8.801573e-09, 8.811972e-09, 8.821614e-09, 
    8.840658e-09, 8.865099e-09, 8.907979e-09, 8.945293e-09, 8.979362e-09, 
    8.976865e-09, 8.977745e-09, 8.985355e-09, 8.966503e-09, 8.98845e-09, 
    8.992133e-09, 8.982503e-09, 9.038398e-09, 9.022428e-09, 9.03877e-09, 
    9.028372e-09, 8.767077e-09, 8.780028e-09, 8.773029e-09, 8.78619e-09, 
    8.776918e-09, 8.818145e-09, 8.830508e-09, 8.888359e-09, 8.864617e-09, 
    8.902406e-09, 8.868457e-09, 8.874472e-09, 8.903636e-09, 8.870292e-09, 
    8.943235e-09, 8.893777e-09, 8.98565e-09, 8.936254e-09, 8.988747e-09, 
    8.979215e-09, 8.994997e-09, 9.009131e-09, 9.026916e-09, 9.059732e-09, 
    9.052133e-09, 9.079579e-09, 8.799337e-09, 8.816136e-09, 8.814658e-09, 
    8.832241e-09, 8.845245e-09, 8.873432e-09, 8.918644e-09, 8.901643e-09, 
    8.932858e-09, 8.939125e-09, 8.891702e-09, 8.920817e-09, 8.827381e-09, 
    8.842473e-09, 8.833488e-09, 8.800662e-09, 8.905558e-09, 8.85172e-09, 
    8.951145e-09, 8.921974e-09, 9.007116e-09, 8.964769e-09, 9.04795e-09, 
    9.083511e-09, 9.11699e-09, 9.156111e-09, 8.825307e-09, 8.813891e-09, 
    8.834332e-09, 8.862613e-09, 8.888859e-09, 8.923752e-09, 8.927325e-09, 
    8.933862e-09, 8.950797e-09, 8.965036e-09, 8.935928e-09, 8.968605e-09, 
    8.845972e-09, 8.910233e-09, 8.809574e-09, 8.83988e-09, 8.860947e-09, 
    8.851706e-09, 8.8997e-09, 8.911011e-09, 8.956984e-09, 8.933219e-09, 
    9.074732e-09, 9.012115e-09, 9.185906e-09, 9.137329e-09, 8.809902e-09, 
    8.825268e-09, 8.878748e-09, 8.853301e-09, 8.926083e-09, 8.944e-09, 
    8.958567e-09, 8.977188e-09, 8.979199e-09, 8.990232e-09, 8.972153e-09, 
    8.989518e-09, 8.923828e-09, 8.953181e-09, 8.872636e-09, 8.892238e-09, 
    8.88322e-09, 8.873329e-09, 8.903859e-09, 8.936385e-09, 8.937082e-09, 
    8.947512e-09, 8.976901e-09, 8.926379e-09, 9.082811e-09, 8.98619e-09, 
    8.842024e-09, 8.87162e-09, 8.87585e-09, 8.864385e-09, 8.942203e-09, 
    8.914005e-09, 8.989963e-09, 8.969433e-09, 9.003072e-09, 8.986356e-09, 
    8.983896e-09, 8.962428e-09, 8.949062e-09, 8.915298e-09, 8.887827e-09, 
    8.866047e-09, 8.871112e-09, 8.895038e-09, 8.938375e-09, 8.97938e-09, 
    8.970397e-09, 9.000516e-09, 8.920805e-09, 8.954227e-09, 8.941308e-09, 
    8.974993e-09, 8.901191e-09, 8.96403e-09, 8.885129e-09, 8.892046e-09, 
    8.913445e-09, 8.956492e-09, 8.966019e-09, 8.976189e-09, 8.969914e-09, 
    8.939476e-09, 8.93449e-09, 8.912926e-09, 8.90697e-09, 8.890541e-09, 
    8.876938e-09, 8.889366e-09, 8.902417e-09, 8.939489e-09, 8.972901e-09, 
    9.009332e-09, 9.01825e-09, 9.060817e-09, 9.026163e-09, 9.083349e-09, 
    9.034726e-09, 9.118903e-09, 8.967675e-09, 9.033299e-09, 8.914419e-09, 
    8.927225e-09, 8.950386e-09, 9.003517e-09, 8.974835e-09, 9.00838e-09, 
    8.934295e-09, 8.895862e-09, 8.885921e-09, 8.867372e-09, 8.886345e-09, 
    8.884802e-09, 8.902959e-09, 8.897125e-09, 8.94072e-09, 8.917302e-09, 
    8.983834e-09, 9.008116e-09, 9.076702e-09, 9.118752e-09, 9.161566e-09, 
    9.180468e-09, 9.186222e-09, 9.188628e-09 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.182616, 6.210857, 6.20536, 6.228186, 6.215517, 6.230473, 6.188334, 
    6.211982, 6.196878, 6.185153, 6.272632, 6.229205, 6.317922, 6.290085, 
    6.360148, 6.313587, 6.369561, 6.358799, 6.391214, 6.381917, 6.423494, 
    6.395508, 6.445103, 6.416802, 6.421226, 6.394587, 6.237926, 6.267216, 
    6.236194, 6.240365, 6.238492, 6.215779, 6.204354, 6.180459, 6.184793, 
    6.202343, 6.242241, 6.228678, 6.262888, 6.262114, 6.300333, 6.283084, 
    6.34753, 6.329173, 6.382306, 6.368918, 6.381677, 6.377806, 6.381727, 
    6.362101, 6.370505, 6.35325, 6.286313, 6.305942, 6.24751, 6.21254, 
    6.189371, 6.172965, 6.175282, 6.179703, 6.202446, 6.223874, 6.240235, 
    6.251194, 6.262003, 6.294799, 6.312192, 6.351248, 6.344186, 6.35615, 
    6.367588, 6.386822, 6.383654, 6.392137, 6.355832, 6.379948, 6.340167, 
    6.351033, 6.264955, 6.232335, 6.218511, 6.206418, 6.177065, 6.197327, 
    6.189335, 6.208356, 6.220463, 6.214473, 6.251493, 6.237085, 6.313224, 
    6.28036, 6.366253, 6.345635, 6.371201, 6.358147, 6.380524, 6.360383, 
    6.395295, 6.402914, 6.397707, 6.417717, 6.359267, 6.381678, 6.214305, 
    6.215282, 6.219832, 6.199845, 6.198624, 6.180341, 6.196606, 6.203541, 
    6.221164, 6.231604, 6.241538, 6.263412, 6.2879, 6.322235, 6.346971, 
    6.363584, 6.353393, 6.36239, 6.352333, 6.347622, 6.400059, 6.370584, 
    6.414836, 6.412383, 6.392339, 6.412659, 6.215968, 6.210348, 6.190866, 
    6.20611, 6.178351, 6.193881, 6.202822, 6.237389, 6.244996, 6.252059, 
    6.26602, 6.283966, 6.315524, 6.343057, 6.368253, 6.366405, 6.367055, 
    6.372693, 6.358736, 6.374986, 6.377717, 6.37058, 6.412054, 6.400189, 
    6.412331, 6.404603, 6.212174, 6.221633, 6.216521, 6.226136, 6.219362, 
    6.249522, 6.258582, 6.301078, 6.283613, 6.311419, 6.286433, 6.290857, 
    6.312332, 6.287781, 6.341539, 6.305068, 6.372912, 6.336387, 6.375205, 
    6.368144, 6.379837, 6.39032, 6.403522, 6.427927, 6.422271, 6.44271, 
    6.235749, 6.248048, 6.246963, 6.259847, 6.269386, 6.29009, 6.323386, 
    6.310852, 6.333871, 6.338499, 6.303531, 6.324989, 6.256286, 6.267357, 
    6.260763, 6.23672, 6.313742, 6.274143, 6.34738, 6.32584, 6.388825, 
    6.357458, 6.419158, 6.445649, 6.470628, 6.499903, 6.254765, 6.2464, 
    6.261379, 6.282144, 6.30144, 6.327153, 6.329786, 6.334612, 6.347121, 
    6.35765, 6.336141, 6.360291, 6.269931, 6.317185, 6.243242, 6.265455, 
    6.280917, 6.274129, 6.30942, 6.317756, 6.351698, 6.334137, 6.439107, 
    6.39254, 6.522237, 6.485841, 6.24348, 6.254735, 6.294003, 6.2753, 
    6.328871, 6.342101, 6.352865, 6.366645, 6.368133, 6.376307, 6.362916, 
    6.375777, 6.327208, 6.348885, 6.289505, 6.303927, 6.297289, 6.290014, 
    6.312484, 6.33648, 6.336989, 6.344697, 6.366451, 6.329088, 6.445138, 
    6.373327, 6.267021, 6.288764, 6.29187, 6.28344, 6.340774, 6.319963, 
    6.376107, 6.360903, 6.385824, 6.373434, 6.371612, 6.355721, 6.34584, 
    6.320918, 6.300682, 6.284661, 6.288384, 6.30599, 6.337949, 6.368269, 
    6.36162, 6.383928, 6.324977, 6.349659, 6.340114, 6.365019, 6.31052, 
    6.356923, 6.298693, 6.303785, 6.319551, 6.351337, 6.358377, 6.365906, 
    6.361259, 6.33876, 6.335077, 6.319167, 6.314779, 6.302676, 6.292667, 
    6.301812, 6.311425, 6.338768, 6.363472, 6.390471, 6.397086, 6.428745, 
    6.402971, 6.44554, 6.409346, 6.472073, 6.359612, 6.408276, 6.320268, 
    6.329713, 6.346823, 6.386161, 6.364902, 6.389767, 6.334933, 6.306599, 
    6.299276, 6.285635, 6.299589, 6.298453, 6.311821, 6.307523, 6.339677, 
    6.322393, 6.371567, 6.38957, 6.440567, 6.471951, 6.503982, 6.518155, 
    6.522471, 6.524277,
  3.950761, 3.970177, 3.966397, 3.982093, 3.97338, 3.983666, 3.954691, 
    3.970951, 3.960565, 3.952504, 4.012669, 3.982794, 4.043364, 4.024673, 
    4.071574, 4.040469, 4.077863, 4.07067, 4.092332, 4.086119, 4.113914, 
    4.095202, 4.12836, 4.109437, 4.112396, 4.094586, 3.988791, 4.008944, 
    3.9876, 3.990469, 3.989181, 3.973561, 3.965707, 3.949277, 3.952256, 
    3.964323, 3.99176, 3.982431, 4.005961, 4.005428, 4.031615, 4.019855, 
    4.063141, 4.050877, 4.086378, 4.077432, 4.085958, 4.083371, 4.085992, 
    4.072877, 4.078493, 4.066963, 4.022078, 4.035361, 3.995384, 3.971336, 
    3.955404, 3.944125, 3.945719, 3.948758, 3.964394, 3.979127, 3.990379, 
    3.997916, 4.005352, 4.02792, 4.039537, 4.065627, 4.060906, 4.068902, 
    4.076543, 4.089397, 4.087279, 4.09295, 4.068687, 4.084804, 4.05822, 
    4.065481, 4.007388, 3.984946, 3.975441, 3.967124, 3.946944, 3.960874, 
    3.955379, 3.968456, 3.976781, 3.972662, 3.998123, 3.988213, 4.040226, 
    4.017982, 4.075651, 4.061875, 4.078957, 4.070234, 4.085188, 4.071728, 
    4.09506, 4.100153, 4.096673, 4.110048, 4.070983, 4.08596, 3.972547, 
    3.973219, 3.976348, 3.962606, 3.961765, 3.949196, 3.960378, 3.965147, 
    3.977263, 3.984443, 3.991275, 4.006322, 4.02317, 4.046244, 4.062767, 
    4.073867, 4.067058, 4.073069, 4.06635, 4.063202, 4.098246, 4.078547, 
    4.108123, 4.106482, 4.093085, 4.106667, 3.97369, 3.969826, 3.956431, 
    3.966911, 3.947828, 3.958505, 3.964653, 3.988423, 3.993654, 3.998512, 
    4.008116, 4.020463, 4.04176, 4.060153, 4.076987, 4.075752, 4.076187, 
    4.079955, 4.070628, 4.081487, 4.083313, 4.078542, 4.106262, 4.098331, 
    4.106447, 4.101281, 3.971081, 3.977586, 3.974071, 3.980683, 3.976025, 
    3.996768, 4.003001, 4.032113, 4.02022, 4.039019, 4.02216, 4.025205, 
    4.039632, 4.023088, 4.059141, 4.034779, 4.080101, 4.0557, 4.081634, 
    4.076914, 4.084728, 4.091735, 4.100559, 4.116876, 4.113093, 4.126759, 
    3.987293, 3.995754, 3.995006, 4.003869, 4.010432, 4.024676, 4.047011, 
    4.038639, 4.054015, 4.057107, 4.033749, 4.048083, 4.00142, 4.009037, 
    4.004499, 3.987962, 4.040571, 4.013706, 4.063041, 4.048651, 4.090736, 
    4.069776, 4.111012, 4.128727, 4.145428, 4.165013, 4.000373, 3.994619, 
    4.004923, 4.01921, 4.032353, 4.049528, 4.051287, 4.054511, 4.062867, 
    4.069902, 4.055533, 4.071667, 4.01081, 4.042871, 3.992448, 4.007729, 
    4.018366, 4.013695, 4.037682, 4.04325, 4.065927, 4.054193, 4.124353, 
    4.093221, 4.179954, 4.155606, 3.992611, 4.000352, 4.027369, 4.0145, 
    4.050675, 4.059514, 4.066705, 4.075914, 4.076907, 4.08237, 4.073421, 
    4.082015, 4.049565, 4.064046, 4.024273, 4.034015, 4.02958, 4.024623, 
    4.039729, 4.05576, 4.056098, 4.061249, 4.075791, 4.05082, 4.12839, 
    4.080385, 4.008804, 4.023766, 4.025901, 4.0201, 4.058627, 4.044725, 
    4.082236, 4.072076, 4.08873, 4.08045, 4.079232, 4.068613, 4.062012, 
    4.045363, 4.031847, 4.02094, 4.023502, 4.035392, 4.056741, 4.076999, 
    4.072556, 4.087463, 4.048074, 4.064564, 4.058187, 4.074827, 4.038418, 
    4.069423, 4.030518, 4.033919, 4.04445, 4.065687, 4.070388, 4.07542, 
    4.072314, 4.057283, 4.054822, 4.044192, 4.041263, 4.033178, 4.026449, 
    4.032601, 4.039023, 4.057288, 4.073794, 4.091836, 4.096257, 4.117426, 
    4.100194, 4.128659, 4.104461, 4.1464, 4.071218, 4.103741, 4.044928, 
    4.051238, 4.06267, 4.088958, 4.074749, 4.091368, 4.054725, 4.0358, 
    4.030908, 4.021611, 4.031116, 4.030357, 4.039286, 4.036415, 4.057895, 
    4.046348, 4.079203, 4.091235, 4.125327, 4.146315, 4.167739, 4.177221, 
    4.18011, 4.181318,
  3.270926, 3.288148, 3.284794, 3.29872, 3.290989, 3.300116, 3.274411, 
    3.288834, 3.279621, 3.272471, 3.32586, 3.299342, 3.353538, 3.33652, 
    3.37937, 3.350888, 3.385132, 3.378543, 3.39839, 3.392696, 3.41817, 
    3.40102, 3.431417, 3.414067, 3.416779, 3.400455, 3.304665, 3.322552, 
    3.303607, 3.306154, 3.30501, 3.29115, 3.284182, 3.269609, 3.272251, 
    3.282954, 3.307299, 3.29902, 3.319905, 3.319432, 3.342784, 3.332242, 
    3.371647, 3.360416, 3.392934, 3.384737, 3.392549, 3.390179, 3.39258, 
    3.380564, 3.385709, 3.375147, 3.334215, 3.346213, 3.310515, 3.289176, 
    3.275043, 3.265041, 3.266454, 3.269149, 3.283017, 3.296088, 3.306073, 
    3.312764, 3.319364, 3.339404, 3.350035, 3.373923, 3.369601, 3.376923, 
    3.383923, 3.3957, 3.393759, 3.398955, 3.376727, 3.391491, 3.367141, 
    3.37379, 3.321171, 3.301251, 3.292818, 3.285439, 3.267541, 3.279895, 
    3.275021, 3.286621, 3.294007, 3.290352, 3.312947, 3.304151, 3.350666, 
    3.330578, 3.383106, 3.370487, 3.386134, 3.378144, 3.391843, 3.379512, 
    3.400889, 3.405557, 3.402367, 3.414627, 3.37883, 3.39255, 3.29025, 
    3.290846, 3.293622, 3.281431, 3.280685, 3.269537, 3.279455, 3.283685, 
    3.294435, 3.300806, 3.306869, 3.320225, 3.335186, 3.356175, 3.371305, 
    3.381472, 3.375234, 3.380741, 3.374586, 3.371703, 3.403808, 3.385758, 
    3.412862, 3.411358, 3.399079, 3.411528, 3.291265, 3.287836, 3.275954, 
    3.28525, 3.268325, 3.277793, 3.283247, 3.304337, 3.30898, 3.313293, 
    3.321818, 3.332781, 3.352071, 3.368911, 3.38433, 3.383198, 3.383597, 
    3.387048, 3.378505, 3.388452, 3.390124, 3.385754, 3.411157, 3.403887, 
    3.411326, 3.406591, 3.28895, 3.294721, 3.291602, 3.297469, 3.293336, 
    3.311744, 3.317276, 3.34324, 3.332566, 3.349561, 3.334289, 3.336992, 
    3.350121, 3.335112, 3.367983, 3.345679, 3.387182, 3.364832, 3.388586, 
    3.384263, 3.391422, 3.397843, 3.405929, 3.420886, 3.417419, 3.429949, 
    3.303335, 3.310844, 3.31018, 3.318048, 3.323874, 3.336523, 3.356878, 
    3.349213, 3.36329, 3.366122, 3.344738, 3.357859, 3.315874, 3.322636, 
    3.318607, 3.303928, 3.350982, 3.326781, 3.371556, 3.358379, 3.396927, 
    3.377723, 3.415511, 3.431753, 3.447074, 3.465045, 3.314944, 3.309837, 
    3.318983, 3.331668, 3.34346, 3.359182, 3.360792, 3.363744, 3.371396, 
    3.37784, 3.36468, 3.379456, 3.32421, 3.353087, 3.30791, 3.321475, 
    3.330919, 3.326771, 3.348338, 3.353435, 3.374198, 3.363453, 3.427742, 
    3.399203, 3.478761, 3.456412, 3.308054, 3.314926, 3.338915, 3.327487, 
    3.360232, 3.368325, 3.374911, 3.383346, 3.384256, 3.389261, 3.381063, 
    3.388936, 3.359215, 3.372476, 3.336165, 3.34498, 3.340922, 3.336476, 
    3.350211, 3.364887, 3.365198, 3.369914, 3.383231, 3.360365, 3.431443, 
    3.38744, 3.322429, 3.335714, 3.33761, 3.332459, 3.367513, 3.354785, 
    3.389138, 3.379831, 3.395089, 3.387501, 3.386386, 3.376659, 3.370613, 
    3.355368, 3.342997, 3.333205, 3.33548, 3.346241, 3.365786, 3.38434, 
    3.380271, 3.393928, 3.357851, 3.37295, 3.36711, 3.38235, 3.349011, 
    3.377399, 3.341781, 3.344893, 3.354532, 3.373978, 3.378285, 3.382894, 
    3.380049, 3.366282, 3.364029, 3.354297, 3.351615, 3.344215, 3.338098, 
    3.343687, 3.349565, 3.366287, 3.381404, 3.397934, 3.401986, 3.42139, 
    3.405594, 3.43169, 3.409503, 3.447964, 3.379043, 3.408845, 3.35497, 
    3.360747, 3.371215, 3.395297, 3.382279, 3.397505, 3.36394, 3.346615, 
    3.342137, 3.333801, 3.342328, 3.341634, 3.349806, 3.347178, 3.366843, 
    3.35627, 3.386359, 3.397383, 3.428636, 3.447887, 3.467548, 3.476253, 
    3.478904, 3.480014,
  2.994152, 3.010521, 3.007335, 3.020567, 3.013221, 3.021894, 2.997474, 
    3.011173, 3.002422, 2.995633, 3.046373, 3.021158, 3.072721, 3.056519, 
    3.097337, 3.070196, 3.10283, 3.096548, 3.115477, 3.110045, 3.134356, 
    3.117986, 3.147009, 3.130439, 3.133028, 3.117448, 3.026217, 3.043226, 
    3.025213, 3.027633, 3.026546, 3.013373, 3.006753, 2.992861, 2.995424, 
    3.005588, 3.028722, 3.020852, 3.04071, 3.04026, 3.062481, 3.052447, 
    3.089975, 3.079274, 3.110272, 3.102455, 3.109905, 3.107644, 3.109934, 
    3.098475, 3.103381, 3.093311, 3.054325, 3.065745, 3.03178, 3.011497, 
    2.998074, 2.988379, 2.989765, 2.992409, 3.005647, 3.018066, 3.027557, 
    3.033918, 3.040195, 3.059262, 3.069385, 3.092144, 3.088025, 3.095003, 
    3.101678, 3.112911, 3.111059, 3.116016, 3.094817, 3.108895, 3.085681, 
    3.092018, 3.041913, 3.022973, 3.014957, 3.007948, 2.990831, 3.002681, 
    2.998054, 3.009071, 3.016088, 3.012616, 3.034092, 3.025729, 3.069985, 
    3.050864, 3.100899, 3.08887, 3.103787, 3.096168, 3.109232, 3.097472, 
    3.117862, 3.122316, 3.119272, 3.130974, 3.096822, 3.109906, 3.012519, 
    3.013085, 3.015723, 3.004141, 3.003433, 2.99279, 3.002264, 3.006281, 
    3.016495, 3.02255, 3.028313, 3.041015, 3.055248, 3.075233, 3.089649, 
    3.099341, 3.093395, 3.098644, 3.092776, 3.090029, 3.120647, 3.103427, 
    3.129289, 3.127853, 3.116135, 3.128015, 3.013482, 3.010225, 2.99894, 
    3.007769, 2.9916, 3.000686, 3.005865, 3.025906, 3.03032, 3.034421, 
    3.042529, 3.05296, 3.071324, 3.087367, 3.102066, 3.100987, 3.101367, 
    3.104658, 3.096512, 3.105997, 3.107592, 3.103424, 3.127661, 3.120723, 
    3.127823, 3.123303, 3.011283, 3.016767, 3.013803, 3.019378, 3.01545, 
    3.032948, 3.038209, 3.062915, 3.052755, 3.068934, 3.054395, 3.056968, 
    3.069466, 3.055179, 3.086483, 3.065237, 3.104786, 3.083479, 3.106125, 
    3.102002, 3.108829, 3.114955, 3.122672, 3.13695, 3.133639, 3.145607, 
    3.024954, 3.032092, 3.031462, 3.038943, 3.044485, 3.056522, 3.075902, 
    3.068603, 3.082012, 3.084709, 3.064342, 3.076837, 3.036875, 3.043307, 
    3.039475, 3.025518, 3.070287, 3.047251, 3.089888, 3.077332, 3.114081, 
    3.095766, 3.131818, 3.147329, 3.161972, 3.179158, 3.035992, 3.031136, 
    3.039833, 3.051901, 3.063125, 3.078098, 3.079632, 3.082444, 3.089736, 
    3.095878, 3.083335, 3.097419, 3.044803, 3.072291, 3.029303, 3.042202, 
    3.051188, 3.047242, 3.067769, 3.072623, 3.092406, 3.082167, 3.143497, 
    3.116252, 3.192284, 3.1709, 3.029441, 3.035974, 3.058798, 3.047922, 
    3.079098, 3.086809, 3.093087, 3.101128, 3.101996, 3.106768, 3.098951, 
    3.106459, 3.07813, 3.090765, 3.056181, 3.064573, 3.060709, 3.056477, 
    3.069553, 3.083533, 3.083829, 3.088323, 3.101016, 3.079225, 3.147032, 
    3.105031, 3.043111, 3.055751, 3.057557, 3.052654, 3.086035, 3.073909, 
    3.106652, 3.097776, 3.112328, 3.105091, 3.104027, 3.094753, 3.08899, 
    3.074465, 3.062684, 3.053364, 3.055529, 3.065773, 3.084389, 3.102076, 
    3.098195, 3.11122, 3.07683, 3.091217, 3.085651, 3.100179, 3.06841, 
    3.095456, 3.061526, 3.064489, 3.073669, 3.092196, 3.096303, 3.100696, 
    3.097984, 3.084862, 3.082715, 3.073445, 3.07089, 3.063844, 3.058021, 
    3.063342, 3.068937, 3.084867, 3.099276, 3.115042, 3.118909, 3.13743, 
    3.12235, 3.147267, 3.12608, 3.162822, 3.097024, 3.125453, 3.074086, 
    3.079589, 3.089563, 3.112525, 3.10011, 3.114632, 3.082631, 3.066128, 
    3.061866, 3.053931, 3.062047, 3.061387, 3.069167, 3.066665, 3.085397, 
    3.075324, 3.104001, 3.114516, 3.144352, 3.162749, 3.181554, 3.189883, 
    3.192422, 3.193483,
  2.977715, 2.994344, 2.991104, 3.004567, 2.997091, 3.005917, 2.981078, 
    2.995006, 2.986108, 2.979208, 3.03086, 3.005168, 3.057434, 3.041213, 
    3.0818, 3.054938, 3.087245, 3.08102, 3.099787, 3.094399, 3.11853, 
    3.102276, 3.131109, 3.11464, 3.117211, 3.101742, 3.01032, 3.027651, 
    3.009297, 3.011761, 3.010655, 2.997246, 2.990511, 2.976447, 2.978995, 
    2.989326, 3.01287, 3.004857, 3.025087, 3.024629, 3.0473, 3.037058, 
    3.07451, 3.063917, 3.094623, 3.086873, 3.094259, 3.092017, 3.094288, 
    3.082929, 3.087791, 3.077813, 3.038974, 3.050538, 3.015986, 2.995336, 
    2.981688, 2.972041, 2.973403, 2.976002, 2.989387, 3.002022, 3.011684, 
    3.018165, 3.024563, 3.044013, 3.054135, 3.076657, 3.072579, 3.079489, 
    3.086103, 3.09724, 3.095404, 3.100322, 3.079305, 3.093258, 3.070258, 
    3.076532, 3.026311, 3.007017, 2.998857, 2.991726, 2.974451, 2.986372, 
    2.981667, 2.992869, 3.000008, 2.996475, 3.018342, 3.009823, 3.054729, 
    3.035442, 3.085331, 3.073415, 3.088193, 3.080643, 3.093591, 3.081936, 
    3.102153, 3.106573, 3.103552, 3.115171, 3.081291, 3.09426, 2.996376, 
    2.996953, 2.999637, 2.987855, 2.987135, 2.976377, 2.985947, 2.990032, 
    3.000422, 3.006585, 3.012455, 3.025398, 3.039916, 3.059919, 3.074186, 
    3.083787, 3.077896, 3.083096, 3.077284, 3.074563, 3.104917, 3.087837, 
    3.113497, 3.112072, 3.100439, 3.112232, 2.997357, 2.994043, 2.982568, 
    2.991545, 2.975208, 2.984343, 2.989608, 3.010003, 3.014499, 3.018677, 
    3.026942, 3.037582, 3.056053, 3.071927, 3.086488, 3.085418, 3.085795, 
    3.089057, 3.080984, 3.090384, 3.091965, 3.087834, 3.111881, 3.104992, 
    3.112041, 3.107554, 2.99512, 3.000699, 2.997683, 3.003357, 2.999359, 
    3.017176, 3.022537, 3.04774, 3.037372, 3.05369, 3.039046, 3.041672, 
    3.054216, 3.039846, 3.071051, 3.050035, 3.089184, 3.068078, 3.090511, 
    3.086425, 3.093193, 3.099268, 3.106927, 3.121109, 3.117819, 3.129714, 
    3.009033, 3.016304, 3.015662, 3.023286, 3.028937, 3.041216, 3.060582, 
    3.053364, 3.066626, 3.069296, 3.049151, 3.061506, 3.021178, 3.027735, 
    3.023828, 3.009607, 3.055027, 3.031756, 3.074423, 3.061996, 3.098402, 
    3.080245, 3.116009, 3.131427, 3.146, 3.163124, 3.020278, 3.01533, 
    3.024194, 3.0365, 3.047949, 3.062753, 3.064271, 3.067054, 3.074273, 
    3.080356, 3.067936, 3.081883, 3.029259, 3.05701, 3.013462, 3.026608, 
    3.035773, 3.031748, 3.052539, 3.057338, 3.076917, 3.06678, 3.127616, 
    3.100555, 3.176219, 3.154892, 3.013603, 3.02026, 3.04354, 3.032442, 
    3.063743, 3.071375, 3.077591, 3.085558, 3.086418, 3.091149, 3.0834, 
    3.090842, 3.062785, 3.075292, 3.040869, 3.049379, 3.045491, 3.041171, 
    3.054303, 3.068131, 3.068425, 3.072873, 3.085445, 3.063869, 3.13113, 
    3.089424, 3.027535, 3.040429, 3.042273, 3.037269, 3.070609, 3.05861, 
    3.091033, 3.082237, 3.096662, 3.089486, 3.088432, 3.079241, 3.073534, 
    3.05916, 3.047507, 3.037994, 3.040204, 3.050565, 3.068979, 3.086497, 
    3.082651, 3.095564, 3.061499, 3.075739, 3.070228, 3.084617, 3.053173, 
    3.079936, 3.046326, 3.049297, 3.058372, 3.076709, 3.080777, 3.08513, 
    3.082443, 3.069447, 3.067322, 3.058151, 3.055624, 3.048659, 3.042747, 
    3.048163, 3.053694, 3.069452, 3.083723, 3.099355, 3.103192, 3.121584, 
    3.106607, 3.131364, 3.110308, 3.146844, 3.081491, 3.109687, 3.058785, 
    3.064229, 3.074101, 3.096858, 3.084549, 3.098948, 3.067239, 3.050916, 
    3.046672, 3.038572, 3.046858, 3.046183, 3.053921, 3.051448, 3.069976, 
    3.06001, 3.088406, 3.098833, 3.128467, 3.146773, 3.165513, 3.173823, 
    3.176357, 3.177417,
  2.97641, 2.994802, 2.991215, 3.006129, 2.997844, 3.007627, 2.980127, 
    2.995535, 2.985687, 2.978059, 3.035337, 3.006797, 3.065332, 3.046869, 
    3.093514, 3.062451, 3.099825, 3.09261, 3.114383, 3.108126, 3.136191, 
    3.117277, 3.150863, 3.13166, 3.134655, 3.116655, 3.012512, 3.031767, 
    3.011376, 3.014111, 3.012883, 2.998015, 2.990559, 2.975009, 2.977824, 
    2.989248, 3.015342, 3.006452, 3.028916, 3.028406, 3.053657, 3.042239, 
    3.085071, 3.072821, 3.108387, 3.099394, 3.107964, 3.105362, 3.107998, 
    3.094822, 3.100459, 3.088896, 3.044374, 3.057376, 3.018802, 2.9959, 
    2.980801, 2.970106, 2.971648, 2.974518, 2.989315, 3.003308, 3.014026, 
    3.021222, 3.028333, 3.049989, 3.061525, 3.087557, 3.082837, 3.090837, 
    3.098501, 3.111426, 3.109293, 3.115005, 3.090624, 3.106801, 3.080153, 
    3.087413, 3.030277, 3.008847, 2.9998, 2.991904, 2.972805, 2.985979, 
    2.980778, 2.993169, 3.001076, 2.997162, 3.021419, 3.01196, 3.062211, 
    3.04044, 3.097606, 3.083805, 3.100925, 3.092174, 3.107189, 3.093671, 
    3.117133, 3.122272, 3.118759, 3.132279, 3.092924, 3.107965, 2.997053, 
    2.997691, 3.000664, 2.98762, 2.986824, 2.974932, 2.98551, 2.990029, 
    3.001535, 3.008368, 3.014881, 3.029261, 3.045424, 3.068202, 3.084697, 
    3.095816, 3.088992, 3.095016, 3.088283, 3.085133, 3.120346, 3.100512, 
    3.13033, 3.12867, 3.115141, 3.128857, 2.998139, 2.994469, 2.981773, 
    2.991703, 2.973641, 2.983736, 2.98956, 3.012159, 3.017151, 3.021791, 
    3.030979, 3.042823, 3.063739, 3.082083, 3.098948, 3.097708, 3.098144, 
    3.101927, 3.092568, 3.103467, 3.105301, 3.100509, 3.128448, 3.120434, 
    3.128635, 3.123413, 2.995661, 3.001842, 2.9985, 3.004788, 3.000357, 
    3.020123, 3.026081, 3.05415, 3.042589, 3.061011, 3.044454, 3.04738, 
    3.061618, 3.045345, 3.081069, 3.056795, 3.102074, 3.07763, 3.103614, 
    3.098874, 3.106726, 3.113781, 3.122683, 3.139197, 3.135363, 3.149235, 
    3.011084, 3.019155, 3.018442, 3.026913, 3.033198, 3.046873, 3.068968, 
    3.060635, 3.075953, 3.07904, 3.055776, 3.070035, 3.02457, 3.03186, 
    3.027516, 3.01172, 3.062555, 3.036335, 3.084971, 3.070602, 3.112774, 
    3.091712, 3.133255, 3.151234, 3.168177, 3.187602, 3.02357, 3.018073, 
    3.027922, 3.041618, 3.05439, 3.071476, 3.07323, 3.076447, 3.084797, 
    3.091841, 3.077466, 3.09361, 3.033556, 3.064843, 3.015999, 3.030607, 
    3.040808, 3.036326, 3.059684, 3.065223, 3.087858, 3.07613, 3.146785, 
    3.115276, 3.202493, 3.178257, 3.016156, 3.02355, 3.049462, 3.037099, 
    3.07262, 3.081444, 3.088639, 3.097869, 3.098867, 3.104354, 3.095369, 
    3.103998, 3.071512, 3.085976, 3.046485, 3.056039, 3.051639, 3.046822, 
    3.061719, 3.077692, 3.078032, 3.083177, 3.097738, 3.072765, 3.150886, 
    3.102352, 3.031639, 3.045995, 3.04805, 3.042475, 3.080558, 3.066691, 
    3.10422, 3.09402, 3.110754, 3.102425, 3.101202, 3.09055, 3.083942, 
    3.067325, 3.053887, 3.043282, 3.045744, 3.057407, 3.078672, 3.098958, 
    3.0945, 3.109478, 3.070027, 3.086494, 3.080117, 3.096779, 3.060415, 
    3.091353, 3.052569, 3.055945, 3.066416, 3.087616, 3.092328, 3.097373, 
    3.094259, 3.079214, 3.076757, 3.066161, 3.063244, 3.055209, 3.048579, 
    3.054637, 3.061016, 3.079219, 3.095742, 3.113882, 3.118341, 3.139751, 
    3.122311, 3.15116, 3.126616, 3.169132, 3.093155, 3.125894, 3.066893, 
    3.073181, 3.084598, 3.110981, 3.0967, 3.113408, 3.076661, 3.057812, 
    3.052956, 3.043926, 3.053163, 3.05241, 3.061279, 3.058425, 3.079826, 
    3.068307, 3.101171, 3.113275, 3.147779, 3.169052, 3.190317, 3.199766, 
    3.20265, 3.203856,
  3.255228, 3.278703, 3.274116, 3.293223, 3.282598, 3.295146, 3.259963, 
    3.279643, 3.267055, 3.257328, 3.330405, 3.294079, 3.368177, 3.344887, 
    3.403971, 3.364535, 3.412028, 3.402818, 3.430673, 3.422649, 3.458757, 
    3.434388, 3.477758, 3.452906, 3.456772, 3.43359, 3.301424, 3.32593, 
    3.299963, 3.303481, 3.301901, 3.282818, 3.273277, 3.253444, 3.257029, 
    3.271602, 3.305065, 3.293637, 3.322361, 3.321723, 3.353435, 3.339067, 
    3.393216, 3.377659, 3.422983, 3.411477, 3.422441, 3.419109, 3.422485, 
    3.40564, 3.412838, 3.398085, 3.34175, 3.358125, 3.30952, 3.280109, 
    3.260822, 3.247258, 3.249169, 3.252819, 3.271688, 3.289602, 3.303371, 
    3.31264, 3.321631, 3.348815, 3.363365, 3.396379, 3.390374, 3.400558, 
    3.410336, 3.426878, 3.424145, 3.43147, 3.400286, 3.420952, 3.386963, 
    3.396196, 3.324064, 3.296712, 3.285105, 3.274997, 3.250641, 3.267427, 
    3.260792, 3.276615, 3.286741, 3.281725, 3.312894, 3.300714, 3.364231, 
    3.336807, 3.409193, 3.391605, 3.413434, 3.402262, 3.421448, 3.404171, 
    3.434203, 3.44081, 3.436293, 3.453705, 3.403219, 3.422442, 3.281585, 
    3.282403, 3.286213, 3.269522, 3.268506, 3.253347, 3.266828, 3.2726, 
    3.287329, 3.296098, 3.304471, 3.322793, 3.343069, 3.371808, 3.39274, 
    3.406909, 3.398207, 3.405887, 3.397304, 3.393295, 3.438333, 3.412906, 
    3.45119, 3.44905, 3.431645, 3.449291, 3.282976, 3.278278, 3.262061, 
    3.27474, 3.251703, 3.264564, 3.272, 3.30097, 3.307394, 3.313373, 
    3.324944, 3.3398, 3.366162, 3.389416, 3.410907, 3.409323, 3.409881, 
    3.414715, 3.402765, 3.416684, 3.419032, 3.412902, 3.448764, 3.438446, 
    3.449005, 3.442279, 3.279804, 3.287722, 3.283439, 3.291501, 3.285819, 
    3.311223, 3.318814, 3.354056, 3.339507, 3.362715, 3.34185, 3.34553, 
    3.363481, 3.342971, 3.388127, 3.357393, 3.414903, 3.38376, 3.416873, 
    3.410813, 3.420856, 3.4299, 3.441339, 3.462643, 3.457687, 3.475646, 
    3.299588, 3.309975, 3.309057, 3.319855, 3.327723, 3.344892, 3.372778, 
    3.36224, 3.381631, 3.385549, 3.356108, 3.374129, 3.316926, 3.326047, 
    3.320609, 3.300406, 3.364665, 3.331656, 3.393088, 3.374847, 3.428608, 
    3.401673, 3.454965, 3.47824, 3.500414, 3.526686, 3.315667, 3.308582, 
    3.321118, 3.338286, 3.35436, 3.375955, 3.378178, 3.382258, 3.392868, 
    3.401838, 3.383552, 3.404093, 3.328172, 3.367558, 3.305911, 3.324477, 
    3.337269, 3.331645, 3.36104, 3.368038, 3.396763, 3.381856, 3.472469, 
    3.431818, 3.546572, 3.514027, 3.306113, 3.315642, 3.348151, 3.332614, 
    3.377405, 3.388604, 3.397757, 3.409529, 3.410804, 3.41782, 3.406337, 
    3.417364, 3.376001, 3.394368, 3.344404, 3.356439, 3.350893, 3.344829, 
    3.36361, 3.383839, 3.384271, 3.390808, 3.409361, 3.377589, 3.477788, 
    3.415259, 3.32577, 3.343788, 3.346374, 3.339363, 3.387478, 3.369896, 
    3.417648, 3.404617, 3.426017, 3.415351, 3.413788, 3.400192, 3.391779, 
    3.370699, 3.353725, 3.340378, 3.343472, 3.358165, 3.385083, 3.41092, 
    3.405229, 3.424382, 3.37412, 3.395027, 3.386918, 3.408137, 3.361962, 
    3.401216, 3.352065, 3.35632, 3.369548, 3.396456, 3.402459, 3.408896, 
    3.404921, 3.385771, 3.382652, 3.369225, 3.365537, 3.355393, 3.347039, 
    3.354671, 3.362721, 3.385778, 3.406813, 3.430029, 3.435755, 3.463359, 
    3.44086, 3.478143, 3.446403, 3.501702, 3.403513, 3.445472, 3.370152, 
    3.378116, 3.392614, 3.426307, 3.408037, 3.429421, 3.382529, 3.358676, 
    3.352552, 3.341187, 3.352813, 3.351864, 3.363053, 3.35945, 3.386549, 
    3.371942, 3.413749, 3.429251, 3.473757, 3.501594, 3.530372, 3.54297, 
    3.546779, 3.548374,
  3.812406, 3.852937, 3.844965, 3.878337, 3.859725, 3.88172, 3.820528, 
    3.854572, 3.832743, 3.816005, 3.945441, 3.879843, 4.016919, 3.972602, 
    4.084902, 4.009935, 4.100404, 4.082693, 4.136674, 4.120996, 4.192387, 
    4.143969, 4.230847, 4.18067, 4.188406, 4.1424, 3.892799, 3.937108, 
    3.890217, 3.89644, 3.893644, 3.860109, 3.843509, 3.809353, 3.815492, 
    3.840606, 3.899247, 3.879064, 3.930483, 3.929301, 3.988773, 3.961651, 
    4.064367, 4.034976, 4.121647, 4.099342, 4.120593, 4.114114, 4.120677, 
    4.088106, 4.101969, 4.073642, 3.966692, 3.997694, 3.90716, 3.855384, 
    3.822004, 3.798792, 3.802051, 3.808284, 3.840755, 3.871978, 3.896246, 
    3.912715, 3.929131, 3.980019, 4.007695, 4.070389, 4.058971, 4.078366, 
    4.097142, 4.129247, 4.123911, 4.138238, 4.077847, 4.117694, 4.052509, 
    4.07004, 3.933642, 3.88448, 3.864103, 3.846494, 3.804561, 3.833386, 
    3.821953, 3.849304, 3.866965, 3.858202, 3.913168, 3.891545, 4.009353, 
    3.95741, 4.094939, 4.061306, 4.103121, 4.081627, 4.11866, 4.085287, 
    4.143606, 4.156632, 4.147718, 4.182267, 4.083461, 4.120594, 3.857958, 
    3.859383, 3.866041, 3.837007, 3.835249, 3.809186, 3.832352, 3.842335, 
    3.867995, 3.883397, 3.898195, 3.931284, 3.969176, 4.023901, 4.063463, 
    4.090543, 4.073874, 4.088581, 4.072152, 4.064517, 4.151739, 4.1021, 
    4.177246, 4.172981, 4.138581, 4.173461, 3.860385, 3.852197, 3.824136, 
    3.846048, 3.806376, 3.828447, 3.841296, 3.891997, 3.90338, 3.914023, 
    3.935276, 3.963027, 4.013052, 4.057153, 4.098241, 4.09519, 4.096263, 
    4.105597, 4.082591, 4.10941, 4.113964, 4.102092, 4.172411, 4.151961, 
    4.17289, 4.159537, 3.854853, 3.868683, 3.861193, 3.875311, 3.865351, 
    3.910191, 3.923916, 3.989953, 3.962476, 4.006454, 3.966881, 3.973814, 
    4.007918, 3.968991, 4.054713, 3.996298, 4.105961, 4.046458, 4.109776, 
    4.098061, 4.117509, 4.135159, 4.157679, 4.200201, 4.190239, 4.226541, 
    3.889554, 3.907969, 3.906336, 3.925842, 3.940444, 3.972611, 4.025768, 
    4.005546, 4.042444, 4.049837, 3.993853, 4.028356, 3.920427, 3.937326, 
    3.927238, 3.891, 4.010185, 3.947776, 4.064125, 4.029701, 4.132629, 
    4.0805, 4.184786, 4.231831, 4.27755, 4.332259, 3.918119, 3.90549, 
    3.928179, 3.960185, 3.99053, 4.031777, 4.03595, 4.043626, 4.063705, 
    4.080815, 4.046065, 4.085137, 3.94128, 4.015731, 3.900748, 3.93441, 
    3.958277, 3.947755, 4.003252, 4.016653, 4.07112, 4.042868, 4.220078, 
    4.13892, 4.374619, 4.30607, 3.901105, 3.918074, 3.978764, 3.949564, 
    4.034498, 4.055614, 4.073017, 4.095586, 4.098042, 4.111611, 4.089445, 
    4.110728, 4.031864, 4.066558, 3.971691, 3.994484, 3.983952, 3.972491, 
    4.008164, 4.046607, 4.047422, 4.059793, 4.095263, 4.034842, 4.230909, 
    4.106649, 3.936811, 3.97053, 3.975406, 3.962205, 4.053483, 4.020221, 
    4.111279, 4.086141, 4.127565, 4.106829, 4.103804, 4.077666, 4.061638, 
    4.021765, 3.989325, 3.964112, 3.969935, 3.99777, 4.048955, 4.098268, 
    4.087317, 4.124373, 4.028338, 4.067812, 4.052424, 4.092906, 4.005013, 
    4.079625, 3.986174, 3.994257, 4.019553, 4.070534, 4.082005, 4.094367, 
    4.086725, 4.050255, 4.044368, 4.018932, 4.011854, 3.992493, 3.976662, 
    3.99112, 4.006464, 4.050269, 4.09036, 4.135413, 4.146659, 4.201644, 
    4.156731, 4.231634, 4.167716, 4.280234, 4.084024, 4.165867, 4.020713, 
    4.035833, 4.063223, 4.128132, 4.092713, 4.134222, 4.044137, 3.998742, 
    3.987098, 3.965633, 3.987592, 3.985793, 4.0071, 4.000218, 4.051725, 
    4.024158, 4.103729, 4.133888, 4.222695, 4.280008, 4.339909, 4.366786, 
    4.375069, 4.378547,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24855.56, 24876.36, 24872.28, 24889.3, 24879.82, 24891.02, 24859.74, 
    24877.19, 24866.02, 24857.41, 24923.11, 24890.07, 24958.46, 24936.61, 
    24991.94, 24955.03, 24999.53, 24990.86, 25017.19, 25009.57, 25044.06, 
    25020.72, 25062.45, 25038.44, 25042.15, 25019.96, 24896.65, 24918.95, 
    24895.34, 24898.49, 24897.07, 24880.02, 24871.54, 24853.98, 24857.15, 
    24870.05, 24899.91, 24889.67, 24915.64, 24915.05, 24944.61, 24931.17, 
    24981.86, 24967.35, 25009.89, 24999.01, 25009.37, 25006.22, 25009.42, 
    24993.51, 25000.29, 24986.42, 24933.68, 24949.01, 24903.91, 24877.61, 
    24860.5, 24848.52, 24850.21, 24853.43, 24870.12, 24886.07, 24898.39, 
    24906.72, 24914.96, 24940.28, 24953.93, 24984.82, 24979.2, 24988.74, 
    24997.94, 25013.58, 25010.99, 25017.95, 24988.48, 25007.96, 24976.01, 
    24984.65, 24917.22, 24892.43, 24882.06, 24873.06, 24851.51, 24866.35, 
    24860.47, 24874.5, 24883.52, 24879.05, 24906.95, 24896.01, 24954.74, 
    24929.06, 24996.86, 24980.35, 25000.86, 24990.34, 25008.43, 24992.13, 
    25020.55, 25026.85, 25022.54, 25039.21, 24991.24, 25009.38, 24878.92, 
    24879.65, 24883.04, 24868.21, 24867.3, 24853.9, 24865.82, 24870.93, 
    24884.04, 24891.88, 24899.38, 24916.04, 24934.91, 24961.88, 24981.41, 
    24994.71, 24986.53, 24993.75, 24985.69, 24981.93, 25024.48, 25000.36, 
    25036.79, 25034.74, 25018.11, 25034.97, 24880.16, 24875.98, 24861.6, 
    24872.84, 24852.45, 24863.81, 24870.4, 24896.24, 24902, 24907.38, 
    24918.03, 24931.86, 24956.56, 24978.3, 24998.47, 24996.98, 24997.51, 
    25002.07, 24990.81, 25003.93, 25006.15, 25000.35, 25034.46, 25024.59, 
    25034.69, 25028.25, 24877.34, 24884.39, 24880.57, 24887.77, 24882.69, 
    24905.45, 24912.35, 24945.2, 24931.58, 24953.32, 24933.77, 24937.21, 
    24954.04, 24934.82, 24977.1, 24948.32, 25002.24, 24973.03, 25004.11, 
    24998.38, 25007.87, 25016.45, 25027.36, 25047.81, 25043.04, 25060.4, 
    24895, 24904.32, 24903.5, 24913.32, 24920.61, 24936.61, 24962.8, 
    24952.87, 24971.04, 24974.7, 24947.12, 24964.07, 24910.6, 24919.06, 
    24914.01, 24895.73, 24955.15, 24924.27, 24981.74, 24964.73, 25015.22, 
    24989.79, 25040.42, 25062.92, 25084.58, 25110.33, 24909.45, 24903.07, 
    24914.48, 24930.45, 24945.48, 24965.76, 24967.83, 24971.63, 24981.53, 
    24989.94, 24972.83, 24992.06, 24921.03, 24957.88, 24900.67, 24917.6, 
    24929.5, 24924.26, 24951.75, 24958.33, 24985.18, 24971.25, 25057.31, 
    25018.28, 25130.15, 25097.97, 24900.85, 24909.42, 24939.66, 24925.16, 
    24967.11, 24977.54, 24986.11, 24997.17, 24998.38, 25005, 24994.17, 
    25004.57, 24965.81, 24982.94, 24936.16, 24947.43, 24942.23, 24936.55, 
    24954.16, 24973.1, 24973.5, 24979.61, 24997.02, 24967.28, 25062.48, 
    25002.58, 24918.8, 24935.58, 24938, 24931.45, 24976.49, 24960.08, 
    25004.84, 24992.55, 25012.77, 25002.67, 25001.19, 24988.39, 24980.51, 
    24960.84, 24944.88, 24932.4, 24935.29, 24949.05, 24974.26, 24998.49, 
    24993.13, 25011.21, 24964.06, 24983.55, 24975.97, 24995.86, 24952.61, 
    24989.36, 24943.33, 24947.32, 24959.75, 24984.89, 24990.52, 24996.58, 
    24992.84, 24974.9, 24971.99, 24959.45, 24955.97, 24946.45, 24938.62, 
    24945.77, 24953.33, 24974.91, 24994.62, 25016.58, 25022.03, 25048.5, 
    25026.9, 25062.82, 25032.2, 25085.84, 24991.51, 25031.31, 24960.32, 
    24967.77, 24981.29, 25013.04, 24995.77, 25016, 24971.88, 24949.53, 
    24943.79, 24933.15, 24944.03, 24943.14, 24953.64, 24950.25, 24975.63, 
    24962.01, 25001.15, 25015.84, 25058.56, 25085.74, 25113.93, 25126.5, 
    25130.36, 25131.97 ;

 HCSOI =
  24855.56, 24876.36, 24872.28, 24889.3, 24879.82, 24891.02, 24859.74, 
    24877.19, 24866.02, 24857.41, 24923.11, 24890.07, 24958.46, 24936.61, 
    24991.94, 24955.03, 24999.53, 24990.86, 25017.19, 25009.57, 25044.06, 
    25020.72, 25062.45, 25038.44, 25042.15, 25019.96, 24896.65, 24918.95, 
    24895.34, 24898.49, 24897.07, 24880.02, 24871.54, 24853.98, 24857.15, 
    24870.05, 24899.91, 24889.67, 24915.64, 24915.05, 24944.61, 24931.17, 
    24981.86, 24967.35, 25009.89, 24999.01, 25009.37, 25006.22, 25009.42, 
    24993.51, 25000.29, 24986.42, 24933.68, 24949.01, 24903.91, 24877.61, 
    24860.5, 24848.52, 24850.21, 24853.43, 24870.12, 24886.07, 24898.39, 
    24906.72, 24914.96, 24940.28, 24953.93, 24984.82, 24979.2, 24988.74, 
    24997.94, 25013.58, 25010.99, 25017.95, 24988.48, 25007.96, 24976.01, 
    24984.65, 24917.22, 24892.43, 24882.06, 24873.06, 24851.51, 24866.35, 
    24860.47, 24874.5, 24883.52, 24879.05, 24906.95, 24896.01, 24954.74, 
    24929.06, 24996.86, 24980.35, 25000.86, 24990.34, 25008.43, 24992.13, 
    25020.55, 25026.85, 25022.54, 25039.21, 24991.24, 25009.38, 24878.92, 
    24879.65, 24883.04, 24868.21, 24867.3, 24853.9, 24865.82, 24870.93, 
    24884.04, 24891.88, 24899.38, 24916.04, 24934.91, 24961.88, 24981.41, 
    24994.71, 24986.53, 24993.75, 24985.69, 24981.93, 25024.48, 25000.36, 
    25036.79, 25034.74, 25018.11, 25034.97, 24880.16, 24875.98, 24861.6, 
    24872.84, 24852.45, 24863.81, 24870.4, 24896.24, 24902, 24907.38, 
    24918.03, 24931.86, 24956.56, 24978.3, 24998.47, 24996.98, 24997.51, 
    25002.07, 24990.81, 25003.93, 25006.15, 25000.35, 25034.46, 25024.59, 
    25034.69, 25028.25, 24877.34, 24884.39, 24880.57, 24887.77, 24882.69, 
    24905.45, 24912.35, 24945.2, 24931.58, 24953.32, 24933.77, 24937.21, 
    24954.04, 24934.82, 24977.1, 24948.32, 25002.24, 24973.03, 25004.11, 
    24998.38, 25007.87, 25016.45, 25027.36, 25047.81, 25043.04, 25060.4, 
    24895, 24904.32, 24903.5, 24913.32, 24920.61, 24936.61, 24962.8, 
    24952.87, 24971.04, 24974.7, 24947.12, 24964.07, 24910.6, 24919.06, 
    24914.01, 24895.73, 24955.15, 24924.27, 24981.74, 24964.73, 25015.22, 
    24989.79, 25040.42, 25062.92, 25084.58, 25110.33, 24909.45, 24903.07, 
    24914.48, 24930.45, 24945.48, 24965.76, 24967.83, 24971.63, 24981.53, 
    24989.94, 24972.83, 24992.06, 24921.03, 24957.88, 24900.67, 24917.6, 
    24929.5, 24924.26, 24951.75, 24958.33, 24985.18, 24971.25, 25057.31, 
    25018.28, 25130.15, 25097.97, 24900.85, 24909.42, 24939.66, 24925.16, 
    24967.11, 24977.54, 24986.11, 24997.17, 24998.38, 25005, 24994.17, 
    25004.57, 24965.81, 24982.94, 24936.16, 24947.43, 24942.23, 24936.55, 
    24954.16, 24973.1, 24973.5, 24979.61, 24997.02, 24967.28, 25062.48, 
    25002.58, 24918.8, 24935.58, 24938, 24931.45, 24976.49, 24960.08, 
    25004.84, 24992.55, 25012.77, 25002.67, 25001.19, 24988.39, 24980.51, 
    24960.84, 24944.88, 24932.4, 24935.29, 24949.05, 24974.26, 24998.49, 
    24993.13, 25011.21, 24964.06, 24983.55, 24975.97, 24995.86, 24952.61, 
    24989.36, 24943.33, 24947.32, 24959.75, 24984.89, 24990.52, 24996.58, 
    24992.84, 24974.9, 24971.99, 24959.45, 24955.97, 24946.45, 24938.62, 
    24945.77, 24953.33, 24974.91, 24994.62, 25016.58, 25022.03, 25048.5, 
    25026.9, 25062.82, 25032.2, 25085.84, 24991.51, 25031.31, 24960.32, 
    24967.77, 24981.29, 25013.04, 24995.77, 25016, 24971.88, 24949.53, 
    24943.79, 24933.15, 24944.03, 24943.14, 24953.64, 24950.25, 24975.63, 
    24962.01, 25001.15, 25015.84, 25058.56, 25085.74, 25113.93, 25126.5, 
    25130.36, 25131.97 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.194416e-08, 6.221921e-08, 6.216575e-08, 6.238761e-08, 6.226454e-08, 
    6.240981e-08, 6.199993e-08, 6.223013e-08, 6.208317e-08, 6.196893e-08, 
    6.281821e-08, 6.239751e-08, 6.325536e-08, 6.298698e-08, 6.366125e-08, 
    6.321359e-08, 6.375153e-08, 6.364835e-08, 6.395895e-08, 6.386996e-08, 
    6.426725e-08, 6.400002e-08, 6.447324e-08, 6.420344e-08, 6.424563e-08, 
    6.39912e-08, 6.248218e-08, 6.276583e-08, 6.246538e-08, 6.250582e-08, 
    6.248767e-08, 6.226708e-08, 6.215591e-08, 6.192315e-08, 6.19654e-08, 
    6.213637e-08, 6.2524e-08, 6.239242e-08, 6.272409e-08, 6.27166e-08, 
    6.308589e-08, 6.291938e-08, 6.354018e-08, 6.336372e-08, 6.387368e-08, 
    6.374542e-08, 6.386765e-08, 6.383059e-08, 6.386814e-08, 6.368003e-08, 
    6.376062e-08, 6.359511e-08, 6.295056e-08, 6.313996e-08, 6.25751e-08, 
    6.223551e-08, 6.201002e-08, 6.185e-08, 6.187263e-08, 6.191575e-08, 
    6.213737e-08, 6.234576e-08, 6.250459e-08, 6.261083e-08, 6.271553e-08, 
    6.303241e-08, 6.320018e-08, 6.357585e-08, 6.350807e-08, 6.362291e-08, 
    6.373266e-08, 6.39169e-08, 6.388658e-08, 6.396775e-08, 6.361989e-08, 
    6.385107e-08, 6.346945e-08, 6.357381e-08, 6.274394e-08, 6.242792e-08, 
    6.229357e-08, 6.217602e-08, 6.189002e-08, 6.208752e-08, 6.200966e-08, 
    6.219491e-08, 6.231262e-08, 6.22544e-08, 6.261374e-08, 6.247403e-08, 
    6.321012e-08, 6.289304e-08, 6.371985e-08, 6.352198e-08, 6.376729e-08, 
    6.364211e-08, 6.38566e-08, 6.366356e-08, 6.399797e-08, 6.407078e-08, 
    6.402102e-08, 6.421219e-08, 6.365286e-08, 6.386765e-08, 6.225277e-08, 
    6.226226e-08, 6.23065e-08, 6.211204e-08, 6.210015e-08, 6.192198e-08, 
    6.208052e-08, 6.214803e-08, 6.231944e-08, 6.242083e-08, 6.251722e-08, 
    6.272915e-08, 6.296587e-08, 6.329692e-08, 6.353481e-08, 6.369427e-08, 
    6.359649e-08, 6.368282e-08, 6.358631e-08, 6.354109e-08, 6.40435e-08, 
    6.376137e-08, 6.41847e-08, 6.416128e-08, 6.396969e-08, 6.416391e-08, 
    6.226892e-08, 6.221429e-08, 6.202459e-08, 6.217304e-08, 6.190258e-08, 
    6.205396e-08, 6.214101e-08, 6.247694e-08, 6.255076e-08, 6.26192e-08, 
    6.27544e-08, 6.29279e-08, 6.32323e-08, 6.349719e-08, 6.373904e-08, 
    6.372132e-08, 6.372756e-08, 6.378159e-08, 6.364776e-08, 6.380356e-08, 
    6.38297e-08, 6.376134e-08, 6.415814e-08, 6.404477e-08, 6.416078e-08, 
    6.408697e-08, 6.223205e-08, 6.232399e-08, 6.227431e-08, 6.236773e-08, 
    6.230191e-08, 6.259458e-08, 6.268234e-08, 6.309303e-08, 6.292449e-08, 
    6.319274e-08, 6.295173e-08, 6.299444e-08, 6.320148e-08, 6.296477e-08, 
    6.348257e-08, 6.313149e-08, 6.378369e-08, 6.343302e-08, 6.380566e-08, 
    6.3738e-08, 6.385004e-08, 6.395038e-08, 6.407663e-08, 6.430958e-08, 
    6.425564e-08, 6.445048e-08, 6.246106e-08, 6.258032e-08, 6.256982e-08, 
    6.269464e-08, 6.278695e-08, 6.298706e-08, 6.330801e-08, 6.318732e-08, 
    6.340892e-08, 6.345341e-08, 6.311675e-08, 6.332343e-08, 6.266014e-08, 
    6.276728e-08, 6.27035e-08, 6.247047e-08, 6.321512e-08, 6.283292e-08, 
    6.353874e-08, 6.333165e-08, 6.393607e-08, 6.363545e-08, 6.422594e-08, 
    6.447839e-08, 6.471606e-08, 6.499378e-08, 6.264541e-08, 6.256438e-08, 
    6.270949e-08, 6.291025e-08, 6.309657e-08, 6.334428e-08, 6.336963e-08, 
    6.341604e-08, 6.353626e-08, 6.363734e-08, 6.34307e-08, 6.366268e-08, 
    6.279212e-08, 6.32483e-08, 6.253374e-08, 6.274887e-08, 6.289842e-08, 
    6.283283e-08, 6.317353e-08, 6.325383e-08, 6.358018e-08, 6.341148e-08, 
    6.441608e-08, 6.397156e-08, 6.52053e-08, 6.486045e-08, 6.253607e-08, 
    6.264514e-08, 6.302479e-08, 6.284415e-08, 6.336082e-08, 6.348802e-08, 
    6.359143e-08, 6.372361e-08, 6.373789e-08, 6.381621e-08, 6.368786e-08, 
    6.381114e-08, 6.334481e-08, 6.355319e-08, 6.298141e-08, 6.312055e-08, 
    6.305654e-08, 6.298632e-08, 6.320305e-08, 6.343395e-08, 6.34389e-08, 
    6.351294e-08, 6.372157e-08, 6.336292e-08, 6.447343e-08, 6.378752e-08, 
    6.276409e-08, 6.297419e-08, 6.300422e-08, 6.292283e-08, 6.347526e-08, 
    6.327508e-08, 6.38143e-08, 6.366856e-08, 6.390736e-08, 6.37887e-08, 
    6.377123e-08, 6.361883e-08, 6.352395e-08, 6.328425e-08, 6.308925e-08, 
    6.293464e-08, 6.297059e-08, 6.314043e-08, 6.344808e-08, 6.373917e-08, 
    6.367541e-08, 6.388921e-08, 6.332336e-08, 6.356061e-08, 6.34689e-08, 
    6.370803e-08, 6.318411e-08, 6.36302e-08, 6.307009e-08, 6.31192e-08, 
    6.327111e-08, 6.357669e-08, 6.364433e-08, 6.371651e-08, 6.367197e-08, 
    6.34559e-08, 6.34205e-08, 6.326741e-08, 6.322514e-08, 6.310851e-08, 
    6.301195e-08, 6.310017e-08, 6.319282e-08, 6.345599e-08, 6.369318e-08, 
    6.39518e-08, 6.401511e-08, 6.431729e-08, 6.407128e-08, 6.447725e-08, 
    6.413207e-08, 6.472964e-08, 6.365608e-08, 6.412193e-08, 6.327802e-08, 
    6.336893e-08, 6.353335e-08, 6.391052e-08, 6.370691e-08, 6.394504e-08, 
    6.341912e-08, 6.314629e-08, 6.307572e-08, 6.294403e-08, 6.307872e-08, 
    6.306777e-08, 6.319667e-08, 6.315525e-08, 6.346473e-08, 6.329849e-08, 
    6.377079e-08, 6.394317e-08, 6.443005e-08, 6.472857e-08, 6.503251e-08, 
    6.51667e-08, 6.520754e-08, 6.522462e-08 ;

 HR_vr =
  2.705586e-07, 2.712941e-07, 2.711512e-07, 2.717439e-07, 2.714153e-07, 
    2.718033e-07, 2.707078e-07, 2.713232e-07, 2.709305e-07, 2.70625e-07, 
    2.728924e-07, 2.717704e-07, 2.740571e-07, 2.733427e-07, 2.751362e-07, 
    2.739459e-07, 2.75376e-07, 2.751021e-07, 2.759267e-07, 2.756906e-07, 
    2.767435e-07, 2.760356e-07, 2.772891e-07, 2.765747e-07, 2.766864e-07, 
    2.760122e-07, 2.719966e-07, 2.727528e-07, 2.719517e-07, 2.720596e-07, 
    2.720112e-07, 2.71422e-07, 2.711247e-07, 2.705025e-07, 2.706155e-07, 
    2.710726e-07, 2.721081e-07, 2.71757e-07, 2.726422e-07, 2.726222e-07, 
    2.736062e-07, 2.731627e-07, 2.748147e-07, 2.743456e-07, 2.757004e-07, 
    2.753599e-07, 2.756844e-07, 2.75586e-07, 2.756857e-07, 2.751862e-07, 
    2.754003e-07, 2.749607e-07, 2.732457e-07, 2.737501e-07, 2.722446e-07, 
    2.713374e-07, 2.707348e-07, 2.703067e-07, 2.703673e-07, 2.704826e-07, 
    2.710753e-07, 2.716323e-07, 2.720565e-07, 2.7234e-07, 2.726193e-07, 
    2.734634e-07, 2.739102e-07, 2.749094e-07, 2.747294e-07, 2.750345e-07, 
    2.753261e-07, 2.75815e-07, 2.757346e-07, 2.759499e-07, 2.750266e-07, 
    2.756403e-07, 2.746268e-07, 2.749041e-07, 2.726944e-07, 2.718517e-07, 
    2.714926e-07, 2.711787e-07, 2.704138e-07, 2.70942e-07, 2.707338e-07, 
    2.712293e-07, 2.715438e-07, 2.713883e-07, 2.723478e-07, 2.719748e-07, 
    2.739367e-07, 2.730924e-07, 2.752921e-07, 2.747664e-07, 2.75418e-07, 
    2.750856e-07, 2.75655e-07, 2.751426e-07, 2.760301e-07, 2.762231e-07, 
    2.760912e-07, 2.76598e-07, 2.751142e-07, 2.756843e-07, 2.713839e-07, 
    2.714092e-07, 2.715275e-07, 2.710076e-07, 2.709758e-07, 2.704993e-07, 
    2.709234e-07, 2.711039e-07, 2.715621e-07, 2.718328e-07, 2.720901e-07, 
    2.726556e-07, 2.732864e-07, 2.741678e-07, 2.748004e-07, 2.752242e-07, 
    2.749644e-07, 2.751937e-07, 2.749374e-07, 2.748172e-07, 2.761507e-07, 
    2.754022e-07, 2.765251e-07, 2.764631e-07, 2.75955e-07, 2.764701e-07, 
    2.71427e-07, 2.712811e-07, 2.707738e-07, 2.711708e-07, 2.704474e-07, 
    2.708523e-07, 2.71085e-07, 2.719825e-07, 2.721797e-07, 2.723623e-07, 
    2.727229e-07, 2.731854e-07, 2.739959e-07, 2.747004e-07, 2.753431e-07, 
    2.75296e-07, 2.753126e-07, 2.75456e-07, 2.751006e-07, 2.755143e-07, 
    2.755836e-07, 2.754022e-07, 2.764548e-07, 2.761543e-07, 2.764618e-07, 
    2.762661e-07, 2.713286e-07, 2.715742e-07, 2.714415e-07, 2.71691e-07, 
    2.715151e-07, 2.722964e-07, 2.725305e-07, 2.73625e-07, 2.731763e-07, 
    2.738906e-07, 2.732489e-07, 2.733626e-07, 2.739135e-07, 2.732837e-07, 
    2.746614e-07, 2.737273e-07, 2.754615e-07, 2.745295e-07, 2.755199e-07, 
    2.753403e-07, 2.756377e-07, 2.759039e-07, 2.762387e-07, 2.768558e-07, 
    2.76713e-07, 2.772289e-07, 2.719403e-07, 2.722584e-07, 2.722306e-07, 
    2.725636e-07, 2.728097e-07, 2.73343e-07, 2.741974e-07, 2.738763e-07, 
    2.744659e-07, 2.745841e-07, 2.736885e-07, 2.742383e-07, 2.724715e-07, 
    2.727571e-07, 2.725872e-07, 2.719653e-07, 2.739501e-07, 2.729321e-07, 
    2.748109e-07, 2.742603e-07, 2.758659e-07, 2.750677e-07, 2.766344e-07, 
    2.773025e-07, 2.779315e-07, 2.786648e-07, 2.724322e-07, 2.722161e-07, 
    2.726032e-07, 2.731382e-07, 2.736346e-07, 2.742939e-07, 2.743614e-07, 
    2.744847e-07, 2.748044e-07, 2.750729e-07, 2.745236e-07, 2.751403e-07, 
    2.72823e-07, 2.740385e-07, 2.721342e-07, 2.727079e-07, 2.731067e-07, 
    2.72932e-07, 2.738396e-07, 2.740533e-07, 2.74921e-07, 2.744727e-07, 
    2.771375e-07, 2.759598e-07, 2.792231e-07, 2.783128e-07, 2.721405e-07, 
    2.724316e-07, 2.734434e-07, 2.729622e-07, 2.743379e-07, 2.746761e-07, 
    2.74951e-07, 2.753019e-07, 2.753399e-07, 2.755478e-07, 2.752071e-07, 
    2.755344e-07, 2.742953e-07, 2.748493e-07, 2.73328e-07, 2.736985e-07, 
    2.735281e-07, 2.733411e-07, 2.739182e-07, 2.745322e-07, 2.745456e-07, 
    2.747423e-07, 2.752958e-07, 2.743435e-07, 2.772889e-07, 2.75471e-07, 
    2.727488e-07, 2.733085e-07, 2.733887e-07, 2.731719e-07, 2.746422e-07, 
    2.741098e-07, 2.755428e-07, 2.751559e-07, 2.757898e-07, 2.754748e-07, 
    2.754285e-07, 2.750238e-07, 2.747716e-07, 2.741342e-07, 2.736151e-07, 
    2.732034e-07, 2.732992e-07, 2.737514e-07, 2.745698e-07, 2.753433e-07, 
    2.751739e-07, 2.757417e-07, 2.742383e-07, 2.748689e-07, 2.746252e-07, 
    2.752606e-07, 2.738677e-07, 2.750533e-07, 2.735642e-07, 2.73695e-07, 
    2.740992e-07, 2.749115e-07, 2.750915e-07, 2.752831e-07, 2.751649e-07, 
    2.745906e-07, 2.744966e-07, 2.740895e-07, 2.739769e-07, 2.736665e-07, 
    2.734094e-07, 2.736443e-07, 2.738908e-07, 2.745909e-07, 2.752211e-07, 
    2.759076e-07, 2.760756e-07, 2.768759e-07, 2.762241e-07, 2.772989e-07, 
    2.763847e-07, 2.779667e-07, 2.751223e-07, 2.763583e-07, 2.741177e-07, 
    2.743595e-07, 2.747964e-07, 2.757979e-07, 2.752577e-07, 2.758895e-07, 
    2.744929e-07, 2.737669e-07, 2.735792e-07, 2.732284e-07, 2.735872e-07, 
    2.73558e-07, 2.739012e-07, 2.73791e-07, 2.746142e-07, 2.741721e-07, 
    2.754273e-07, 2.758846e-07, 2.771748e-07, 2.779643e-07, 2.787673e-07, 
    2.791214e-07, 2.792291e-07, 2.792742e-07,
  2.344915e-07, 2.353864e-07, 2.352125e-07, 2.359338e-07, 2.355338e-07, 
    2.36006e-07, 2.34673e-07, 2.354218e-07, 2.349439e-07, 2.345722e-07, 
    2.37332e-07, 2.35966e-07, 2.387497e-07, 2.378798e-07, 2.400639e-07, 
    2.386143e-07, 2.40356e-07, 2.400223e-07, 2.410267e-07, 2.40739e-07, 
    2.420222e-07, 2.411594e-07, 2.42687e-07, 2.418163e-07, 2.419525e-07, 
    2.411309e-07, 2.362412e-07, 2.37162e-07, 2.361866e-07, 2.363179e-07, 
    2.36259e-07, 2.35542e-07, 2.351804e-07, 2.344231e-07, 2.345607e-07, 
    2.351169e-07, 2.36377e-07, 2.359495e-07, 2.370269e-07, 2.370026e-07, 
    2.382006e-07, 2.376606e-07, 2.396722e-07, 2.391009e-07, 2.407511e-07, 
    2.403363e-07, 2.407315e-07, 2.406117e-07, 2.407331e-07, 2.401248e-07, 
    2.403854e-07, 2.3985e-07, 2.377617e-07, 2.383758e-07, 2.36543e-07, 
    2.354392e-07, 2.347059e-07, 2.34185e-07, 2.342586e-07, 2.34399e-07, 
    2.351202e-07, 2.357979e-07, 2.36314e-07, 2.366591e-07, 2.369991e-07, 
    2.380269e-07, 2.385709e-07, 2.397876e-07, 2.395683e-07, 2.399399e-07, 
    2.40295e-07, 2.408907e-07, 2.407928e-07, 2.410551e-07, 2.399302e-07, 
    2.406779e-07, 2.394433e-07, 2.397811e-07, 2.370909e-07, 2.360649e-07, 
    2.35628e-07, 2.352459e-07, 2.343153e-07, 2.34958e-07, 2.347047e-07, 
    2.353074e-07, 2.356901e-07, 2.355009e-07, 2.366686e-07, 2.362147e-07, 
    2.386031e-07, 2.375751e-07, 2.402536e-07, 2.396133e-07, 2.40407e-07, 
    2.400022e-07, 2.406958e-07, 2.400716e-07, 2.411527e-07, 2.413879e-07, 
    2.412272e-07, 2.418447e-07, 2.400369e-07, 2.407315e-07, 2.354955e-07, 
    2.355264e-07, 2.356703e-07, 2.350378e-07, 2.349991e-07, 2.344193e-07, 
    2.349353e-07, 2.351549e-07, 2.357124e-07, 2.360419e-07, 2.36355e-07, 
    2.370433e-07, 2.378113e-07, 2.388845e-07, 2.396548e-07, 2.401709e-07, 
    2.398545e-07, 2.401338e-07, 2.398216e-07, 2.396752e-07, 2.412998e-07, 
    2.403878e-07, 2.417559e-07, 2.416803e-07, 2.410613e-07, 2.416888e-07, 
    2.355481e-07, 2.353705e-07, 2.347533e-07, 2.352363e-07, 2.343562e-07, 
    2.348489e-07, 2.35132e-07, 2.362241e-07, 2.36464e-07, 2.366863e-07, 
    2.371252e-07, 2.376882e-07, 2.386751e-07, 2.395331e-07, 2.403157e-07, 
    2.402584e-07, 2.402786e-07, 2.404533e-07, 2.400204e-07, 2.405243e-07, 
    2.406088e-07, 2.403878e-07, 2.416701e-07, 2.41304e-07, 2.416787e-07, 
    2.414403e-07, 2.354282e-07, 2.357271e-07, 2.355656e-07, 2.358693e-07, 
    2.356553e-07, 2.366062e-07, 2.368912e-07, 2.382236e-07, 2.376771e-07, 
    2.385469e-07, 2.377656e-07, 2.37904e-07, 2.38575e-07, 2.378078e-07, 
    2.394856e-07, 2.383482e-07, 2.404601e-07, 2.393251e-07, 2.405311e-07, 
    2.403123e-07, 2.406746e-07, 2.409989e-07, 2.414069e-07, 2.42159e-07, 
    2.419849e-07, 2.426136e-07, 2.361726e-07, 2.3656e-07, 2.36526e-07, 
    2.369313e-07, 2.372309e-07, 2.378801e-07, 2.389204e-07, 2.385294e-07, 
    2.392473e-07, 2.393913e-07, 2.383007e-07, 2.389704e-07, 2.368192e-07, 
    2.371669e-07, 2.3696e-07, 2.362031e-07, 2.386194e-07, 2.3738e-07, 
    2.396675e-07, 2.38997e-07, 2.409527e-07, 2.399805e-07, 2.41889e-07, 
    2.427035e-07, 2.434699e-07, 2.443641e-07, 2.367714e-07, 2.365083e-07, 
    2.369795e-07, 2.376309e-07, 2.382352e-07, 2.390379e-07, 2.391201e-07, 
    2.392703e-07, 2.396596e-07, 2.399867e-07, 2.393177e-07, 2.400687e-07, 
    2.372473e-07, 2.387269e-07, 2.364087e-07, 2.371071e-07, 2.375925e-07, 
    2.373798e-07, 2.384847e-07, 2.387449e-07, 2.398017e-07, 2.392556e-07, 
    2.425024e-07, 2.410673e-07, 2.450448e-07, 2.439349e-07, 2.364163e-07, 
    2.367706e-07, 2.380024e-07, 2.374165e-07, 2.390915e-07, 2.395034e-07, 
    2.398381e-07, 2.402657e-07, 2.403119e-07, 2.405652e-07, 2.401502e-07, 
    2.405489e-07, 2.390396e-07, 2.397144e-07, 2.378618e-07, 2.38313e-07, 
    2.381055e-07, 2.378778e-07, 2.385804e-07, 2.393282e-07, 2.393444e-07, 
    2.39584e-07, 2.402587e-07, 2.390983e-07, 2.426872e-07, 2.40472e-07, 
    2.371567e-07, 2.378383e-07, 2.379358e-07, 2.376718e-07, 2.394621e-07, 
    2.388138e-07, 2.405591e-07, 2.400877e-07, 2.408599e-07, 2.404763e-07, 
    2.404198e-07, 2.399268e-07, 2.396197e-07, 2.388435e-07, 2.382115e-07, 
    2.377101e-07, 2.378267e-07, 2.383774e-07, 2.39374e-07, 2.403161e-07, 
    2.401098e-07, 2.408013e-07, 2.389702e-07, 2.397383e-07, 2.394414e-07, 
    2.402154e-07, 2.38519e-07, 2.399632e-07, 2.381494e-07, 2.383086e-07, 
    2.388009e-07, 2.397903e-07, 2.400093e-07, 2.402428e-07, 2.400988e-07, 
    2.393993e-07, 2.392848e-07, 2.38789e-07, 2.386519e-07, 2.38274e-07, 
    2.379609e-07, 2.382469e-07, 2.385472e-07, 2.393997e-07, 2.401673e-07, 
    2.410035e-07, 2.412081e-07, 2.421836e-07, 2.413894e-07, 2.426994e-07, 
    2.415854e-07, 2.435133e-07, 2.400471e-07, 2.415529e-07, 2.388233e-07, 
    2.391178e-07, 2.3965e-07, 2.4087e-07, 2.402117e-07, 2.409816e-07, 
    2.392803e-07, 2.383963e-07, 2.381676e-07, 2.377406e-07, 2.381774e-07, 
    2.381419e-07, 2.385597e-07, 2.384255e-07, 2.39428e-07, 2.388896e-07, 
    2.404183e-07, 2.409756e-07, 2.425477e-07, 2.4351e-07, 2.44489e-07, 
    2.449207e-07, 2.450521e-07, 2.45107e-07,
  2.19386e-07, 2.203636e-07, 2.201737e-07, 2.209618e-07, 2.205247e-07, 
    2.210407e-07, 2.195843e-07, 2.204024e-07, 2.198802e-07, 2.194741e-07, 
    2.224903e-07, 2.20997e-07, 2.240406e-07, 2.230892e-07, 2.254785e-07, 
    2.238926e-07, 2.257981e-07, 2.254329e-07, 2.265322e-07, 2.262174e-07, 
    2.276225e-07, 2.266776e-07, 2.283505e-07, 2.273969e-07, 2.275461e-07, 
    2.266463e-07, 2.212978e-07, 2.223044e-07, 2.212381e-07, 2.213817e-07, 
    2.213172e-07, 2.205337e-07, 2.201386e-07, 2.193113e-07, 2.194616e-07, 
    2.200692e-07, 2.214462e-07, 2.20979e-07, 2.221565e-07, 2.2213e-07, 
    2.234399e-07, 2.228494e-07, 2.250498e-07, 2.244247e-07, 2.262305e-07, 
    2.257766e-07, 2.262092e-07, 2.26078e-07, 2.262109e-07, 2.255451e-07, 
    2.258303e-07, 2.252444e-07, 2.2296e-07, 2.236316e-07, 2.216277e-07, 
    2.204215e-07, 2.196202e-07, 2.190512e-07, 2.191317e-07, 2.19285e-07, 
    2.200728e-07, 2.208133e-07, 2.213773e-07, 2.217545e-07, 2.221261e-07, 
    2.232502e-07, 2.23845e-07, 2.251761e-07, 2.249361e-07, 2.253428e-07, 
    2.257314e-07, 2.263835e-07, 2.262762e-07, 2.265634e-07, 2.253321e-07, 
    2.261505e-07, 2.247993e-07, 2.25169e-07, 2.222267e-07, 2.211051e-07, 
    2.206278e-07, 2.202102e-07, 2.191935e-07, 2.198956e-07, 2.196189e-07, 
    2.202773e-07, 2.206955e-07, 2.204887e-07, 2.217649e-07, 2.212688e-07, 
    2.238803e-07, 2.227559e-07, 2.256861e-07, 2.249854e-07, 2.25854e-07, 
    2.254108e-07, 2.261701e-07, 2.254868e-07, 2.266703e-07, 2.269278e-07, 
    2.267518e-07, 2.274279e-07, 2.254489e-07, 2.262091e-07, 2.204829e-07, 
    2.205166e-07, 2.206738e-07, 2.199828e-07, 2.199405e-07, 2.193072e-07, 
    2.198708e-07, 2.201107e-07, 2.207198e-07, 2.210799e-07, 2.214222e-07, 
    2.221745e-07, 2.230143e-07, 2.24188e-07, 2.250308e-07, 2.255955e-07, 
    2.252493e-07, 2.255549e-07, 2.252132e-07, 2.250531e-07, 2.268313e-07, 
    2.25833e-07, 2.273307e-07, 2.272479e-07, 2.265702e-07, 2.272572e-07, 
    2.205403e-07, 2.203462e-07, 2.19672e-07, 2.201996e-07, 2.192382e-07, 
    2.197764e-07, 2.200857e-07, 2.212791e-07, 2.215413e-07, 2.217842e-07, 
    2.222641e-07, 2.228796e-07, 2.23959e-07, 2.248975e-07, 2.25754e-07, 
    2.256913e-07, 2.257134e-07, 2.259046e-07, 2.254308e-07, 2.259824e-07, 
    2.260749e-07, 2.258329e-07, 2.272368e-07, 2.268359e-07, 2.272461e-07, 
    2.269851e-07, 2.204093e-07, 2.207359e-07, 2.205594e-07, 2.208913e-07, 
    2.206575e-07, 2.216968e-07, 2.220083e-07, 2.234652e-07, 2.228675e-07, 
    2.238187e-07, 2.229642e-07, 2.231156e-07, 2.238496e-07, 2.230104e-07, 
    2.248457e-07, 2.236015e-07, 2.25912e-07, 2.246701e-07, 2.259898e-07, 
    2.257503e-07, 2.261469e-07, 2.265019e-07, 2.269485e-07, 2.277722e-07, 
    2.275815e-07, 2.282702e-07, 2.212228e-07, 2.216462e-07, 2.21609e-07, 
    2.22052e-07, 2.223796e-07, 2.230895e-07, 2.242273e-07, 2.237995e-07, 
    2.245849e-07, 2.247425e-07, 2.235494e-07, 2.242819e-07, 2.219295e-07, 
    2.223097e-07, 2.220834e-07, 2.212561e-07, 2.23898e-07, 2.225427e-07, 
    2.250447e-07, 2.243111e-07, 2.264513e-07, 2.253872e-07, 2.274765e-07, 
    2.283687e-07, 2.292083e-07, 2.301884e-07, 2.218773e-07, 2.215896e-07, 
    2.221047e-07, 2.22817e-07, 2.234778e-07, 2.243558e-07, 2.244457e-07, 
    2.246101e-07, 2.25036e-07, 2.253939e-07, 2.24662e-07, 2.254837e-07, 
    2.223978e-07, 2.240157e-07, 2.214808e-07, 2.222444e-07, 2.22775e-07, 
    2.225423e-07, 2.237507e-07, 2.240353e-07, 2.251915e-07, 2.245939e-07, 
    2.281485e-07, 2.265768e-07, 2.309346e-07, 2.297179e-07, 2.214891e-07, 
    2.218763e-07, 2.232233e-07, 2.225825e-07, 2.244145e-07, 2.248651e-07, 
    2.252313e-07, 2.256993e-07, 2.257499e-07, 2.260271e-07, 2.255728e-07, 
    2.260092e-07, 2.243577e-07, 2.250959e-07, 2.230694e-07, 2.235628e-07, 
    2.233359e-07, 2.230869e-07, 2.238553e-07, 2.246735e-07, 2.246911e-07, 
    2.249534e-07, 2.256919e-07, 2.244219e-07, 2.28351e-07, 2.259254e-07, 
    2.222985e-07, 2.230438e-07, 2.231503e-07, 2.228617e-07, 2.248199e-07, 
    2.241106e-07, 2.260204e-07, 2.255045e-07, 2.263497e-07, 2.259298e-07, 
    2.258679e-07, 2.253284e-07, 2.249923e-07, 2.241431e-07, 2.234518e-07, 
    2.229036e-07, 2.230311e-07, 2.236333e-07, 2.247236e-07, 2.257544e-07, 
    2.255287e-07, 2.262855e-07, 2.242817e-07, 2.251222e-07, 2.247973e-07, 
    2.256442e-07, 2.237882e-07, 2.253684e-07, 2.233839e-07, 2.23558e-07, 
    2.240965e-07, 2.251791e-07, 2.254187e-07, 2.256742e-07, 2.255165e-07, 
    2.247513e-07, 2.246259e-07, 2.240835e-07, 2.239336e-07, 2.235202e-07, 
    2.231777e-07, 2.234906e-07, 2.23819e-07, 2.247516e-07, 2.255916e-07, 
    2.265069e-07, 2.267309e-07, 2.277993e-07, 2.269295e-07, 2.283645e-07, 
    2.271443e-07, 2.29256e-07, 2.254602e-07, 2.271086e-07, 2.241211e-07, 
    2.244432e-07, 2.250256e-07, 2.263608e-07, 2.256402e-07, 2.26483e-07, 
    2.24621e-07, 2.23654e-07, 2.234039e-07, 2.229369e-07, 2.234145e-07, 
    2.233757e-07, 2.238327e-07, 2.236859e-07, 2.247826e-07, 2.241936e-07, 
    2.258664e-07, 2.264764e-07, 2.28198e-07, 2.292524e-07, 2.303252e-07, 
    2.307985e-07, 2.309425e-07, 2.310027e-07,
  2.09813e-07, 2.108176e-07, 2.106223e-07, 2.114325e-07, 2.109831e-07, 
    2.115136e-07, 2.100167e-07, 2.108574e-07, 2.103207e-07, 2.099035e-07, 
    2.130047e-07, 2.114687e-07, 2.146002e-07, 2.136207e-07, 2.160814e-07, 
    2.144478e-07, 2.164108e-07, 2.160343e-07, 2.171674e-07, 2.168428e-07, 
    2.18292e-07, 2.173173e-07, 2.190432e-07, 2.180592e-07, 2.182131e-07, 
    2.172851e-07, 2.117778e-07, 2.128134e-07, 2.117164e-07, 2.118641e-07, 
    2.117979e-07, 2.109924e-07, 2.105864e-07, 2.097363e-07, 2.098906e-07, 
    2.10515e-07, 2.119305e-07, 2.114501e-07, 2.12661e-07, 2.126337e-07, 
    2.139817e-07, 2.133739e-07, 2.156396e-07, 2.149957e-07, 2.168564e-07, 
    2.163884e-07, 2.168344e-07, 2.166992e-07, 2.168361e-07, 2.161499e-07, 
    2.164439e-07, 2.1584e-07, 2.134878e-07, 2.141791e-07, 2.121171e-07, 
    2.108771e-07, 2.100536e-07, 2.094691e-07, 2.095517e-07, 2.097092e-07, 
    2.105187e-07, 2.112797e-07, 2.118596e-07, 2.122475e-07, 2.126298e-07, 
    2.137865e-07, 2.143989e-07, 2.157698e-07, 2.155224e-07, 2.159415e-07, 
    2.163419e-07, 2.17014e-07, 2.169034e-07, 2.171995e-07, 2.159305e-07, 
    2.167739e-07, 2.153815e-07, 2.157623e-07, 2.127335e-07, 2.115797e-07, 
    2.110891e-07, 2.106598e-07, 2.096153e-07, 2.103366e-07, 2.100522e-07, 
    2.107288e-07, 2.111586e-07, 2.109461e-07, 2.122581e-07, 2.11748e-07, 
    2.144351e-07, 2.132778e-07, 2.162952e-07, 2.155732e-07, 2.164682e-07, 
    2.160115e-07, 2.167941e-07, 2.160898e-07, 2.173098e-07, 2.175754e-07, 
    2.173939e-07, 2.180912e-07, 2.160508e-07, 2.168344e-07, 2.109401e-07, 
    2.109748e-07, 2.111363e-07, 2.104262e-07, 2.103827e-07, 2.09732e-07, 
    2.103111e-07, 2.105576e-07, 2.111836e-07, 2.115538e-07, 2.119057e-07, 
    2.126795e-07, 2.135436e-07, 2.147519e-07, 2.1562e-07, 2.162018e-07, 
    2.158451e-07, 2.1616e-07, 2.158079e-07, 2.156429e-07, 2.174758e-07, 
    2.164467e-07, 2.179909e-07, 2.179055e-07, 2.172066e-07, 2.179151e-07, 
    2.109991e-07, 2.107996e-07, 2.101068e-07, 2.10649e-07, 2.096612e-07, 
    2.102141e-07, 2.10532e-07, 2.117587e-07, 2.120282e-07, 2.122781e-07, 
    2.127717e-07, 2.13405e-07, 2.145161e-07, 2.154827e-07, 2.163652e-07, 
    2.163005e-07, 2.163233e-07, 2.165204e-07, 2.160321e-07, 2.166006e-07, 
    2.16696e-07, 2.164465e-07, 2.17894e-07, 2.174805e-07, 2.179036e-07, 
    2.176344e-07, 2.108644e-07, 2.112002e-07, 2.110188e-07, 2.113599e-07, 
    2.111196e-07, 2.121882e-07, 2.125086e-07, 2.140078e-07, 2.133926e-07, 
    2.143717e-07, 2.13492e-07, 2.136479e-07, 2.144036e-07, 2.135396e-07, 
    2.154294e-07, 2.141482e-07, 2.165281e-07, 2.152486e-07, 2.166082e-07, 
    2.163614e-07, 2.167701e-07, 2.171362e-07, 2.175967e-07, 2.184464e-07, 
    2.182496e-07, 2.189602e-07, 2.117007e-07, 2.121361e-07, 2.120978e-07, 
    2.125535e-07, 2.128905e-07, 2.13621e-07, 2.147924e-07, 2.143519e-07, 
    2.151606e-07, 2.15323e-07, 2.140944e-07, 2.148487e-07, 2.124276e-07, 
    2.128187e-07, 2.125858e-07, 2.11735e-07, 2.144534e-07, 2.130584e-07, 
    2.156343e-07, 2.148787e-07, 2.17084e-07, 2.159873e-07, 2.181413e-07, 
    2.19062e-07, 2.199286e-07, 2.209411e-07, 2.123738e-07, 2.120779e-07, 
    2.126077e-07, 2.133406e-07, 2.140207e-07, 2.149247e-07, 2.150173e-07, 
    2.151866e-07, 2.156253e-07, 2.159941e-07, 2.152401e-07, 2.160866e-07, 
    2.129094e-07, 2.145745e-07, 2.119661e-07, 2.127515e-07, 2.132974e-07, 
    2.13058e-07, 2.143016e-07, 2.145947e-07, 2.157856e-07, 2.1517e-07, 
    2.188347e-07, 2.172135e-07, 2.21712e-07, 2.20455e-07, 2.119746e-07, 
    2.123728e-07, 2.137587e-07, 2.130993e-07, 2.149851e-07, 2.154493e-07, 
    2.158266e-07, 2.163089e-07, 2.16361e-07, 2.166467e-07, 2.161785e-07, 
    2.166282e-07, 2.149267e-07, 2.156871e-07, 2.136003e-07, 2.141082e-07, 
    2.138746e-07, 2.136183e-07, 2.144093e-07, 2.15252e-07, 2.1527e-07, 
    2.155402e-07, 2.163015e-07, 2.149928e-07, 2.190439e-07, 2.165421e-07, 
    2.128071e-07, 2.13574e-07, 2.136836e-07, 2.133865e-07, 2.154027e-07, 
    2.146722e-07, 2.166397e-07, 2.16108e-07, 2.169792e-07, 2.165463e-07, 
    2.164826e-07, 2.159266e-07, 2.155804e-07, 2.147057e-07, 2.13994e-07, 
    2.134296e-07, 2.135609e-07, 2.141808e-07, 2.153036e-07, 2.163657e-07, 
    2.16133e-07, 2.16913e-07, 2.148484e-07, 2.157142e-07, 2.153795e-07, 
    2.16252e-07, 2.143402e-07, 2.159681e-07, 2.139241e-07, 2.141033e-07, 
    2.146577e-07, 2.157728e-07, 2.160196e-07, 2.16283e-07, 2.161205e-07, 
    2.153321e-07, 2.152029e-07, 2.146442e-07, 2.1449e-07, 2.140643e-07, 
    2.137118e-07, 2.140338e-07, 2.14372e-07, 2.153324e-07, 2.161979e-07, 
    2.171414e-07, 2.173723e-07, 2.184745e-07, 2.175772e-07, 2.190578e-07, 
    2.17799e-07, 2.199781e-07, 2.160625e-07, 2.17762e-07, 2.14683e-07, 
    2.150147e-07, 2.156147e-07, 2.169908e-07, 2.162479e-07, 2.171167e-07, 
    2.151978e-07, 2.142022e-07, 2.139446e-07, 2.134639e-07, 2.139556e-07, 
    2.139156e-07, 2.14386e-07, 2.142349e-07, 2.153643e-07, 2.147576e-07, 
    2.16481e-07, 2.171099e-07, 2.188857e-07, 2.199742e-07, 2.210822e-07, 
    2.215713e-07, 2.217202e-07, 2.217824e-07,
  2.025419e-07, 2.034944e-07, 2.033092e-07, 2.040779e-07, 2.036514e-07, 
    2.041549e-07, 2.02735e-07, 2.035323e-07, 2.030232e-07, 2.026276e-07, 
    2.055712e-07, 2.041122e-07, 2.070885e-07, 2.061566e-07, 2.08499e-07, 
    2.069435e-07, 2.088129e-07, 2.084541e-07, 2.095343e-07, 2.092247e-07, 
    2.106076e-07, 2.096772e-07, 2.113251e-07, 2.103854e-07, 2.105323e-07, 
    2.096466e-07, 2.044057e-07, 2.053895e-07, 2.043474e-07, 2.044876e-07, 
    2.044247e-07, 2.036602e-07, 2.032752e-07, 2.024691e-07, 2.026154e-07, 
    2.032075e-07, 2.045507e-07, 2.040945e-07, 2.052445e-07, 2.052185e-07, 
    2.065e-07, 2.05922e-07, 2.08078e-07, 2.074648e-07, 2.092377e-07, 
    2.087916e-07, 2.092167e-07, 2.090878e-07, 2.092184e-07, 2.085642e-07, 
    2.088444e-07, 2.082689e-07, 2.060302e-07, 2.066877e-07, 2.047278e-07, 
    2.03551e-07, 2.027699e-07, 2.02216e-07, 2.022943e-07, 2.024435e-07, 
    2.032109e-07, 2.039329e-07, 2.044833e-07, 2.048517e-07, 2.052147e-07, 
    2.063144e-07, 2.068969e-07, 2.082021e-07, 2.079664e-07, 2.083656e-07, 
    2.087472e-07, 2.09388e-07, 2.092825e-07, 2.09565e-07, 2.083551e-07, 
    2.091591e-07, 2.078322e-07, 2.081949e-07, 2.053136e-07, 2.042176e-07, 
    2.037521e-07, 2.033448e-07, 2.023545e-07, 2.030383e-07, 2.027687e-07, 
    2.034102e-07, 2.03818e-07, 2.036163e-07, 2.048617e-07, 2.043774e-07, 
    2.069314e-07, 2.058306e-07, 2.087027e-07, 2.080148e-07, 2.088676e-07, 
    2.084323e-07, 2.091783e-07, 2.085069e-07, 2.096701e-07, 2.099236e-07, 
    2.097504e-07, 2.104158e-07, 2.084697e-07, 2.092167e-07, 2.036106e-07, 
    2.036435e-07, 2.037968e-07, 2.031232e-07, 2.03082e-07, 2.024651e-07, 
    2.03014e-07, 2.032479e-07, 2.038416e-07, 2.04193e-07, 2.045271e-07, 
    2.05262e-07, 2.060834e-07, 2.072328e-07, 2.080593e-07, 2.086137e-07, 
    2.082737e-07, 2.085739e-07, 2.082384e-07, 2.080811e-07, 2.098286e-07, 
    2.088471e-07, 2.103201e-07, 2.102385e-07, 2.095717e-07, 2.102477e-07, 
    2.036666e-07, 2.034773e-07, 2.028204e-07, 2.033345e-07, 2.023979e-07, 
    2.029221e-07, 2.032236e-07, 2.043875e-07, 2.046434e-07, 2.048807e-07, 
    2.053496e-07, 2.059516e-07, 2.070084e-07, 2.079286e-07, 2.087694e-07, 
    2.087077e-07, 2.087294e-07, 2.089174e-07, 2.08452e-07, 2.089938e-07, 
    2.090847e-07, 2.088469e-07, 2.102276e-07, 2.09833e-07, 2.102368e-07, 
    2.099798e-07, 2.035389e-07, 2.038574e-07, 2.036853e-07, 2.04009e-07, 
    2.037809e-07, 2.047954e-07, 2.050998e-07, 2.065248e-07, 2.059397e-07, 
    2.06871e-07, 2.060343e-07, 2.061825e-07, 2.069014e-07, 2.060795e-07, 
    2.078779e-07, 2.066584e-07, 2.089246e-07, 2.077058e-07, 2.090011e-07, 
    2.087657e-07, 2.091554e-07, 2.095045e-07, 2.099439e-07, 2.10755e-07, 
    2.105671e-07, 2.112458e-07, 2.043325e-07, 2.047459e-07, 2.047095e-07, 
    2.051423e-07, 2.054625e-07, 2.061569e-07, 2.072713e-07, 2.068521e-07, 
    2.076218e-07, 2.077764e-07, 2.066071e-07, 2.073249e-07, 2.050227e-07, 
    2.053944e-07, 2.051731e-07, 2.043651e-07, 2.069487e-07, 2.056221e-07, 
    2.08073e-07, 2.073534e-07, 2.094547e-07, 2.084093e-07, 2.104637e-07, 
    2.113432e-07, 2.121714e-07, 2.131403e-07, 2.049716e-07, 2.046906e-07, 
    2.051938e-07, 2.058904e-07, 2.06537e-07, 2.073973e-07, 2.074854e-07, 
    2.076466e-07, 2.080644e-07, 2.084158e-07, 2.076976e-07, 2.085038e-07, 
    2.054806e-07, 2.070639e-07, 2.045844e-07, 2.053305e-07, 2.058493e-07, 
    2.056217e-07, 2.068042e-07, 2.070831e-07, 2.082171e-07, 2.076307e-07, 
    2.111261e-07, 2.095783e-07, 2.138784e-07, 2.126751e-07, 2.045925e-07, 
    2.049706e-07, 2.062879e-07, 2.05661e-07, 2.074547e-07, 2.078967e-07, 
    2.082561e-07, 2.087157e-07, 2.087654e-07, 2.090378e-07, 2.085914e-07, 
    2.090201e-07, 2.073991e-07, 2.081232e-07, 2.061372e-07, 2.066203e-07, 
    2.06398e-07, 2.061543e-07, 2.069067e-07, 2.077089e-07, 2.07726e-07, 
    2.079834e-07, 2.087089e-07, 2.07462e-07, 2.11326e-07, 2.089382e-07, 
    2.053832e-07, 2.061123e-07, 2.062165e-07, 2.05934e-07, 2.078524e-07, 
    2.071569e-07, 2.090311e-07, 2.085243e-07, 2.093548e-07, 2.089421e-07, 
    2.088813e-07, 2.083514e-07, 2.080216e-07, 2.071888e-07, 2.065116e-07, 
    2.059749e-07, 2.060997e-07, 2.066893e-07, 2.07758e-07, 2.087699e-07, 
    2.085481e-07, 2.092917e-07, 2.073246e-07, 2.08149e-07, 2.078304e-07, 
    2.086615e-07, 2.06841e-07, 2.083912e-07, 2.064451e-07, 2.066156e-07, 
    2.071431e-07, 2.08205e-07, 2.0844e-07, 2.086911e-07, 2.085362e-07, 
    2.077851e-07, 2.076621e-07, 2.071303e-07, 2.069835e-07, 2.065784e-07, 
    2.062432e-07, 2.065495e-07, 2.068713e-07, 2.077854e-07, 2.086099e-07, 
    2.095095e-07, 2.097298e-07, 2.10782e-07, 2.099254e-07, 2.113394e-07, 
    2.101372e-07, 2.12219e-07, 2.084811e-07, 2.101018e-07, 2.071671e-07, 
    2.074829e-07, 2.080543e-07, 2.093659e-07, 2.086576e-07, 2.09486e-07, 
    2.076573e-07, 2.067097e-07, 2.064646e-07, 2.060076e-07, 2.064751e-07, 
    2.06437e-07, 2.068846e-07, 2.067407e-07, 2.078158e-07, 2.072382e-07, 
    2.088798e-07, 2.094795e-07, 2.111747e-07, 2.122151e-07, 2.132753e-07, 
    2.137436e-07, 2.138862e-07, 2.139458e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.194416e-08, 6.221921e-08, 6.216575e-08, 6.238761e-08, 6.226454e-08, 
    6.240981e-08, 6.199993e-08, 6.223013e-08, 6.208317e-08, 6.196893e-08, 
    6.281821e-08, 6.239751e-08, 6.325536e-08, 6.298698e-08, 6.366125e-08, 
    6.321359e-08, 6.375153e-08, 6.364835e-08, 6.395895e-08, 6.386996e-08, 
    6.426725e-08, 6.400002e-08, 6.447324e-08, 6.420344e-08, 6.424563e-08, 
    6.39912e-08, 6.248218e-08, 6.276583e-08, 6.246538e-08, 6.250582e-08, 
    6.248767e-08, 6.226708e-08, 6.215591e-08, 6.192315e-08, 6.19654e-08, 
    6.213637e-08, 6.2524e-08, 6.239242e-08, 6.272409e-08, 6.27166e-08, 
    6.308589e-08, 6.291938e-08, 6.354018e-08, 6.336372e-08, 6.387368e-08, 
    6.374542e-08, 6.386765e-08, 6.383059e-08, 6.386814e-08, 6.368003e-08, 
    6.376062e-08, 6.359511e-08, 6.295056e-08, 6.313996e-08, 6.25751e-08, 
    6.223551e-08, 6.201002e-08, 6.185e-08, 6.187263e-08, 6.191575e-08, 
    6.213737e-08, 6.234576e-08, 6.250459e-08, 6.261083e-08, 6.271553e-08, 
    6.303241e-08, 6.320018e-08, 6.357585e-08, 6.350807e-08, 6.362291e-08, 
    6.373266e-08, 6.39169e-08, 6.388658e-08, 6.396775e-08, 6.361989e-08, 
    6.385107e-08, 6.346945e-08, 6.357381e-08, 6.274394e-08, 6.242792e-08, 
    6.229357e-08, 6.217602e-08, 6.189002e-08, 6.208752e-08, 6.200966e-08, 
    6.219491e-08, 6.231262e-08, 6.22544e-08, 6.261374e-08, 6.247403e-08, 
    6.321012e-08, 6.289304e-08, 6.371985e-08, 6.352198e-08, 6.376729e-08, 
    6.364211e-08, 6.38566e-08, 6.366356e-08, 6.399797e-08, 6.407078e-08, 
    6.402102e-08, 6.421219e-08, 6.365286e-08, 6.386765e-08, 6.225277e-08, 
    6.226226e-08, 6.23065e-08, 6.211204e-08, 6.210015e-08, 6.192198e-08, 
    6.208052e-08, 6.214803e-08, 6.231944e-08, 6.242083e-08, 6.251722e-08, 
    6.272915e-08, 6.296587e-08, 6.329692e-08, 6.353481e-08, 6.369427e-08, 
    6.359649e-08, 6.368282e-08, 6.358631e-08, 6.354109e-08, 6.40435e-08, 
    6.376137e-08, 6.41847e-08, 6.416128e-08, 6.396969e-08, 6.416391e-08, 
    6.226892e-08, 6.221429e-08, 6.202459e-08, 6.217304e-08, 6.190258e-08, 
    6.205396e-08, 6.214101e-08, 6.247694e-08, 6.255076e-08, 6.26192e-08, 
    6.27544e-08, 6.29279e-08, 6.32323e-08, 6.349719e-08, 6.373904e-08, 
    6.372132e-08, 6.372756e-08, 6.378159e-08, 6.364776e-08, 6.380356e-08, 
    6.38297e-08, 6.376134e-08, 6.415814e-08, 6.404477e-08, 6.416078e-08, 
    6.408697e-08, 6.223205e-08, 6.232399e-08, 6.227431e-08, 6.236773e-08, 
    6.230191e-08, 6.259458e-08, 6.268234e-08, 6.309303e-08, 6.292449e-08, 
    6.319274e-08, 6.295173e-08, 6.299444e-08, 6.320148e-08, 6.296477e-08, 
    6.348257e-08, 6.313149e-08, 6.378369e-08, 6.343302e-08, 6.380566e-08, 
    6.3738e-08, 6.385004e-08, 6.395038e-08, 6.407663e-08, 6.430958e-08, 
    6.425564e-08, 6.445048e-08, 6.246106e-08, 6.258032e-08, 6.256982e-08, 
    6.269464e-08, 6.278695e-08, 6.298706e-08, 6.330801e-08, 6.318732e-08, 
    6.340892e-08, 6.345341e-08, 6.311675e-08, 6.332343e-08, 6.266014e-08, 
    6.276728e-08, 6.27035e-08, 6.247047e-08, 6.321512e-08, 6.283292e-08, 
    6.353874e-08, 6.333165e-08, 6.393607e-08, 6.363545e-08, 6.422594e-08, 
    6.447839e-08, 6.471606e-08, 6.499378e-08, 6.264541e-08, 6.256438e-08, 
    6.270949e-08, 6.291025e-08, 6.309657e-08, 6.334428e-08, 6.336963e-08, 
    6.341604e-08, 6.353626e-08, 6.363734e-08, 6.34307e-08, 6.366268e-08, 
    6.279212e-08, 6.32483e-08, 6.253374e-08, 6.274887e-08, 6.289842e-08, 
    6.283283e-08, 6.317353e-08, 6.325383e-08, 6.358018e-08, 6.341148e-08, 
    6.441608e-08, 6.397156e-08, 6.52053e-08, 6.486045e-08, 6.253607e-08, 
    6.264514e-08, 6.302479e-08, 6.284415e-08, 6.336082e-08, 6.348802e-08, 
    6.359143e-08, 6.372361e-08, 6.373789e-08, 6.381621e-08, 6.368786e-08, 
    6.381114e-08, 6.334481e-08, 6.355319e-08, 6.298141e-08, 6.312055e-08, 
    6.305654e-08, 6.298632e-08, 6.320305e-08, 6.343395e-08, 6.34389e-08, 
    6.351294e-08, 6.372157e-08, 6.336292e-08, 6.447343e-08, 6.378752e-08, 
    6.276409e-08, 6.297419e-08, 6.300422e-08, 6.292283e-08, 6.347526e-08, 
    6.327508e-08, 6.38143e-08, 6.366856e-08, 6.390736e-08, 6.37887e-08, 
    6.377123e-08, 6.361883e-08, 6.352395e-08, 6.328425e-08, 6.308925e-08, 
    6.293464e-08, 6.297059e-08, 6.314043e-08, 6.344808e-08, 6.373917e-08, 
    6.367541e-08, 6.388921e-08, 6.332336e-08, 6.356061e-08, 6.34689e-08, 
    6.370803e-08, 6.318411e-08, 6.36302e-08, 6.307009e-08, 6.31192e-08, 
    6.327111e-08, 6.357669e-08, 6.364433e-08, 6.371651e-08, 6.367197e-08, 
    6.34559e-08, 6.34205e-08, 6.326741e-08, 6.322514e-08, 6.310851e-08, 
    6.301195e-08, 6.310017e-08, 6.319282e-08, 6.345599e-08, 6.369318e-08, 
    6.39518e-08, 6.401511e-08, 6.431729e-08, 6.407128e-08, 6.447725e-08, 
    6.413207e-08, 6.472964e-08, 6.365608e-08, 6.412193e-08, 6.327802e-08, 
    6.336893e-08, 6.353335e-08, 6.391052e-08, 6.370691e-08, 6.394504e-08, 
    6.341912e-08, 6.314629e-08, 6.307572e-08, 6.294403e-08, 6.307872e-08, 
    6.306777e-08, 6.319667e-08, 6.315525e-08, 6.346473e-08, 6.329849e-08, 
    6.377079e-08, 6.394317e-08, 6.443005e-08, 6.472857e-08, 6.503251e-08, 
    6.51667e-08, 6.520754e-08, 6.522462e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.681104e-13, 9.707342e-13, 9.702246e-13, 9.723389e-13, 9.711665e-13, 
    9.725504e-13, 9.686429e-13, 9.70838e-13, 9.694371e-13, 9.683471e-13, 
    9.764359e-13, 9.724333e-13, 9.805901e-13, 9.780419e-13, 9.84439e-13, 
    9.801932e-13, 9.852943e-13, 9.843174e-13, 9.872582e-13, 9.864161e-13, 
    9.901719e-13, 9.876468e-13, 9.921177e-13, 9.895696e-13, 9.899681e-13, 
    9.875633e-13, 9.7324e-13, 9.759378e-13, 9.730799e-13, 9.734648e-13, 
    9.732923e-13, 9.711905e-13, 9.701301e-13, 9.679102e-13, 9.683135e-13, 
    9.699442e-13, 9.736379e-13, 9.723851e-13, 9.755428e-13, 9.754715e-13, 
    9.789815e-13, 9.773996e-13, 9.832922e-13, 9.816191e-13, 9.864514e-13, 
    9.85237e-13, 9.863941e-13, 9.860434e-13, 9.863988e-13, 9.846174e-13, 
    9.853807e-13, 9.83813e-13, 9.776958e-13, 9.794949e-13, 9.741246e-13, 
    9.708887e-13, 9.687391e-13, 9.67212e-13, 9.674279e-13, 9.678393e-13, 
    9.699537e-13, 9.719406e-13, 9.734535e-13, 9.744651e-13, 9.754612e-13, 
    9.784723e-13, 9.800662e-13, 9.836301e-13, 9.82988e-13, 9.840761e-13, 
    9.851161e-13, 9.868602e-13, 9.865733e-13, 9.873413e-13, 9.840479e-13, 
    9.862369e-13, 9.82622e-13, 9.836112e-13, 9.757294e-13, 9.727233e-13, 
    9.714423e-13, 9.703225e-13, 9.675938e-13, 9.694783e-13, 9.687355e-13, 
    9.705029e-13, 9.716248e-13, 9.7107e-13, 9.744927e-13, 9.731625e-13, 
    9.801606e-13, 9.771488e-13, 9.849949e-13, 9.831198e-13, 9.854441e-13, 
    9.842585e-13, 9.862894e-13, 9.844618e-13, 9.876273e-13, 9.883157e-13, 
    9.878452e-13, 9.896528e-13, 9.843603e-13, 9.863939e-13, 9.710544e-13, 
    9.711448e-13, 9.715666e-13, 9.697122e-13, 9.695989e-13, 9.67899e-13, 
    9.694118e-13, 9.700555e-13, 9.7169e-13, 9.726558e-13, 9.735737e-13, 
    9.755907e-13, 9.77841e-13, 9.809848e-13, 9.832414e-13, 9.847526e-13, 
    9.838262e-13, 9.846441e-13, 9.837297e-13, 9.833011e-13, 9.880576e-13, 
    9.853878e-13, 9.893929e-13, 9.891715e-13, 9.873595e-13, 9.891965e-13, 
    9.712084e-13, 9.706877e-13, 9.688782e-13, 9.702944e-13, 9.677139e-13, 
    9.691583e-13, 9.699883e-13, 9.731897e-13, 9.738932e-13, 9.745446e-13, 
    9.75831e-13, 9.774806e-13, 9.803716e-13, 9.828846e-13, 9.851767e-13, 
    9.850088e-13, 9.850679e-13, 9.855795e-13, 9.843119e-13, 9.857875e-13, 
    9.860348e-13, 9.853878e-13, 9.891419e-13, 9.8807e-13, 9.891669e-13, 
    9.884691e-13, 9.708571e-13, 9.717332e-13, 9.712597e-13, 9.721498e-13, 
    9.715226e-13, 9.743097e-13, 9.751447e-13, 9.790488e-13, 9.774479e-13, 
    9.799959e-13, 9.777072e-13, 9.781127e-13, 9.800779e-13, 9.77831e-13, 
    9.827456e-13, 9.794138e-13, 9.855993e-13, 9.822751e-13, 9.858074e-13, 
    9.851668e-13, 9.862276e-13, 9.871769e-13, 9.883713e-13, 9.905725e-13, 
    9.900631e-13, 9.919032e-13, 9.73039e-13, 9.741741e-13, 9.740747e-13, 
    9.752625e-13, 9.761404e-13, 9.780428e-13, 9.810904e-13, 9.79945e-13, 
    9.820479e-13, 9.824696e-13, 9.792749e-13, 9.812365e-13, 9.74934e-13, 
    9.759528e-13, 9.753466e-13, 9.731283e-13, 9.802082e-13, 9.765771e-13, 
    9.832786e-13, 9.813147e-13, 9.870416e-13, 9.841947e-13, 9.897825e-13, 
    9.921658e-13, 9.944088e-13, 9.970244e-13, 9.74794e-13, 9.740228e-13, 
    9.754039e-13, 9.773123e-13, 9.79083e-13, 9.814344e-13, 9.816752e-13, 
    9.821152e-13, 9.832554e-13, 9.842133e-13, 9.822539e-13, 9.844534e-13, 
    9.761881e-13, 9.805235e-13, 9.737309e-13, 9.757776e-13, 9.772001e-13, 
    9.765767e-13, 9.798141e-13, 9.805764e-13, 9.836712e-13, 9.820722e-13, 
    9.915773e-13, 9.873767e-13, 9.990156e-13, 9.957689e-13, 9.737533e-13, 
    9.747916e-13, 9.78401e-13, 9.766843e-13, 9.815917e-13, 9.827977e-13, 
    9.837783e-13, 9.850302e-13, 9.851656e-13, 9.859071e-13, 9.846919e-13, 
    9.858593e-13, 9.814395e-13, 9.834157e-13, 9.779893e-13, 9.793108e-13, 
    9.787031e-13, 9.78036e-13, 9.800944e-13, 9.822847e-13, 9.823322e-13, 
    9.830339e-13, 9.850087e-13, 9.816115e-13, 9.921174e-13, 9.856334e-13, 
    9.759232e-13, 9.779198e-13, 9.782058e-13, 9.774325e-13, 9.826768e-13, 
    9.807779e-13, 9.858892e-13, 9.84509e-13, 9.867701e-13, 9.856468e-13, 
    9.854814e-13, 9.840378e-13, 9.831385e-13, 9.808648e-13, 9.790134e-13, 
    9.775448e-13, 9.778864e-13, 9.794995e-13, 9.824187e-13, 9.851775e-13, 
    9.845734e-13, 9.865984e-13, 9.812361e-13, 9.834858e-13, 9.826162e-13, 
    9.848829e-13, 9.799144e-13, 9.841435e-13, 9.788318e-13, 9.792982e-13, 
    9.807402e-13, 9.836377e-13, 9.842794e-13, 9.84963e-13, 9.845413e-13, 
    9.824929e-13, 9.821575e-13, 9.807053e-13, 9.803037e-13, 9.791968e-13, 
    9.782794e-13, 9.791173e-13, 9.799968e-13, 9.824941e-13, 9.847419e-13, 
    9.871904e-13, 9.877895e-13, 9.906442e-13, 9.883195e-13, 9.921533e-13, 
    9.888926e-13, 9.94535e-13, 9.843895e-13, 9.887982e-13, 9.80806e-13, 
    9.816685e-13, 9.83227e-13, 9.867991e-13, 9.848722e-13, 9.87126e-13, 
    9.821445e-13, 9.795547e-13, 9.788852e-13, 9.77634e-13, 9.789138e-13, 
    9.788098e-13, 9.800338e-13, 9.796405e-13, 9.82577e-13, 9.810002e-13, 
    9.85477e-13, 9.871084e-13, 9.917101e-13, 9.94526e-13, 9.9739e-13, 
    9.986528e-13, 9.99037e-13, 9.991976e-13 ;

 LITR1C =
  3.066829e-05, 3.066817e-05, 3.066819e-05, 3.06681e-05, 3.066815e-05, 
    3.066809e-05, 3.066827e-05, 3.066817e-05, 3.066823e-05, 3.066828e-05, 
    3.066791e-05, 3.06681e-05, 3.066772e-05, 3.066784e-05, 3.066755e-05, 
    3.066774e-05, 3.066751e-05, 3.066756e-05, 3.066742e-05, 3.066746e-05, 
    3.066729e-05, 3.06674e-05, 3.06672e-05, 3.066732e-05, 3.06673e-05, 
    3.066741e-05, 3.066806e-05, 3.066794e-05, 3.066807e-05, 3.066805e-05, 
    3.066806e-05, 3.066815e-05, 3.06682e-05, 3.06683e-05, 3.066828e-05, 
    3.066821e-05, 3.066804e-05, 3.06681e-05, 3.066795e-05, 3.066796e-05, 
    3.06678e-05, 3.066787e-05, 3.06676e-05, 3.066768e-05, 3.066746e-05, 
    3.066751e-05, 3.066746e-05, 3.066748e-05, 3.066746e-05, 3.066754e-05, 
    3.066751e-05, 3.066758e-05, 3.066786e-05, 3.066778e-05, 3.066802e-05, 
    3.066816e-05, 3.066826e-05, 3.066833e-05, 3.066832e-05, 3.06683e-05, 
    3.066821e-05, 3.066812e-05, 3.066805e-05, 3.0668e-05, 3.066796e-05, 
    3.066782e-05, 3.066775e-05, 3.066759e-05, 3.066762e-05, 3.066757e-05, 
    3.066752e-05, 3.066744e-05, 3.066746e-05, 3.066742e-05, 3.066757e-05, 
    3.066747e-05, 3.066763e-05, 3.066759e-05, 3.066795e-05, 3.066808e-05, 
    3.066814e-05, 3.066819e-05, 3.066831e-05, 3.066823e-05, 3.066826e-05, 
    3.066818e-05, 3.066813e-05, 3.066816e-05, 3.0668e-05, 3.066806e-05, 
    3.066775e-05, 3.066788e-05, 3.066752e-05, 3.066761e-05, 3.066751e-05, 
    3.066756e-05, 3.066747e-05, 3.066755e-05, 3.066741e-05, 3.066738e-05, 
    3.06674e-05, 3.066731e-05, 3.066755e-05, 3.066746e-05, 3.066816e-05, 
    3.066815e-05, 3.066814e-05, 3.066822e-05, 3.066822e-05, 3.06683e-05, 
    3.066823e-05, 3.06682e-05, 3.066813e-05, 3.066808e-05, 3.066804e-05, 
    3.066795e-05, 3.066785e-05, 3.066771e-05, 3.06676e-05, 3.066754e-05, 
    3.066758e-05, 3.066754e-05, 3.066758e-05, 3.06676e-05, 3.066739e-05, 
    3.066751e-05, 3.066733e-05, 3.066734e-05, 3.066742e-05, 3.066734e-05, 
    3.066815e-05, 3.066817e-05, 3.066826e-05, 3.066819e-05, 3.066831e-05, 
    3.066824e-05, 3.06682e-05, 3.066806e-05, 3.066803e-05, 3.0668e-05, 
    3.066794e-05, 3.066787e-05, 3.066774e-05, 3.066762e-05, 3.066752e-05, 
    3.066752e-05, 3.066752e-05, 3.06675e-05, 3.066756e-05, 3.066749e-05, 
    3.066748e-05, 3.066751e-05, 3.066734e-05, 3.066739e-05, 3.066734e-05, 
    3.066737e-05, 3.066816e-05, 3.066812e-05, 3.066815e-05, 3.066811e-05, 
    3.066814e-05, 3.066801e-05, 3.066797e-05, 3.066779e-05, 3.066787e-05, 
    3.066775e-05, 3.066786e-05, 3.066784e-05, 3.066775e-05, 3.066785e-05, 
    3.066763e-05, 3.066778e-05, 3.06675e-05, 3.066765e-05, 3.066749e-05, 
    3.066752e-05, 3.066747e-05, 3.066743e-05, 3.066737e-05, 3.066727e-05, 
    3.06673e-05, 3.066721e-05, 3.066807e-05, 3.066802e-05, 3.066802e-05, 
    3.066797e-05, 3.066793e-05, 3.066784e-05, 3.06677e-05, 3.066775e-05, 
    3.066766e-05, 3.066764e-05, 3.066779e-05, 3.06677e-05, 3.066798e-05, 
    3.066794e-05, 3.066796e-05, 3.066806e-05, 3.066774e-05, 3.066791e-05, 
    3.06676e-05, 3.066769e-05, 3.066743e-05, 3.066756e-05, 3.066731e-05, 
    3.06672e-05, 3.06671e-05, 3.066698e-05, 3.066799e-05, 3.066802e-05, 
    3.066796e-05, 3.066787e-05, 3.066779e-05, 3.066769e-05, 3.066768e-05, 
    3.066766e-05, 3.06676e-05, 3.066756e-05, 3.066765e-05, 3.066755e-05, 
    3.066792e-05, 3.066773e-05, 3.066804e-05, 3.066794e-05, 3.066788e-05, 
    3.066791e-05, 3.066776e-05, 3.066772e-05, 3.066759e-05, 3.066766e-05, 
    3.066723e-05, 3.066742e-05, 3.066689e-05, 3.066704e-05, 3.066803e-05, 
    3.066799e-05, 3.066782e-05, 3.06679e-05, 3.066768e-05, 3.066763e-05, 
    3.066758e-05, 3.066752e-05, 3.066752e-05, 3.066748e-05, 3.066754e-05, 
    3.066749e-05, 3.066769e-05, 3.06676e-05, 3.066784e-05, 3.066778e-05, 
    3.066781e-05, 3.066784e-05, 3.066775e-05, 3.066765e-05, 3.066764e-05, 
    3.066762e-05, 3.066752e-05, 3.066768e-05, 3.06672e-05, 3.06675e-05, 
    3.066794e-05, 3.066784e-05, 3.066783e-05, 3.066787e-05, 3.066763e-05, 
    3.066772e-05, 3.066748e-05, 3.066755e-05, 3.066744e-05, 3.06675e-05, 
    3.06675e-05, 3.066757e-05, 3.066761e-05, 3.066771e-05, 3.06678e-05, 
    3.066786e-05, 3.066785e-05, 3.066778e-05, 3.066764e-05, 3.066752e-05, 
    3.066755e-05, 3.066745e-05, 3.06677e-05, 3.066759e-05, 3.066763e-05, 
    3.066753e-05, 3.066776e-05, 3.066756e-05, 3.06678e-05, 3.066778e-05, 
    3.066772e-05, 3.066759e-05, 3.066756e-05, 3.066753e-05, 3.066755e-05, 
    3.066764e-05, 3.066766e-05, 3.066772e-05, 3.066774e-05, 3.066779e-05, 
    3.066783e-05, 3.066779e-05, 3.066775e-05, 3.066764e-05, 3.066754e-05, 
    3.066743e-05, 3.06674e-05, 3.066727e-05, 3.066738e-05, 3.06672e-05, 
    3.066735e-05, 3.06671e-05, 3.066755e-05, 3.066735e-05, 3.066771e-05, 
    3.066768e-05, 3.06676e-05, 3.066744e-05, 3.066753e-05, 3.066743e-05, 
    3.066766e-05, 3.066777e-05, 3.06678e-05, 3.066786e-05, 3.06678e-05, 
    3.06678e-05, 3.066775e-05, 3.066777e-05, 3.066763e-05, 3.066771e-05, 
    3.06675e-05, 3.066743e-05, 3.066722e-05, 3.06671e-05, 3.066696e-05, 
    3.066691e-05, 3.066689e-05, 3.066688e-05 ;

 LITR1C_TO_SOIL1C =
  6.448038e-13, 6.46551e-13, 6.462117e-13, 6.476196e-13, 6.468389e-13, 
    6.477605e-13, 6.451584e-13, 6.466202e-13, 6.456873e-13, 6.449615e-13, 
    6.503479e-13, 6.476824e-13, 6.531142e-13, 6.514173e-13, 6.556772e-13, 
    6.5285e-13, 6.562468e-13, 6.555963e-13, 6.575546e-13, 6.569939e-13, 
    6.594949e-13, 6.578134e-13, 6.607906e-13, 6.590938e-13, 6.593591e-13, 
    6.577578e-13, 6.482197e-13, 6.500162e-13, 6.481131e-13, 6.483694e-13, 
    6.482545e-13, 6.468549e-13, 6.461487e-13, 6.446705e-13, 6.449391e-13, 
    6.46025e-13, 6.484847e-13, 6.476504e-13, 6.497531e-13, 6.497057e-13, 
    6.520431e-13, 6.509896e-13, 6.549136e-13, 6.537995e-13, 6.570173e-13, 
    6.562086e-13, 6.569792e-13, 6.567457e-13, 6.569823e-13, 6.557961e-13, 
    6.563044e-13, 6.552604e-13, 6.511869e-13, 6.523849e-13, 6.488088e-13, 
    6.46654e-13, 6.452224e-13, 6.442055e-13, 6.443493e-13, 6.446233e-13, 
    6.460313e-13, 6.473544e-13, 6.483619e-13, 6.490355e-13, 6.496989e-13, 
    6.51704e-13, 6.527654e-13, 6.551385e-13, 6.54711e-13, 6.554356e-13, 
    6.561281e-13, 6.572896e-13, 6.570986e-13, 6.576099e-13, 6.554168e-13, 
    6.568746e-13, 6.544673e-13, 6.55126e-13, 6.498775e-13, 6.478756e-13, 
    6.470225e-13, 6.462768e-13, 6.444598e-13, 6.457147e-13, 6.452201e-13, 
    6.463969e-13, 6.471441e-13, 6.467747e-13, 6.490539e-13, 6.48168e-13, 
    6.528282e-13, 6.508226e-13, 6.560474e-13, 6.547988e-13, 6.563466e-13, 
    6.55557e-13, 6.569095e-13, 6.556924e-13, 6.578004e-13, 6.582588e-13, 
    6.579455e-13, 6.591492e-13, 6.556248e-13, 6.569791e-13, 6.467642e-13, 
    6.468245e-13, 6.471053e-13, 6.458705e-13, 6.45795e-13, 6.44663e-13, 
    6.456705e-13, 6.460991e-13, 6.471875e-13, 6.478306e-13, 6.484419e-13, 
    6.497851e-13, 6.512836e-13, 6.533771e-13, 6.548797e-13, 6.558861e-13, 
    6.552692e-13, 6.558138e-13, 6.552049e-13, 6.549195e-13, 6.580869e-13, 
    6.56309e-13, 6.589761e-13, 6.588287e-13, 6.57622e-13, 6.588454e-13, 
    6.468668e-13, 6.465201e-13, 6.453151e-13, 6.462582e-13, 6.445398e-13, 
    6.455016e-13, 6.460543e-13, 6.481862e-13, 6.486546e-13, 6.490884e-13, 
    6.499451e-13, 6.510436e-13, 6.529687e-13, 6.546421e-13, 6.561685e-13, 
    6.560568e-13, 6.560961e-13, 6.564367e-13, 6.555926e-13, 6.565752e-13, 
    6.567399e-13, 6.56309e-13, 6.58809e-13, 6.580952e-13, 6.588256e-13, 
    6.58361e-13, 6.466328e-13, 6.472163e-13, 6.46901e-13, 6.474937e-13, 
    6.47076e-13, 6.48932e-13, 6.494881e-13, 6.520879e-13, 6.510218e-13, 
    6.527185e-13, 6.511944e-13, 6.514645e-13, 6.527731e-13, 6.512769e-13, 
    6.545496e-13, 6.523309e-13, 6.564499e-13, 6.542363e-13, 6.565885e-13, 
    6.561619e-13, 6.568683e-13, 6.575005e-13, 6.582958e-13, 6.597616e-13, 
    6.594224e-13, 6.606478e-13, 6.480859e-13, 6.488417e-13, 6.487755e-13, 
    6.495665e-13, 6.501512e-13, 6.514179e-13, 6.534474e-13, 6.526846e-13, 
    6.54085e-13, 6.543658e-13, 6.522385e-13, 6.535447e-13, 6.493477e-13, 
    6.500262e-13, 6.496225e-13, 6.481453e-13, 6.528599e-13, 6.504419e-13, 
    6.549045e-13, 6.535968e-13, 6.574103e-13, 6.555146e-13, 6.592356e-13, 
    6.608226e-13, 6.623162e-13, 6.640581e-13, 6.492545e-13, 6.48741e-13, 
    6.496607e-13, 6.509315e-13, 6.521106e-13, 6.536765e-13, 6.538368e-13, 
    6.541299e-13, 6.548891e-13, 6.55527e-13, 6.542222e-13, 6.556868e-13, 
    6.501829e-13, 6.530699e-13, 6.485465e-13, 6.499095e-13, 6.508568e-13, 
    6.504416e-13, 6.525975e-13, 6.531051e-13, 6.55166e-13, 6.541012e-13, 
    6.604307e-13, 6.576336e-13, 6.65384e-13, 6.632219e-13, 6.485615e-13, 
    6.492529e-13, 6.516565e-13, 6.505133e-13, 6.537812e-13, 6.545844e-13, 
    6.552373e-13, 6.560709e-13, 6.561612e-13, 6.566549e-13, 6.558457e-13, 
    6.566231e-13, 6.536799e-13, 6.549959e-13, 6.513823e-13, 6.522624e-13, 
    6.518576e-13, 6.514134e-13, 6.527841e-13, 6.542426e-13, 6.542743e-13, 
    6.547416e-13, 6.560566e-13, 6.537944e-13, 6.607904e-13, 6.564727e-13, 
    6.500065e-13, 6.51336e-13, 6.515265e-13, 6.510116e-13, 6.545038e-13, 
    6.532393e-13, 6.566429e-13, 6.557239e-13, 6.572296e-13, 6.564815e-13, 
    6.563714e-13, 6.554101e-13, 6.548112e-13, 6.532972e-13, 6.520643e-13, 
    6.510863e-13, 6.513138e-13, 6.52388e-13, 6.543319e-13, 6.561691e-13, 
    6.557668e-13, 6.571152e-13, 6.535444e-13, 6.550424e-13, 6.544635e-13, 
    6.559728e-13, 6.526642e-13, 6.554805e-13, 6.519434e-13, 6.522539e-13, 
    6.532142e-13, 6.551436e-13, 6.55571e-13, 6.560262e-13, 6.557454e-13, 
    6.543813e-13, 6.54158e-13, 6.53191e-13, 6.529236e-13, 6.521864e-13, 
    6.515755e-13, 6.521335e-13, 6.527191e-13, 6.543821e-13, 6.558789e-13, 
    6.575094e-13, 6.579084e-13, 6.598094e-13, 6.582613e-13, 6.608143e-13, 
    6.58643e-13, 6.624003e-13, 6.556443e-13, 6.585801e-13, 6.53258e-13, 
    6.538324e-13, 6.548701e-13, 6.572489e-13, 6.559657e-13, 6.574665e-13, 
    6.541493e-13, 6.524247e-13, 6.519789e-13, 6.511457e-13, 6.519979e-13, 
    6.519287e-13, 6.527438e-13, 6.524819e-13, 6.544373e-13, 6.533873e-13, 
    6.563685e-13, 6.574548e-13, 6.605192e-13, 6.623943e-13, 6.643015e-13, 
    6.651424e-13, 6.653982e-13, 6.655052e-13 ;

 LITR1C_vr =
  0.001751191, 0.001751184, 0.001751186, 0.00175118, 0.001751183, 0.00175118, 
    0.00175119, 0.001751184, 0.001751188, 0.001751191, 0.00175117, 
    0.00175118, 0.001751159, 0.001751165, 0.001751149, 0.00175116, 
    0.001751147, 0.001751149, 0.001751142, 0.001751144, 0.001751134, 
    0.001751141, 0.001751129, 0.001751136, 0.001751135, 0.001751141, 
    0.001751178, 0.001751171, 0.001751178, 0.001751177, 0.001751178, 
    0.001751183, 0.001751186, 0.001751192, 0.001751191, 0.001751186, 
    0.001751177, 0.00175118, 0.001751172, 0.001751172, 0.001751163, 
    0.001751167, 0.001751152, 0.001751156, 0.001751144, 0.001751147, 
    0.001751144, 0.001751145, 0.001751144, 0.001751148, 0.001751146, 
    0.00175115, 0.001751166, 0.001751162, 0.001751175, 0.001751184, 
    0.001751189, 0.001751193, 0.001751193, 0.001751192, 0.001751186, 
    0.001751181, 0.001751177, 0.001751175, 0.001751172, 0.001751164, 
    0.00175116, 0.001751151, 0.001751153, 0.00175115, 0.001751147, 
    0.001751143, 0.001751143, 0.001751141, 0.00175115, 0.001751144, 
    0.001751153, 0.001751151, 0.001751171, 0.001751179, 0.001751182, 
    0.001751185, 0.001751192, 0.001751188, 0.001751189, 0.001751185, 
    0.001751182, 0.001751183, 0.001751175, 0.001751178, 0.00175116, 
    0.001751168, 0.001751147, 0.001751152, 0.001751146, 0.001751149, 
    0.001751144, 0.001751149, 0.001751141, 0.001751139, 0.00175114, 
    0.001751135, 0.001751149, 0.001751144, 0.001751183, 0.001751183, 
    0.001751182, 0.001751187, 0.001751187, 0.001751192, 0.001751188, 
    0.001751186, 0.001751182, 0.001751179, 0.001751177, 0.001751172, 
    0.001751166, 0.001751158, 0.001751152, 0.001751148, 0.00175115, 
    0.001751148, 0.001751151, 0.001751152, 0.00175114, 0.001751146, 
    0.001751136, 0.001751137, 0.001751141, 0.001751137, 0.001751183, 
    0.001751184, 0.001751189, 0.001751185, 0.001751192, 0.001751188, 
    0.001751186, 0.001751178, 0.001751176, 0.001751174, 0.001751171, 
    0.001751167, 0.001751159, 0.001751153, 0.001751147, 0.001751147, 
    0.001751147, 0.001751146, 0.001751149, 0.001751145, 0.001751145, 
    0.001751146, 0.001751137, 0.001751139, 0.001751137, 0.001751138, 
    0.001751184, 0.001751182, 0.001751183, 0.001751181, 0.001751182, 
    0.001751175, 0.001751173, 0.001751163, 0.001751167, 0.00175116, 
    0.001751166, 0.001751165, 0.00175116, 0.001751166, 0.001751153, 
    0.001751162, 0.001751146, 0.001751154, 0.001751145, 0.001751147, 
    0.001751144, 0.001751142, 0.001751139, 0.001751133, 0.001751134, 
    0.00175113, 0.001751178, 0.001751175, 0.001751176, 0.001751173, 
    0.00175117, 0.001751165, 0.001751158, 0.00175116, 0.001751155, 
    0.001751154, 0.001751162, 0.001751157, 0.001751173, 0.001751171, 
    0.001751172, 0.001751178, 0.00175116, 0.001751169, 0.001751152, 
    0.001751157, 0.001751142, 0.00175115, 0.001751135, 0.001751129, 
    0.001751123, 0.001751116, 0.001751174, 0.001751176, 0.001751172, 
    0.001751167, 0.001751163, 0.001751157, 0.001751156, 0.001751155, 
    0.001751152, 0.001751149, 0.001751155, 0.001751149, 0.00175117, 
    0.001751159, 0.001751177, 0.001751171, 0.001751168, 0.001751169, 
    0.001751161, 0.001751159, 0.001751151, 0.001751155, 0.00175113, 
    0.001751141, 0.001751111, 0.00175112, 0.001751177, 0.001751174, 
    0.001751164, 0.001751169, 0.001751156, 0.001751153, 0.001751151, 
    0.001751147, 0.001751147, 0.001751145, 0.001751148, 0.001751145, 
    0.001751157, 0.001751152, 0.001751165, 0.001751162, 0.001751164, 
    0.001751165, 0.00175116, 0.001751154, 0.001751154, 0.001751152, 
    0.001751147, 0.001751156, 0.001751129, 0.001751146, 0.001751171, 
    0.001751166, 0.001751165, 0.001751167, 0.001751153, 0.001751158, 
    0.001751145, 0.001751149, 0.001751143, 0.001751146, 0.001751146, 
    0.00175115, 0.001751152, 0.001751158, 0.001751163, 0.001751167, 
    0.001751166, 0.001751162, 0.001751154, 0.001751147, 0.001751148, 
    0.001751143, 0.001751157, 0.001751151, 0.001751154, 0.001751148, 
    0.001751161, 0.00175115, 0.001751163, 0.001751162, 0.001751158, 
    0.001751151, 0.001751149, 0.001751147, 0.001751149, 0.001751154, 
    0.001751155, 0.001751159, 0.00175116, 0.001751162, 0.001751165, 
    0.001751163, 0.00175116, 0.001751154, 0.001751148, 0.001751142, 
    0.00175114, 0.001751133, 0.001751139, 0.001751129, 0.001751137, 
    0.001751123, 0.001751149, 0.001751138, 0.001751158, 0.001751156, 
    0.001751152, 0.001751143, 0.001751148, 0.001751142, 0.001751155, 
    0.001751162, 0.001751163, 0.001751166, 0.001751163, 0.001751163, 
    0.00175116, 0.001751161, 0.001751154, 0.001751158, 0.001751146, 
    0.001751142, 0.00175113, 0.001751123, 0.001751115, 0.001751112, 
    0.001751111, 0.001751111,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.732976e-07, 9.732938e-07, 9.732946e-07, 9.732915e-07, 9.732933e-07, 
    9.732912e-07, 9.732969e-07, 9.732937e-07, 9.732958e-07, 9.732972e-07, 
    9.732856e-07, 9.732914e-07, 9.732797e-07, 9.732834e-07, 9.732742e-07, 
    9.732803e-07, 9.732729e-07, 9.732743e-07, 9.732701e-07, 9.732713e-07, 
    9.732659e-07, 9.732695e-07, 9.732631e-07, 9.732668e-07, 9.732662e-07, 
    9.732696e-07, 9.732903e-07, 9.732863e-07, 9.732905e-07, 9.7329e-07, 
    9.732902e-07, 9.732931e-07, 9.732947e-07, 9.732979e-07, 9.732973e-07, 
    9.73295e-07, 9.732897e-07, 9.732914e-07, 9.732869e-07, 9.73287e-07, 
    9.73282e-07, 9.732843e-07, 9.732757e-07, 9.732782e-07, 9.732713e-07, 
    9.73273e-07, 9.732713e-07, 9.732719e-07, 9.732713e-07, 9.732739e-07, 
    9.732728e-07, 9.732751e-07, 9.732838e-07, 9.732812e-07, 9.732889e-07, 
    9.732936e-07, 9.732967e-07, 9.732989e-07, 9.732986e-07, 9.73298e-07, 
    9.73295e-07, 9.732921e-07, 9.7329e-07, 9.732885e-07, 9.73287e-07, 
    9.732827e-07, 9.732804e-07, 9.732753e-07, 9.732762e-07, 9.732747e-07, 
    9.732731e-07, 9.732706e-07, 9.732711e-07, 9.732699e-07, 9.732747e-07, 
    9.732715e-07, 9.732768e-07, 9.732753e-07, 9.732867e-07, 9.73291e-07, 
    9.732928e-07, 9.732944e-07, 9.732984e-07, 9.732956e-07, 9.732968e-07, 
    9.732942e-07, 9.732926e-07, 9.732934e-07, 9.732885e-07, 9.732904e-07, 
    9.732803e-07, 9.732846e-07, 9.732734e-07, 9.732761e-07, 9.732727e-07, 
    9.732744e-07, 9.732715e-07, 9.732742e-07, 9.732696e-07, 9.732686e-07, 
    9.732693e-07, 9.732667e-07, 9.732743e-07, 9.732713e-07, 9.732934e-07, 
    9.732933e-07, 9.732927e-07, 9.732953e-07, 9.732955e-07, 9.732979e-07, 
    9.732958e-07, 9.732948e-07, 9.732925e-07, 9.732911e-07, 9.732897e-07, 
    9.732869e-07, 9.732836e-07, 9.732792e-07, 9.732759e-07, 9.732737e-07, 
    9.732751e-07, 9.732738e-07, 9.732752e-07, 9.732757e-07, 9.732689e-07, 
    9.732728e-07, 9.73267e-07, 9.732673e-07, 9.732699e-07, 9.732673e-07, 
    9.732931e-07, 9.732939e-07, 9.732966e-07, 9.732945e-07, 9.732981e-07, 
    9.732961e-07, 9.73295e-07, 9.732903e-07, 9.732893e-07, 9.732884e-07, 
    9.732865e-07, 9.732842e-07, 9.7328e-07, 9.732764e-07, 9.732731e-07, 
    9.732734e-07, 9.732732e-07, 9.732726e-07, 9.732744e-07, 9.732722e-07, 
    9.732719e-07, 9.732728e-07, 9.732673e-07, 9.732689e-07, 9.732673e-07, 
    9.732684e-07, 9.732937e-07, 9.732925e-07, 9.732931e-07, 9.732918e-07, 
    9.732927e-07, 9.732887e-07, 9.732875e-07, 9.732819e-07, 9.732842e-07, 
    9.732805e-07, 9.732838e-07, 9.732832e-07, 9.732804e-07, 9.732837e-07, 
    9.732765e-07, 9.732814e-07, 9.732724e-07, 9.732772e-07, 9.732722e-07, 
    9.732731e-07, 9.732715e-07, 9.732702e-07, 9.732685e-07, 9.732653e-07, 
    9.732661e-07, 9.732635e-07, 9.732905e-07, 9.732889e-07, 9.73289e-07, 
    9.732873e-07, 9.732861e-07, 9.732834e-07, 9.732789e-07, 9.732806e-07, 
    9.732776e-07, 9.73277e-07, 9.732815e-07, 9.732787e-07, 9.732878e-07, 
    9.732863e-07, 9.732872e-07, 9.732904e-07, 9.732802e-07, 9.732854e-07, 
    9.732759e-07, 9.732786e-07, 9.732704e-07, 9.732745e-07, 9.732664e-07, 
    9.73263e-07, 9.732598e-07, 9.732561e-07, 9.73288e-07, 9.732892e-07, 
    9.732871e-07, 9.732844e-07, 9.732819e-07, 9.732785e-07, 9.732781e-07, 
    9.732775e-07, 9.732759e-07, 9.732745e-07, 9.732773e-07, 9.732742e-07, 
    9.73286e-07, 9.732797e-07, 9.732895e-07, 9.732865e-07, 9.732846e-07, 
    9.732854e-07, 9.732807e-07, 9.732797e-07, 9.732753e-07, 9.732776e-07, 
    9.732639e-07, 9.732699e-07, 9.732532e-07, 9.732579e-07, 9.732895e-07, 
    9.73288e-07, 9.732828e-07, 9.732853e-07, 9.732782e-07, 9.732765e-07, 
    9.732751e-07, 9.732732e-07, 9.732731e-07, 9.73272e-07, 9.732738e-07, 
    9.732721e-07, 9.732785e-07, 9.732756e-07, 9.732835e-07, 9.732815e-07, 
    9.732823e-07, 9.732834e-07, 9.732804e-07, 9.732772e-07, 9.732772e-07, 
    9.732762e-07, 9.732734e-07, 9.732782e-07, 9.732631e-07, 9.732724e-07, 
    9.732864e-07, 9.732835e-07, 9.732831e-07, 9.732843e-07, 9.732767e-07, 
    9.732794e-07, 9.732721e-07, 9.73274e-07, 9.732707e-07, 9.732724e-07, 
    9.732727e-07, 9.732747e-07, 9.73276e-07, 9.732793e-07, 9.73282e-07, 
    9.73284e-07, 9.732836e-07, 9.732812e-07, 9.732771e-07, 9.732731e-07, 
    9.732739e-07, 9.732711e-07, 9.732787e-07, 9.732755e-07, 9.732768e-07, 
    9.732735e-07, 9.732806e-07, 9.732746e-07, 9.732822e-07, 9.732815e-07, 
    9.732795e-07, 9.732753e-07, 9.732744e-07, 9.732734e-07, 9.73274e-07, 
    9.73277e-07, 9.732775e-07, 9.732795e-07, 9.732801e-07, 9.732817e-07, 
    9.73283e-07, 9.732818e-07, 9.732805e-07, 9.73277e-07, 9.732737e-07, 
    9.732702e-07, 9.732694e-07, 9.732652e-07, 9.732686e-07, 9.73263e-07, 
    9.732678e-07, 9.732596e-07, 9.732743e-07, 9.732679e-07, 9.732794e-07, 
    9.732781e-07, 9.732759e-07, 9.732707e-07, 9.732735e-07, 9.732703e-07, 
    9.732775e-07, 9.732812e-07, 9.732821e-07, 9.732839e-07, 9.732821e-07, 
    9.732822e-07, 9.732805e-07, 9.732811e-07, 9.732769e-07, 9.73279e-07, 
    9.732727e-07, 9.732703e-07, 9.732637e-07, 9.732596e-07, 9.732555e-07, 
    9.732537e-07, 9.732531e-07, 9.732529e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  -1.56858e-25, 7.352717e-25, 3.921449e-25, 8.82326e-26, -5.048866e-25, 
    -3.676358e-25, 3.333231e-25, -3.921449e-25, 1.068595e-24, -1.323489e-25, 
    3.823413e-25, 5.490028e-25, 1.171533e-24, -9.803622e-26, 2.352869e-25, 
    -3.62734e-25, 1.02938e-25, -2.352869e-25, -5.882173e-25, 9.656568e-25, 
    7.205662e-25, -1.56858e-25, -1.862688e-25, -4.705739e-25, -2.009742e-25, 
    -5.146902e-25, 4.264576e-25, -9.803622e-27, 1.107809e-24, 1.147024e-24, 
    -7.842898e-26, 2.450906e-25, 3.578322e-25, -6.323336e-25, 4.803775e-25, 
    -4.901811e-25, -3.921449e-26, 1.960724e-25, 5.19592e-25, -5.048866e-25, 
    3.921449e-26, -2.695996e-25, -2.646978e-25, 3.823413e-25, -2.843051e-25, 
    -9.656568e-25, -3.578322e-25, -1.960724e-25, -4.264576e-25, 2.892069e-25, 
    -4.215557e-25, -4.019485e-25, -2.892069e-25, 4.803775e-25, 2.254833e-25, 
    -1.274471e-25, 4.509666e-25, 4.117521e-25, 9.803622e-27, 8.82326e-26, 
    6.960572e-25, -9.803622e-26, 7.646825e-25, 2.450906e-25, 1.372507e-25, 
    -3.529304e-25, 5.98021e-25, 8.235043e-25, -1.117613e-24, 6.862535e-26, 
    -5.391992e-25, -2.156797e-25, 2.548942e-25, 4.803775e-25, 2.59796e-25, 
    -9.803622e-27, 1.372507e-25, 2.450906e-25, 4.41163e-25, -2.843051e-25, 
    3.872431e-25, -4.901811e-26, -9.803622e-26, 2.941087e-26, 3.921449e-25, 
    3.823413e-25, 3.38225e-25, 0, -6.274318e-25, -1.274471e-25, 
    -4.901811e-26, 2.499924e-25, -3.284213e-25, -2.794032e-25, 4.705739e-25, 
    8.82326e-26, -5.293956e-25, 7.597807e-25, 1.470543e-25, -7.842898e-26, 
    -4.901811e-26, 2.548942e-25, -2.058761e-25, 1.421525e-25, 6.372354e-25, 
    4.901811e-26, -6.911554e-25, -5.293956e-25, 1.274471e-25, 2.646978e-25, 
    -2.941087e-26, -3.62734e-25, 9.509513e-25, -1.078398e-25, -8.82326e-26, 
    8.82326e-26, 2.009742e-25, -3.823413e-25, 2.254833e-25, 2.941087e-25, 
    1.078398e-25, 8.235043e-25, 7.058608e-25, 2.058761e-25, -3.921449e-26, 
    1.56858e-25, 3.62734e-25, 3.039123e-25, 2.254833e-25, 4.460648e-25, 
    8.82326e-26, 7.352717e-26, -2.352869e-25, 1.176435e-25, 4.803775e-25, 
    2.548942e-25, 1.81367e-25, -1.019577e-24, -3.921449e-26, 2.941087e-26, 
    4.901811e-26, -2.941087e-26, 3.921449e-25, -1.421525e-25, -6.127264e-25, 
    -4.019485e-25, 3.235195e-25, -5.882173e-26, -2.156797e-25, 5.391992e-25, 
    -7.940934e-25, -2.646978e-25, -3.431268e-26, -3.823413e-25, 7.891916e-25, 
    -3.921449e-26, -8.82326e-25, -4.509666e-25, -6.862535e-26, -1.715634e-25, 
    1.519561e-25, 8.82326e-26, -1.666616e-25, -4.901811e-26, 5.686101e-25, 
    8.333079e-26, 5.244938e-25, 3.529304e-25, -2.352869e-25, 4.901811e-27, 
    8.529151e-25, -3.529304e-25, -8.82326e-26, 1.078398e-25, -6.862535e-26, 
    2.450906e-25, 2.058761e-25, -3.872431e-25, 4.901811e-26, 9.509513e-25, 
    1.911706e-25, 3.039123e-25, -2.695996e-25, -1.56858e-25, 5.391992e-26, 
    -7.744861e-25, -1.073497e-24, -3.823413e-25, 4.019485e-25, -1.666616e-25, 
    1.200944e-24, 3.921449e-25, -3.823413e-25, 1.764652e-25, 6.372354e-25, 
    -2.009742e-25, 4.41163e-25, 6.862535e-26, -8.431115e-25, 4.117521e-25, 
    -4.264576e-25, -1.81367e-25, 9.215405e-25, 7.058608e-25, -4.41163e-26, 
    6.421373e-25, 7.646825e-25, -4.019485e-25, 5.588064e-25, 4.166539e-25, 
    9.117368e-25, 2.745014e-25, 3.529304e-25, 9.803622e-26, 2.450905e-26, 
    1.372507e-25, 9.313441e-25, 1.421525e-25, 4.852793e-25, 9.803622e-26, 
    -2.450906e-25, -5.490028e-25, 9.803622e-27, 4.705739e-25, -9.411477e-25, 
    -7.548789e-25, 5.44101e-25, 2.303851e-25, -3.235195e-25, 3.480286e-25, 
    -3.431268e-25, -1.960724e-26, -2.450905e-26, 3.431268e-25, -3.725376e-25, 
    -5.784137e-25, -3.725376e-25, -5.686101e-25, -5.146902e-25, 
    -8.921296e-25, -5.882173e-26, -6.176282e-25, -4.41163e-25, 5.244938e-25, 
    5.391992e-25, 2.156797e-25, 3.480286e-25, 3.921449e-26, -5.882173e-26, 
    2.794032e-25, 1.078398e-25, 4.803775e-25, -3.921449e-25, -4.901811e-26, 
    -4.999847e-25, -3.431268e-25, -3.921449e-26, 8.333079e-26, 1.666616e-25, 
    2.941087e-25, 4.019485e-25, 7.842898e-26, 3.039123e-25, 4.901811e-26, 
    -5.882173e-26, -6.568427e-25, -7.25468e-25, 4.901811e-27, 4.509666e-25, 
    -2.646978e-25, -1.764652e-25, 1.009773e-24, -3.921449e-26, 5.244938e-25, 
    1.274471e-25, 1.960724e-25, 1.225453e-25, -7.646825e-25, -5.44101e-25, 
    4.362612e-25, -3.578322e-25, 3.676358e-25, -1.960724e-25, -1.617598e-25, 
    -1.078398e-25, -6.176282e-25, 2.499924e-25, 2.59796e-25, -1.078398e-25, 
    5.293956e-25, 1.960724e-26, 4.068503e-25, 1.176435e-25, -2.843051e-25, 
    4.460648e-25, -1.56858e-25, -3.480286e-25, 7.842898e-26, 1.862688e-25, 
    -6.862535e-26, -2.401887e-25, 6.372354e-25, -4.901811e-26, -3.235195e-25, 
    9.803622e-27, 6.764499e-25, -2.352869e-25, -1.470543e-25, 6.176282e-25, 
    4.215557e-25, 1.862688e-25, -1.960724e-26, -2.941087e-25, 1.470543e-25, 
    9.117368e-25, 5.882173e-26, 1.960724e-25, 9.460495e-25, -3.872431e-25, 
    1.264667e-24, 2.941087e-26, -1.862688e-25, 4.41163e-25, 2.107779e-25, 
    -1.764652e-25, -3.823413e-25, 5.882173e-26, 4.215557e-25, 2.941087e-26, 
    1.666616e-25, 3.921449e-25, 8.333079e-26, 9.803622e-26, -1.666616e-25, 
    -1.225453e-24, 1.862688e-25, 5.882173e-26, 2.401887e-25,
  9.436816e-32, 9.436779e-32, 9.436786e-32, 9.436755e-32, 9.436772e-32, 
    9.436752e-32, 9.436809e-32, 9.436777e-32, 9.436798e-32, 9.436813e-32, 
    9.436696e-32, 9.436754e-32, 9.436636e-32, 9.436673e-32, 9.436581e-32, 
    9.436642e-32, 9.436568e-32, 9.436582e-32, 9.43654e-32, 9.436552e-32, 
    9.436498e-32, 9.436534e-32, 9.43647e-32, 9.436507e-32, 9.436501e-32, 
    9.436535e-32, 9.436742e-32, 9.436703e-32, 9.436745e-32, 9.436739e-32, 
    9.436742e-32, 9.436772e-32, 9.436788e-32, 9.436819e-32, 9.436813e-32, 
    9.43679e-32, 9.436736e-32, 9.436755e-32, 9.436709e-32, 9.43671e-32, 
    9.436659e-32, 9.436682e-32, 9.436597e-32, 9.436621e-32, 9.436552e-32, 
    9.436569e-32, 9.436552e-32, 9.436558e-32, 9.436552e-32, 9.436578e-32, 
    9.436567e-32, 9.436589e-32, 9.436678e-32, 9.436652e-32, 9.436729e-32, 
    9.436776e-32, 9.436808e-32, 9.436829e-32, 9.436826e-32, 9.43682e-32, 
    9.43679e-32, 9.436761e-32, 9.436739e-32, 9.436725e-32, 9.436711e-32, 
    9.436667e-32, 9.436644e-32, 9.436592e-32, 9.436602e-32, 9.436586e-32, 
    9.436571e-32, 9.436545e-32, 9.43655e-32, 9.436539e-32, 9.436587e-32, 
    9.436555e-32, 9.436607e-32, 9.436592e-32, 9.436706e-32, 9.43675e-32, 
    9.436768e-32, 9.436785e-32, 9.436824e-32, 9.436797e-32, 9.436808e-32, 
    9.436782e-32, 9.436766e-32, 9.436773e-32, 9.436724e-32, 9.436743e-32, 
    9.436642e-32, 9.436686e-32, 9.436572e-32, 9.436599e-32, 9.436566e-32, 
    9.436583e-32, 9.436554e-32, 9.43658e-32, 9.436535e-32, 9.436525e-32, 
    9.436531e-32, 9.436505e-32, 9.436582e-32, 9.436552e-32, 9.436774e-32, 
    9.436773e-32, 9.436766e-32, 9.436793e-32, 9.436795e-32, 9.436819e-32, 
    9.436798e-32, 9.436788e-32, 9.436765e-32, 9.436751e-32, 9.436738e-32, 
    9.436708e-32, 9.436676e-32, 9.436631e-32, 9.436598e-32, 9.436576e-32, 
    9.436589e-32, 9.436578e-32, 9.436591e-32, 9.436597e-32, 9.436528e-32, 
    9.436567e-32, 9.436509e-32, 9.436512e-32, 9.436538e-32, 9.436512e-32, 
    9.436772e-32, 9.436779e-32, 9.436805e-32, 9.436785e-32, 9.436822e-32, 
    9.436801e-32, 9.436789e-32, 9.436743e-32, 9.436733e-32, 9.436723e-32, 
    9.436705e-32, 9.436681e-32, 9.436639e-32, 9.436603e-32, 9.43657e-32, 
    9.436572e-32, 9.436572e-32, 9.436564e-32, 9.436582e-32, 9.436561e-32, 
    9.436558e-32, 9.436567e-32, 9.436512e-32, 9.436528e-32, 9.436512e-32, 
    9.436522e-32, 9.436777e-32, 9.436764e-32, 9.436771e-32, 9.436758e-32, 
    9.436767e-32, 9.436727e-32, 9.436715e-32, 9.436658e-32, 9.436682e-32, 
    9.436645e-32, 9.436678e-32, 9.436672e-32, 9.436644e-32, 9.436676e-32, 
    9.436605e-32, 9.436653e-32, 9.436564e-32, 9.436612e-32, 9.436561e-32, 
    9.43657e-32, 9.436555e-32, 9.436541e-32, 9.436524e-32, 9.436492e-32, 
    9.4365e-32, 9.436473e-32, 9.436745e-32, 9.436729e-32, 9.436731e-32, 
    9.436713e-32, 9.436701e-32, 9.436673e-32, 9.436629e-32, 9.436645e-32, 
    9.436615e-32, 9.436609e-32, 9.436655e-32, 9.436627e-32, 9.436718e-32, 
    9.436703e-32, 9.436712e-32, 9.436744e-32, 9.436642e-32, 9.436694e-32, 
    9.436597e-32, 9.436626e-32, 9.436543e-32, 9.436584e-32, 9.436504e-32, 
    9.436469e-32, 9.436437e-32, 9.436399e-32, 9.43672e-32, 9.436731e-32, 
    9.436711e-32, 9.436684e-32, 9.436658e-32, 9.436624e-32, 9.436621e-32, 
    9.436614e-32, 9.436598e-32, 9.436584e-32, 9.436612e-32, 9.436581e-32, 
    9.4367e-32, 9.436637e-32, 9.436735e-32, 9.436706e-32, 9.436685e-32, 
    9.436694e-32, 9.436648e-32, 9.436636e-32, 9.436592e-32, 9.436615e-32, 
    9.436478e-32, 9.436538e-32, 9.43637e-32, 9.436417e-32, 9.436735e-32, 
    9.43672e-32, 9.436668e-32, 9.436693e-32, 9.436622e-32, 9.436604e-32, 
    9.43659e-32, 9.436572e-32, 9.43657e-32, 9.436559e-32, 9.436577e-32, 
    9.43656e-32, 9.436624e-32, 9.436595e-32, 9.436674e-32, 9.436655e-32, 
    9.436664e-32, 9.436673e-32, 9.436644e-32, 9.436612e-32, 9.436611e-32, 
    9.436601e-32, 9.436572e-32, 9.436621e-32, 9.43647e-32, 9.436564e-32, 
    9.436703e-32, 9.436675e-32, 9.436671e-32, 9.436682e-32, 9.436606e-32, 
    9.436634e-32, 9.436559e-32, 9.436579e-32, 9.436547e-32, 9.436563e-32, 
    9.436565e-32, 9.436587e-32, 9.436599e-32, 9.436632e-32, 9.436659e-32, 
    9.43668e-32, 9.436675e-32, 9.436652e-32, 9.43661e-32, 9.43657e-32, 
    9.436579e-32, 9.43655e-32, 9.436627e-32, 9.436594e-32, 9.436607e-32, 
    9.436574e-32, 9.436646e-32, 9.436585e-32, 9.436662e-32, 9.436655e-32, 
    9.436634e-32, 9.436592e-32, 9.436583e-32, 9.436573e-32, 9.436579e-32, 
    9.436609e-32, 9.436614e-32, 9.436635e-32, 9.436641e-32, 9.436656e-32, 
    9.436669e-32, 9.436658e-32, 9.436645e-32, 9.436609e-32, 9.436577e-32, 
    9.436541e-32, 9.436532e-32, 9.436491e-32, 9.436525e-32, 9.436469e-32, 
    9.436517e-32, 9.436435e-32, 9.436581e-32, 9.436518e-32, 9.436633e-32, 
    9.436621e-32, 9.436598e-32, 9.436547e-32, 9.436574e-32, 9.436542e-32, 
    9.436614e-32, 9.436651e-32, 9.436661e-32, 9.436679e-32, 9.436661e-32, 
    9.436662e-32, 9.436644e-32, 9.43665e-32, 9.436608e-32, 9.43663e-32, 
    9.436565e-32, 9.436542e-32, 9.436475e-32, 9.436435e-32, 9.436394e-32, 
    9.436376e-32, 9.43637e-32, 9.436367e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.547479e-14, 4.559802e-14, 4.557408e-14, 4.567338e-14, 4.561832e-14, 
    4.568331e-14, 4.54998e-14, 4.560289e-14, 4.55371e-14, 4.548591e-14, 
    4.586579e-14, 4.567781e-14, 4.606089e-14, 4.594121e-14, 4.624164e-14, 
    4.604225e-14, 4.628181e-14, 4.623593e-14, 4.637404e-14, 4.63345e-14, 
    4.651088e-14, 4.639229e-14, 4.660226e-14, 4.648259e-14, 4.650131e-14, 
    4.638837e-14, 4.57157e-14, 4.584239e-14, 4.570818e-14, 4.572626e-14, 
    4.571815e-14, 4.561944e-14, 4.556964e-14, 4.546539e-14, 4.548433e-14, 
    4.556091e-14, 4.573439e-14, 4.567555e-14, 4.582385e-14, 4.58205e-14, 
    4.598534e-14, 4.591105e-14, 4.618779e-14, 4.610921e-14, 4.633615e-14, 
    4.627912e-14, 4.633346e-14, 4.631699e-14, 4.633368e-14, 4.625003e-14, 
    4.628587e-14, 4.621224e-14, 4.592496e-14, 4.600945e-14, 4.575724e-14, 
    4.560527e-14, 4.550432e-14, 4.54326e-14, 4.544274e-14, 4.546206e-14, 
    4.556136e-14, 4.565468e-14, 4.572573e-14, 4.577323e-14, 4.582002e-14, 
    4.596143e-14, 4.603628e-14, 4.620365e-14, 4.61735e-14, 4.62246e-14, 
    4.627344e-14, 4.635535e-14, 4.634188e-14, 4.637794e-14, 4.622328e-14, 
    4.632608e-14, 4.615631e-14, 4.620277e-14, 4.583261e-14, 4.569143e-14, 
    4.563127e-14, 4.557868e-14, 4.545053e-14, 4.553904e-14, 4.550415e-14, 
    4.558715e-14, 4.563984e-14, 4.561379e-14, 4.577453e-14, 4.571206e-14, 
    4.604072e-14, 4.589927e-14, 4.626774e-14, 4.617969e-14, 4.628885e-14, 
    4.623317e-14, 4.632854e-14, 4.624271e-14, 4.639137e-14, 4.64237e-14, 
    4.640161e-14, 4.64865e-14, 4.623795e-14, 4.633345e-14, 4.561305e-14, 
    4.56173e-14, 4.563711e-14, 4.555002e-14, 4.55447e-14, 4.546487e-14, 
    4.553591e-14, 4.556614e-14, 4.56429e-14, 4.568826e-14, 4.573137e-14, 
    4.58261e-14, 4.593177e-14, 4.607943e-14, 4.61854e-14, 4.625637e-14, 
    4.621286e-14, 4.625128e-14, 4.620833e-14, 4.618821e-14, 4.641158e-14, 
    4.62862e-14, 4.64743e-14, 4.64639e-14, 4.63788e-14, 4.646507e-14, 
    4.562029e-14, 4.559583e-14, 4.551085e-14, 4.557736e-14, 4.545617e-14, 
    4.552401e-14, 4.556299e-14, 4.571333e-14, 4.574637e-14, 4.577696e-14, 
    4.583738e-14, 4.591485e-14, 4.605063e-14, 4.616864e-14, 4.627629e-14, 
    4.626841e-14, 4.627118e-14, 4.62952e-14, 4.623567e-14, 4.630497e-14, 
    4.631659e-14, 4.62862e-14, 4.646251e-14, 4.641217e-14, 4.646368e-14, 
    4.643091e-14, 4.560379e-14, 4.564493e-14, 4.56227e-14, 4.56645e-14, 
    4.563504e-14, 4.576594e-14, 4.580515e-14, 4.59885e-14, 4.591332e-14, 
    4.603298e-14, 4.592549e-14, 4.594454e-14, 4.603683e-14, 4.593131e-14, 
    4.616212e-14, 4.600564e-14, 4.629613e-14, 4.614002e-14, 4.630591e-14, 
    4.627582e-14, 4.632564e-14, 4.637023e-14, 4.642632e-14, 4.652969e-14, 
    4.650577e-14, 4.659219e-14, 4.570626e-14, 4.575957e-14, 4.57549e-14, 
    4.581068e-14, 4.585191e-14, 4.594126e-14, 4.608438e-14, 4.603059e-14, 
    4.612935e-14, 4.614915e-14, 4.599912e-14, 4.609124e-14, 4.579525e-14, 
    4.58431e-14, 4.581463e-14, 4.571045e-14, 4.604295e-14, 4.587242e-14, 
    4.618714e-14, 4.609492e-14, 4.636387e-14, 4.623017e-14, 4.649259e-14, 
    4.660452e-14, 4.670986e-14, 4.68327e-14, 4.578868e-14, 4.575246e-14, 
    4.581732e-14, 4.590695e-14, 4.599011e-14, 4.610054e-14, 4.611185e-14, 
    4.613251e-14, 4.618605e-14, 4.623104e-14, 4.613902e-14, 4.624232e-14, 
    4.585415e-14, 4.605776e-14, 4.573875e-14, 4.583487e-14, 4.590167e-14, 
    4.58724e-14, 4.602444e-14, 4.606025e-14, 4.620558e-14, 4.613049e-14, 
    4.657688e-14, 4.637961e-14, 4.692621e-14, 4.677373e-14, 4.57398e-14, 
    4.578857e-14, 4.595808e-14, 4.587746e-14, 4.610792e-14, 4.616457e-14, 
    4.621061e-14, 4.626941e-14, 4.627577e-14, 4.631059e-14, 4.625352e-14, 
    4.630835e-14, 4.610077e-14, 4.619359e-14, 4.593874e-14, 4.600081e-14, 
    4.597227e-14, 4.594094e-14, 4.60376e-14, 4.614047e-14, 4.61427e-14, 
    4.617566e-14, 4.62684e-14, 4.610886e-14, 4.660225e-14, 4.629774e-14, 
    4.584171e-14, 4.593548e-14, 4.594891e-14, 4.591259e-14, 4.615888e-14, 
    4.606971e-14, 4.630975e-14, 4.624493e-14, 4.635112e-14, 4.629836e-14, 
    4.62906e-14, 4.62228e-14, 4.618056e-14, 4.607379e-14, 4.598684e-14, 
    4.591787e-14, 4.593391e-14, 4.600966e-14, 4.614676e-14, 4.627633e-14, 
    4.624795e-14, 4.634306e-14, 4.609123e-14, 4.619687e-14, 4.615604e-14, 
    4.626249e-14, 4.602915e-14, 4.622776e-14, 4.597831e-14, 4.600021e-14, 
    4.606793e-14, 4.620401e-14, 4.623415e-14, 4.626625e-14, 4.624645e-14, 
    4.615025e-14, 4.61345e-14, 4.60663e-14, 4.604744e-14, 4.599545e-14, 
    4.595237e-14, 4.599172e-14, 4.603302e-14, 4.615031e-14, 4.625587e-14, 
    4.637086e-14, 4.639899e-14, 4.653306e-14, 4.642389e-14, 4.660393e-14, 
    4.64508e-14, 4.671578e-14, 4.623932e-14, 4.644637e-14, 4.607103e-14, 
    4.611154e-14, 4.618472e-14, 4.635248e-14, 4.626199e-14, 4.636783e-14, 
    4.613388e-14, 4.601226e-14, 4.598082e-14, 4.592205e-14, 4.598216e-14, 
    4.597727e-14, 4.603476e-14, 4.601629e-14, 4.61542e-14, 4.608015e-14, 
    4.629039e-14, 4.636701e-14, 4.658312e-14, 4.671536e-14, 4.684986e-14, 
    4.690917e-14, 4.692722e-14, 4.693476e-14 ;

 LITR1N_vr =
  5.55763e-05, 5.557609e-05, 5.557613e-05, 5.557595e-05, 5.557605e-05, 
    5.557594e-05, 5.557626e-05, 5.557607e-05, 5.557619e-05, 5.557628e-05, 
    5.557562e-05, 5.557594e-05, 5.557527e-05, 5.557549e-05, 5.557496e-05, 
    5.557531e-05, 5.557489e-05, 5.557497e-05, 5.557473e-05, 5.55748e-05, 
    5.557449e-05, 5.55747e-05, 5.557433e-05, 5.557454e-05, 5.557451e-05, 
    5.55747e-05, 5.557588e-05, 5.557566e-05, 5.557589e-05, 5.557586e-05, 
    5.557587e-05, 5.557605e-05, 5.557613e-05, 5.557632e-05, 5.557628e-05, 
    5.557615e-05, 5.557585e-05, 5.557595e-05, 5.557569e-05, 5.55757e-05, 
    5.557541e-05, 5.557554e-05, 5.557505e-05, 5.557519e-05, 5.557479e-05, 
    5.55749e-05, 5.55748e-05, 5.557483e-05, 5.55748e-05, 5.557495e-05, 
    5.557488e-05, 5.557501e-05, 5.557551e-05, 5.557536e-05, 5.557581e-05, 
    5.557607e-05, 5.557625e-05, 5.557637e-05, 5.557635e-05, 5.557632e-05, 
    5.557615e-05, 5.557599e-05, 5.557586e-05, 5.557578e-05, 5.55757e-05, 
    5.557545e-05, 5.557532e-05, 5.557503e-05, 5.557508e-05, 5.557499e-05, 
    5.55749e-05, 5.557476e-05, 5.557478e-05, 5.557472e-05, 5.557499e-05, 
    5.557481e-05, 5.557511e-05, 5.557503e-05, 5.557567e-05, 5.557592e-05, 
    5.557603e-05, 5.557612e-05, 5.557634e-05, 5.557619e-05, 5.557625e-05, 
    5.55761e-05, 5.557601e-05, 5.557606e-05, 5.557578e-05, 5.557589e-05, 
    5.557531e-05, 5.557556e-05, 5.557491e-05, 5.557507e-05, 5.557488e-05, 
    5.557498e-05, 5.557481e-05, 5.557496e-05, 5.55747e-05, 5.557464e-05, 
    5.557468e-05, 5.557453e-05, 5.557496e-05, 5.55748e-05, 5.557606e-05, 
    5.557605e-05, 5.557602e-05, 5.557617e-05, 5.557618e-05, 5.557632e-05, 
    5.557619e-05, 5.557614e-05, 5.557601e-05, 5.557593e-05, 5.557585e-05, 
    5.557569e-05, 5.55755e-05, 5.557524e-05, 5.557506e-05, 5.557494e-05, 
    5.557501e-05, 5.557494e-05, 5.557502e-05, 5.557505e-05, 5.557466e-05, 
    5.557488e-05, 5.557455e-05, 5.557457e-05, 5.557472e-05, 5.557457e-05, 
    5.557605e-05, 5.557609e-05, 5.557624e-05, 5.557612e-05, 5.557633e-05, 
    5.557621e-05, 5.557615e-05, 5.557588e-05, 5.557583e-05, 5.557577e-05, 
    5.557567e-05, 5.557553e-05, 5.557529e-05, 5.557509e-05, 5.55749e-05, 
    5.557491e-05, 5.557491e-05, 5.557487e-05, 5.557497e-05, 5.557485e-05, 
    5.557483e-05, 5.557488e-05, 5.557457e-05, 5.557466e-05, 5.557457e-05, 
    5.557463e-05, 5.557607e-05, 5.5576e-05, 5.557604e-05, 5.557597e-05, 
    5.557602e-05, 5.557579e-05, 5.557572e-05, 5.55754e-05, 5.557553e-05, 
    5.557532e-05, 5.557551e-05, 5.557548e-05, 5.557532e-05, 5.55755e-05, 
    5.55751e-05, 5.557537e-05, 5.557486e-05, 5.557514e-05, 5.557485e-05, 
    5.55749e-05, 5.557481e-05, 5.557474e-05, 5.557464e-05, 5.557446e-05, 
    5.55745e-05, 5.557435e-05, 5.55759e-05, 5.55758e-05, 5.557581e-05, 
    5.557571e-05, 5.557564e-05, 5.557549e-05, 5.557523e-05, 5.557533e-05, 
    5.557516e-05, 5.557512e-05, 5.557538e-05, 5.557522e-05, 5.557574e-05, 
    5.557566e-05, 5.557571e-05, 5.557589e-05, 5.557531e-05, 5.557561e-05, 
    5.557506e-05, 5.557522e-05, 5.557475e-05, 5.557498e-05, 5.557452e-05, 
    5.557432e-05, 5.557414e-05, 5.557393e-05, 5.557575e-05, 5.557582e-05, 
    5.55757e-05, 5.557554e-05, 5.55754e-05, 5.55752e-05, 5.557519e-05, 
    5.557515e-05, 5.557506e-05, 5.557498e-05, 5.557514e-05, 5.557496e-05, 
    5.557564e-05, 5.557528e-05, 5.557584e-05, 5.557567e-05, 5.557555e-05, 
    5.557561e-05, 5.557534e-05, 5.557528e-05, 5.557502e-05, 5.557515e-05, 
    5.557438e-05, 5.557472e-05, 5.557376e-05, 5.557403e-05, 5.557584e-05, 
    5.557575e-05, 5.557546e-05, 5.55756e-05, 5.557519e-05, 5.55751e-05, 
    5.557502e-05, 5.557491e-05, 5.55749e-05, 5.557484e-05, 5.557494e-05, 
    5.557484e-05, 5.55752e-05, 5.557504e-05, 5.557549e-05, 5.557538e-05, 
    5.557543e-05, 5.557549e-05, 5.557532e-05, 5.557514e-05, 5.557513e-05, 
    5.557507e-05, 5.557491e-05, 5.557519e-05, 5.557433e-05, 5.557486e-05, 
    5.557566e-05, 5.55755e-05, 5.557547e-05, 5.557554e-05, 5.55751e-05, 
    5.557526e-05, 5.557484e-05, 5.557495e-05, 5.557477e-05, 5.557486e-05, 
    5.557487e-05, 5.557499e-05, 5.557507e-05, 5.557525e-05, 5.55754e-05, 
    5.557553e-05, 5.55755e-05, 5.557536e-05, 5.557512e-05, 5.55749e-05, 
    5.557495e-05, 5.557478e-05, 5.557522e-05, 5.557504e-05, 5.557511e-05, 
    5.557492e-05, 5.557533e-05, 5.557498e-05, 5.557542e-05, 5.557538e-05, 
    5.557526e-05, 5.557503e-05, 5.557497e-05, 5.557492e-05, 5.557495e-05, 
    5.557512e-05, 5.557515e-05, 5.557527e-05, 5.55753e-05, 5.557539e-05, 
    5.557547e-05, 5.55754e-05, 5.557532e-05, 5.557512e-05, 5.557494e-05, 
    5.557474e-05, 5.557468e-05, 5.557445e-05, 5.557464e-05, 5.557433e-05, 
    5.557459e-05, 5.557413e-05, 5.557496e-05, 5.55746e-05, 5.557526e-05, 
    5.557519e-05, 5.557506e-05, 5.557476e-05, 5.557492e-05, 5.557474e-05, 
    5.557515e-05, 5.557536e-05, 5.557542e-05, 5.557552e-05, 5.557541e-05, 
    5.557542e-05, 5.557532e-05, 5.557535e-05, 5.557511e-05, 5.557524e-05, 
    5.557487e-05, 5.557474e-05, 5.557436e-05, 5.557413e-05, 5.55739e-05, 
    5.557379e-05, 5.557376e-05, 5.557375e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.880935e-13, 7.90229e-13, 7.898142e-13, 7.915351e-13, 7.905809e-13, 
    7.917072e-13, 7.885269e-13, 7.903135e-13, 7.891734e-13, 7.882862e-13, 
    7.948696e-13, 7.916119e-13, 7.982507e-13, 7.961767e-13, 8.013833e-13, 
    7.979277e-13, 8.020794e-13, 8.012843e-13, 8.036779e-13, 8.029925e-13, 
    8.060493e-13, 8.039941e-13, 8.076329e-13, 8.055591e-13, 8.058834e-13, 
    8.039262e-13, 7.922685e-13, 7.944642e-13, 7.921382e-13, 7.924515e-13, 
    7.92311e-13, 7.906004e-13, 7.897374e-13, 7.879306e-13, 7.882589e-13, 
    7.89586e-13, 7.925924e-13, 7.915728e-13, 7.941427e-13, 7.940847e-13, 
    7.969416e-13, 7.95654e-13, 8.0045e-13, 7.990882e-13, 8.030212e-13, 
    8.020328e-13, 8.029746e-13, 8.026891e-13, 8.029783e-13, 8.015285e-13, 
    8.021498e-13, 8.008738e-13, 7.958951e-13, 7.973594e-13, 7.929885e-13, 
    7.903548e-13, 7.886052e-13, 7.873623e-13, 7.87538e-13, 7.878729e-13, 
    7.895938e-13, 7.91211e-13, 7.924423e-13, 7.932656e-13, 7.940764e-13, 
    7.965271e-13, 7.978243e-13, 8.007249e-13, 8.002023e-13, 8.010879e-13, 
    8.019344e-13, 8.03354e-13, 8.031205e-13, 8.037455e-13, 8.01065e-13, 
    8.028467e-13, 7.999045e-13, 8.007095e-13, 7.942946e-13, 7.91848e-13, 
    7.908054e-13, 7.898939e-13, 7.876731e-13, 7.892069e-13, 7.886024e-13, 
    7.900407e-13, 7.909538e-13, 7.905024e-13, 7.932881e-13, 7.922054e-13, 
    7.979012e-13, 7.954499e-13, 8.018357e-13, 8.003096e-13, 8.022014e-13, 
    8.012364e-13, 8.028893e-13, 8.014018e-13, 8.039782e-13, 8.045385e-13, 
    8.041556e-13, 8.056268e-13, 8.013192e-13, 8.029744e-13, 7.904896e-13, 
    7.905633e-13, 7.909065e-13, 7.893972e-13, 7.89305e-13, 7.879215e-13, 
    7.891528e-13, 7.896767e-13, 7.91007e-13, 7.91793e-13, 7.925401e-13, 
    7.941817e-13, 7.960132e-13, 7.98572e-13, 8.004086e-13, 8.016385e-13, 
    8.008846e-13, 8.015502e-13, 8.00806e-13, 8.004572e-13, 8.043284e-13, 
    8.021555e-13, 8.054153e-13, 8.052351e-13, 8.037603e-13, 8.052554e-13, 
    7.90615e-13, 7.901912e-13, 7.887184e-13, 7.898711e-13, 7.877708e-13, 
    7.889464e-13, 7.896219e-13, 7.922276e-13, 7.928001e-13, 7.933302e-13, 
    7.943773e-13, 7.957199e-13, 7.980729e-13, 8.001182e-13, 8.019838e-13, 
    8.018471e-13, 8.018952e-13, 8.023115e-13, 8.012799e-13, 8.024808e-13, 
    8.026821e-13, 8.021555e-13, 8.05211e-13, 8.043386e-13, 8.052313e-13, 
    8.046634e-13, 7.90329e-13, 7.910421e-13, 7.906568e-13, 7.913812e-13, 
    7.908707e-13, 7.931392e-13, 7.938187e-13, 7.969963e-13, 7.956934e-13, 
    7.977671e-13, 7.959042e-13, 7.962344e-13, 7.978339e-13, 7.960051e-13, 
    8.000051e-13, 7.972933e-13, 8.023277e-13, 7.996222e-13, 8.024971e-13, 
    8.019757e-13, 8.02839e-13, 8.036117e-13, 8.045838e-13, 8.063754e-13, 
    8.059607e-13, 8.074584e-13, 7.921049e-13, 7.930288e-13, 7.929478e-13, 
    7.939146e-13, 7.946292e-13, 7.961775e-13, 7.986579e-13, 7.977257e-13, 
    7.994372e-13, 7.997804e-13, 7.971803e-13, 7.987768e-13, 7.936472e-13, 
    7.944765e-13, 7.93983e-13, 7.921776e-13, 7.979399e-13, 7.949846e-13, 
    8.004388e-13, 7.988405e-13, 8.035015e-13, 8.011845e-13, 8.057323e-13, 
    8.07672e-13, 8.094977e-13, 8.116265e-13, 7.935333e-13, 7.929057e-13, 
    7.940297e-13, 7.955829e-13, 7.970241e-13, 7.98938e-13, 7.991339e-13, 
    7.99492e-13, 8.0042e-13, 8.011996e-13, 7.996049e-13, 8.01395e-13, 
    7.946679e-13, 7.981965e-13, 7.92668e-13, 7.943338e-13, 7.954915e-13, 
    7.949842e-13, 7.976192e-13, 7.982396e-13, 8.007584e-13, 7.99457e-13, 
    8.071931e-13, 8.037743e-13, 8.132471e-13, 8.106046e-13, 7.926862e-13, 
    7.935314e-13, 7.96469e-13, 7.950719e-13, 7.990658e-13, 8.000475e-13, 
    8.008455e-13, 8.018644e-13, 8.019748e-13, 8.025782e-13, 8.015892e-13, 
    8.025393e-13, 7.98942e-13, 8.005505e-13, 7.961339e-13, 7.972095e-13, 
    7.967149e-13, 7.961719e-13, 7.978472e-13, 7.996299e-13, 7.996686e-13, 
    8.002397e-13, 8.01847e-13, 7.99082e-13, 8.076327e-13, 8.023555e-13, 
    7.944524e-13, 7.960774e-13, 7.963102e-13, 7.956808e-13, 7.999491e-13, 
    7.984036e-13, 8.025636e-13, 8.014403e-13, 8.032806e-13, 8.023663e-13, 
    8.022317e-13, 8.010569e-13, 8.003248e-13, 7.984744e-13, 7.969675e-13, 
    7.957722e-13, 7.960502e-13, 7.97363e-13, 7.99739e-13, 8.019844e-13, 
    8.014927e-13, 8.031408e-13, 7.987765e-13, 8.006074e-13, 7.998998e-13, 
    8.017445e-13, 7.977007e-13, 8.011428e-13, 7.968197e-13, 7.971992e-13, 
    7.983729e-13, 8.007311e-13, 8.012534e-13, 8.018098e-13, 8.014666e-13, 
    7.997994e-13, 7.995264e-13, 7.983445e-13, 7.980177e-13, 7.971167e-13, 
    7.963701e-13, 7.97052e-13, 7.977678e-13, 7.998004e-13, 8.016298e-13, 
    8.036226e-13, 8.041103e-13, 8.064337e-13, 8.045417e-13, 8.076619e-13, 
    8.050081e-13, 8.096003e-13, 8.013431e-13, 8.049313e-13, 7.984265e-13, 
    7.991285e-13, 8.003969e-13, 8.033042e-13, 8.017359e-13, 8.035702e-13, 
    7.995158e-13, 7.97408e-13, 7.968631e-13, 7.958447e-13, 7.968864e-13, 
    7.968017e-13, 7.977979e-13, 7.974779e-13, 7.998679e-13, 7.985845e-13, 
    8.022282e-13, 8.035559e-13, 8.073012e-13, 8.09593e-13, 8.11924e-13, 
    8.129518e-13, 8.132645e-13, 8.133952e-13 ;

 LITR2C =
  1.939604e-05, 1.939602e-05, 1.939603e-05, 1.939601e-05, 1.939602e-05, 
    1.939601e-05, 1.939604e-05, 1.939602e-05, 1.939603e-05, 1.939604e-05, 
    1.939598e-05, 1.939601e-05, 1.939595e-05, 1.939597e-05, 1.939592e-05, 
    1.939595e-05, 1.939591e-05, 1.939592e-05, 1.93959e-05, 1.93959e-05, 
    1.939587e-05, 1.939589e-05, 1.939586e-05, 1.939588e-05, 1.939588e-05, 
    1.939589e-05, 1.9396e-05, 1.939598e-05, 1.939601e-05, 1.9396e-05, 
    1.9396e-05, 1.939602e-05, 1.939603e-05, 1.939604e-05, 1.939604e-05, 
    1.939603e-05, 1.9396e-05, 1.939601e-05, 1.939599e-05, 1.939599e-05, 
    1.939596e-05, 1.939597e-05, 1.939593e-05, 1.939594e-05, 1.93959e-05, 
    1.939591e-05, 1.93959e-05, 1.939591e-05, 1.93959e-05, 1.939592e-05, 
    1.939591e-05, 1.939592e-05, 1.939597e-05, 1.939596e-05, 1.9396e-05, 
    1.939602e-05, 1.939604e-05, 1.939605e-05, 1.939605e-05, 1.939604e-05, 
    1.939603e-05, 1.939601e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.939596e-05, 1.939595e-05, 1.939593e-05, 1.939593e-05, 1.939592e-05, 
    1.939591e-05, 1.93959e-05, 1.93959e-05, 1.93959e-05, 1.939592e-05, 
    1.939591e-05, 1.939593e-05, 1.939593e-05, 1.939599e-05, 1.939601e-05, 
    1.939602e-05, 1.939603e-05, 1.939605e-05, 1.939603e-05, 1.939604e-05, 
    1.939602e-05, 1.939602e-05, 1.939602e-05, 1.939599e-05, 1.9396e-05, 
    1.939595e-05, 1.939597e-05, 1.939591e-05, 1.939593e-05, 1.939591e-05, 
    1.939592e-05, 1.939591e-05, 1.939592e-05, 1.939589e-05, 1.939589e-05, 
    1.939589e-05, 1.939588e-05, 1.939592e-05, 1.93959e-05, 1.939602e-05, 
    1.939602e-05, 1.939602e-05, 1.939603e-05, 1.939603e-05, 1.939604e-05, 
    1.939603e-05, 1.939603e-05, 1.939601e-05, 1.939601e-05, 1.9396e-05, 
    1.939599e-05, 1.939597e-05, 1.939595e-05, 1.939593e-05, 1.939592e-05, 
    1.939592e-05, 1.939592e-05, 1.939592e-05, 1.939593e-05, 1.939589e-05, 
    1.939591e-05, 1.939588e-05, 1.939588e-05, 1.93959e-05, 1.939588e-05, 
    1.939602e-05, 1.939602e-05, 1.939604e-05, 1.939603e-05, 1.939605e-05, 
    1.939603e-05, 1.939603e-05, 1.9396e-05, 1.9396e-05, 1.939599e-05, 
    1.939598e-05, 1.939597e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 
    1.939591e-05, 1.939591e-05, 1.939591e-05, 1.939592e-05, 1.939591e-05, 
    1.939591e-05, 1.939591e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939589e-05, 1.939602e-05, 1.939601e-05, 1.939602e-05, 1.939601e-05, 
    1.939602e-05, 1.939599e-05, 1.939599e-05, 1.939596e-05, 1.939597e-05, 
    1.939595e-05, 1.939597e-05, 1.939597e-05, 1.939595e-05, 1.939597e-05, 
    1.939593e-05, 1.939596e-05, 1.939591e-05, 1.939593e-05, 1.939591e-05, 
    1.939591e-05, 1.939591e-05, 1.93959e-05, 1.939589e-05, 1.939587e-05, 
    1.939588e-05, 1.939586e-05, 1.939601e-05, 1.9396e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939594e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939596e-05, 1.939594e-05, 1.939599e-05, 
    1.939598e-05, 1.939599e-05, 1.9396e-05, 1.939595e-05, 1.939598e-05, 
    1.939593e-05, 1.939594e-05, 1.93959e-05, 1.939592e-05, 1.939588e-05, 
    1.939586e-05, 1.939584e-05, 1.939582e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939597e-05, 1.939596e-05, 1.939594e-05, 1.939594e-05, 
    1.939594e-05, 1.939593e-05, 1.939592e-05, 1.939593e-05, 1.939592e-05, 
    1.939598e-05, 1.939595e-05, 1.9396e-05, 1.939598e-05, 1.939597e-05, 
    1.939598e-05, 1.939595e-05, 1.939595e-05, 1.939592e-05, 1.939594e-05, 
    1.939587e-05, 1.93959e-05, 1.939581e-05, 1.939583e-05, 1.9396e-05, 
    1.939599e-05, 1.939596e-05, 1.939598e-05, 1.939594e-05, 1.939593e-05, 
    1.939592e-05, 1.939591e-05, 1.939591e-05, 1.939591e-05, 1.939592e-05, 
    1.939591e-05, 1.939594e-05, 1.939593e-05, 1.939597e-05, 1.939596e-05, 
    1.939596e-05, 1.939597e-05, 1.939595e-05, 1.939593e-05, 1.939593e-05, 
    1.939593e-05, 1.939591e-05, 1.939594e-05, 1.939586e-05, 1.939591e-05, 
    1.939598e-05, 1.939597e-05, 1.939597e-05, 1.939597e-05, 1.939593e-05, 
    1.939595e-05, 1.939591e-05, 1.939592e-05, 1.93959e-05, 1.939591e-05, 
    1.939591e-05, 1.939592e-05, 1.939593e-05, 1.939595e-05, 1.939596e-05, 
    1.939597e-05, 1.939597e-05, 1.939596e-05, 1.939593e-05, 1.939591e-05, 
    1.939592e-05, 1.93959e-05, 1.939594e-05, 1.939593e-05, 1.939593e-05, 
    1.939591e-05, 1.939595e-05, 1.939592e-05, 1.939596e-05, 1.939596e-05, 
    1.939595e-05, 1.939593e-05, 1.939592e-05, 1.939591e-05, 1.939592e-05, 
    1.939593e-05, 1.939594e-05, 1.939595e-05, 1.939595e-05, 1.939596e-05, 
    1.939597e-05, 1.939596e-05, 1.939595e-05, 1.939593e-05, 1.939592e-05, 
    1.93959e-05, 1.939589e-05, 1.939587e-05, 1.939589e-05, 1.939586e-05, 
    1.939589e-05, 1.939584e-05, 1.939592e-05, 1.939589e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.93959e-05, 1.939591e-05, 1.93959e-05, 
    1.939594e-05, 1.939596e-05, 1.939596e-05, 1.939597e-05, 1.939596e-05, 
    1.939596e-05, 1.939595e-05, 1.939595e-05, 1.939593e-05, 1.939595e-05, 
    1.939591e-05, 1.93959e-05, 1.939586e-05, 1.939584e-05, 1.939582e-05, 
    1.939581e-05, 1.939581e-05, 1.939581e-05 ;

 LITR2C_TO_SOIL1C =
  1.200113e-13, 1.203368e-13, 1.202736e-13, 1.205359e-13, 1.203904e-13, 
    1.205621e-13, 1.200773e-13, 1.203497e-13, 1.201759e-13, 1.200406e-13, 
    1.210442e-13, 1.205476e-13, 1.215596e-13, 1.212434e-13, 1.220371e-13, 
    1.215104e-13, 1.221432e-13, 1.22022e-13, 1.223869e-13, 1.222824e-13, 
    1.227484e-13, 1.224351e-13, 1.229898e-13, 1.226737e-13, 1.227231e-13, 
    1.224248e-13, 1.206477e-13, 1.209824e-13, 1.206278e-13, 1.206756e-13, 
    1.206542e-13, 1.203934e-13, 1.202618e-13, 1.199864e-13, 1.200365e-13, 
    1.202388e-13, 1.20697e-13, 1.205416e-13, 1.209334e-13, 1.209245e-13, 
    1.2136e-13, 1.211638e-13, 1.218949e-13, 1.216873e-13, 1.222868e-13, 
    1.221361e-13, 1.222797e-13, 1.222362e-13, 1.222803e-13, 1.220593e-13, 
    1.22154e-13, 1.219595e-13, 1.212005e-13, 1.214237e-13, 1.207574e-13, 
    1.20356e-13, 1.200893e-13, 1.198998e-13, 1.199266e-13, 1.199776e-13, 
    1.202399e-13, 1.204865e-13, 1.206742e-13, 1.207997e-13, 1.209233e-13, 
    1.212969e-13, 1.214946e-13, 1.219368e-13, 1.218571e-13, 1.219921e-13, 
    1.221211e-13, 1.223375e-13, 1.223019e-13, 1.223972e-13, 1.219886e-13, 
    1.222602e-13, 1.218117e-13, 1.219344e-13, 1.209565e-13, 1.205836e-13, 
    1.204246e-13, 1.202857e-13, 1.199472e-13, 1.20181e-13, 1.200888e-13, 
    1.203081e-13, 1.204473e-13, 1.203785e-13, 1.208031e-13, 1.206381e-13, 
    1.215063e-13, 1.211326e-13, 1.221061e-13, 1.218735e-13, 1.221618e-13, 
    1.220147e-13, 1.222667e-13, 1.2204e-13, 1.224327e-13, 1.225181e-13, 
    1.224597e-13, 1.22684e-13, 1.220274e-13, 1.222797e-13, 1.203765e-13, 
    1.203877e-13, 1.2044e-13, 1.2021e-13, 1.201959e-13, 1.19985e-13, 
    1.201727e-13, 1.202526e-13, 1.204554e-13, 1.205752e-13, 1.206891e-13, 
    1.209393e-13, 1.212185e-13, 1.216086e-13, 1.218885e-13, 1.22076e-13, 
    1.219611e-13, 1.220626e-13, 1.219491e-13, 1.21896e-13, 1.224861e-13, 
    1.221548e-13, 1.226518e-13, 1.226243e-13, 1.223995e-13, 1.226274e-13, 
    1.203956e-13, 1.20331e-13, 1.201065e-13, 1.202822e-13, 1.199621e-13, 
    1.201413e-13, 1.202443e-13, 1.206414e-13, 1.207287e-13, 1.208095e-13, 
    1.209691e-13, 1.211738e-13, 1.215325e-13, 1.218443e-13, 1.221287e-13, 
    1.221078e-13, 1.221152e-13, 1.221786e-13, 1.220214e-13, 1.222044e-13, 
    1.222351e-13, 1.221548e-13, 1.226206e-13, 1.224876e-13, 1.226237e-13, 
    1.225372e-13, 1.20352e-13, 1.204607e-13, 1.20402e-13, 1.205124e-13, 
    1.204346e-13, 1.207804e-13, 1.20884e-13, 1.213684e-13, 1.211698e-13, 
    1.214859e-13, 1.212019e-13, 1.212522e-13, 1.21496e-13, 1.212173e-13, 
    1.21827e-13, 1.214136e-13, 1.221811e-13, 1.217687e-13, 1.222069e-13, 
    1.221274e-13, 1.22259e-13, 1.223768e-13, 1.22525e-13, 1.227981e-13, 
    1.227349e-13, 1.229632e-13, 1.206227e-13, 1.207636e-13, 1.207512e-13, 
    1.208986e-13, 1.210075e-13, 1.212436e-13, 1.216217e-13, 1.214796e-13, 
    1.217405e-13, 1.217928e-13, 1.213964e-13, 1.216398e-13, 1.208578e-13, 
    1.209843e-13, 1.20909e-13, 1.206338e-13, 1.215122e-13, 1.210617e-13, 
    1.218932e-13, 1.216495e-13, 1.2236e-13, 1.220068e-13, 1.227001e-13, 
    1.229958e-13, 1.232741e-13, 1.235986e-13, 1.208405e-13, 1.207448e-13, 
    1.209161e-13, 1.211529e-13, 1.213726e-13, 1.216644e-13, 1.216942e-13, 
    1.217488e-13, 1.218903e-13, 1.220091e-13, 1.21766e-13, 1.220389e-13, 
    1.210134e-13, 1.215513e-13, 1.207086e-13, 1.209625e-13, 1.21139e-13, 
    1.210616e-13, 1.214633e-13, 1.215579e-13, 1.219419e-13, 1.217435e-13, 
    1.229228e-13, 1.224016e-13, 1.238457e-13, 1.234429e-13, 1.207114e-13, 
    1.208402e-13, 1.21288e-13, 1.21075e-13, 1.216839e-13, 1.218335e-13, 
    1.219552e-13, 1.221105e-13, 1.221273e-13, 1.222193e-13, 1.220685e-13, 
    1.222134e-13, 1.21665e-13, 1.219102e-13, 1.212369e-13, 1.214009e-13, 
    1.213255e-13, 1.212427e-13, 1.214981e-13, 1.217698e-13, 1.217757e-13, 
    1.218628e-13, 1.221078e-13, 1.216863e-13, 1.229898e-13, 1.221853e-13, 
    1.209806e-13, 1.212283e-13, 1.212638e-13, 1.211678e-13, 1.218185e-13, 
    1.215829e-13, 1.222171e-13, 1.220458e-13, 1.223264e-13, 1.22187e-13, 
    1.221665e-13, 1.219874e-13, 1.218758e-13, 1.215937e-13, 1.21364e-13, 
    1.211818e-13, 1.212242e-13, 1.214243e-13, 1.217865e-13, 1.221288e-13, 
    1.220538e-13, 1.223051e-13, 1.216398e-13, 1.219189e-13, 1.21811e-13, 
    1.220922e-13, 1.214758e-13, 1.220005e-13, 1.213415e-13, 1.213993e-13, 
    1.215782e-13, 1.219377e-13, 1.220173e-13, 1.221021e-13, 1.220498e-13, 
    1.217957e-13, 1.217541e-13, 1.215739e-13, 1.215241e-13, 1.213867e-13, 
    1.212729e-13, 1.213769e-13, 1.21486e-13, 1.217958e-13, 1.220747e-13, 
    1.223785e-13, 1.224528e-13, 1.22807e-13, 1.225186e-13, 1.229943e-13, 
    1.225897e-13, 1.232898e-13, 1.22031e-13, 1.22578e-13, 1.215864e-13, 
    1.216934e-13, 1.218868e-13, 1.2233e-13, 1.220909e-13, 1.223705e-13, 
    1.217524e-13, 1.214311e-13, 1.213481e-13, 1.211928e-13, 1.213516e-13, 
    1.213387e-13, 1.214906e-13, 1.214418e-13, 1.218061e-13, 1.216105e-13, 
    1.221659e-13, 1.223683e-13, 1.229393e-13, 1.232886e-13, 1.23644e-13, 
    1.238007e-13, 1.238483e-13, 1.238683e-13 ;

 LITR2C_vr =
  0.001107534, 0.001107533, 0.001107533, 0.001107532, 0.001107533, 
    0.001107532, 0.001107534, 0.001107533, 0.001107533, 0.001107534, 
    0.00110753, 0.001107532, 0.001107529, 0.00110753, 0.001107527, 
    0.001107529, 0.001107527, 0.001107527, 0.001107526, 0.001107526, 
    0.001107524, 0.001107526, 0.001107524, 0.001107525, 0.001107525, 
    0.001107526, 0.001107532, 0.001107531, 0.001107532, 0.001107532, 
    0.001107532, 0.001107533, 0.001107533, 0.001107534, 0.001107534, 
    0.001107533, 0.001107532, 0.001107532, 0.001107531, 0.001107531, 
    0.001107529, 0.00110753, 0.001107528, 0.001107528, 0.001107526, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107527, 
    0.001107527, 0.001107527, 0.00110753, 0.001107529, 0.001107531, 
    0.001107533, 0.001107534, 0.001107535, 0.001107534, 0.001107534, 
    0.001107533, 0.001107532, 0.001107532, 0.001107531, 0.001107531, 
    0.00110753, 0.001107529, 0.001107527, 0.001107528, 0.001107527, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107527, 
    0.001107526, 0.001107528, 0.001107527, 0.001107531, 0.001107532, 
    0.001107533, 0.001107533, 0.001107534, 0.001107533, 0.001107534, 
    0.001107533, 0.001107533, 0.001107533, 0.001107531, 0.001107532, 
    0.001107529, 0.00110753, 0.001107527, 0.001107528, 0.001107527, 
    0.001107527, 0.001107526, 0.001107527, 0.001107526, 0.001107525, 
    0.001107526, 0.001107525, 0.001107527, 0.001107526, 0.001107533, 
    0.001107533, 0.001107533, 0.001107533, 0.001107533, 0.001107534, 
    0.001107534, 0.001107533, 0.001107533, 0.001107532, 0.001107532, 
    0.001107531, 0.00110753, 0.001107529, 0.001107528, 0.001107527, 
    0.001107527, 0.001107527, 0.001107527, 0.001107528, 0.001107525, 
    0.001107527, 0.001107525, 0.001107525, 0.001107526, 0.001107525, 
    0.001107533, 0.001107533, 0.001107534, 0.001107533, 0.001107534, 
    0.001107534, 0.001107533, 0.001107532, 0.001107532, 0.001107531, 
    0.001107531, 0.00110753, 0.001107529, 0.001107528, 0.001107527, 
    0.001107527, 0.001107527, 0.001107526, 0.001107527, 0.001107526, 
    0.001107526, 0.001107527, 0.001107525, 0.001107525, 0.001107525, 
    0.001107525, 0.001107533, 0.001107533, 0.001107533, 0.001107532, 
    0.001107533, 0.001107531, 0.001107531, 0.001107529, 0.00110753, 
    0.001107529, 0.00110753, 0.00110753, 0.001107529, 0.00110753, 
    0.001107528, 0.001107529, 0.001107526, 0.001107528, 0.001107526, 
    0.001107527, 0.001107526, 0.001107526, 0.001107525, 0.001107524, 
    0.001107525, 0.001107524, 0.001107532, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.001107528, 0.001107529, 
    0.001107528, 0.001107528, 0.001107529, 0.001107528, 0.001107531, 
    0.001107531, 0.001107531, 0.001107532, 0.001107529, 0.00110753, 
    0.001107528, 0.001107528, 0.001107526, 0.001107527, 0.001107525, 
    0.001107524, 0.001107523, 0.001107522, 0.001107531, 0.001107531, 
    0.001107531, 0.00110753, 0.001107529, 0.001107528, 0.001107528, 
    0.001107528, 0.001107528, 0.001107527, 0.001107528, 0.001107527, 
    0.001107531, 0.001107529, 0.001107532, 0.001107531, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.001107527, 0.001107528, 
    0.001107524, 0.001107526, 0.001107521, 0.001107522, 0.001107532, 
    0.001107531, 0.00110753, 0.00110753, 0.001107528, 0.001107528, 
    0.001107527, 0.001107527, 0.001107527, 0.001107526, 0.001107527, 
    0.001107526, 0.001107528, 0.001107527, 0.00110753, 0.001107529, 
    0.00110753, 0.00110753, 0.001107529, 0.001107528, 0.001107528, 
    0.001107528, 0.001107527, 0.001107528, 0.001107524, 0.001107526, 
    0.001107531, 0.00110753, 0.00110753, 0.00110753, 0.001107528, 
    0.001107529, 0.001107526, 0.001107527, 0.001107526, 0.001107526, 
    0.001107527, 0.001107527, 0.001107528, 0.001107529, 0.001107529, 
    0.00110753, 0.00110753, 0.001107529, 0.001107528, 0.001107527, 
    0.001107527, 0.001107526, 0.001107528, 0.001107527, 0.001107528, 
    0.001107527, 0.001107529, 0.001107527, 0.00110753, 0.001107529, 
    0.001107529, 0.001107527, 0.001107527, 0.001107527, 0.001107527, 
    0.001107528, 0.001107528, 0.001107529, 0.001107529, 0.001107529, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107527, 
    0.001107526, 0.001107526, 0.001107524, 0.001107525, 0.001107524, 
    0.001107525, 0.001107523, 0.001107527, 0.001107525, 0.001107529, 
    0.001107528, 0.001107528, 0.001107526, 0.001107527, 0.001107526, 
    0.001107528, 0.001107529, 0.001107529, 0.00110753, 0.001107529, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107524, 0.001107523, 0.001107521, 
    0.001107521, 0.001107521, 0.001107521,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.68427e-07, 2.684267e-07, 2.684268e-07, 2.684265e-07, 2.684266e-07, 
    2.684265e-07, 2.684269e-07, 2.684267e-07, 2.684268e-07, 2.68427e-07, 
    2.684261e-07, 2.684265e-07, 2.684257e-07, 2.684259e-07, 2.684253e-07, 
    2.684257e-07, 2.684252e-07, 2.684253e-07, 2.68425e-07, 2.684251e-07, 
    2.684247e-07, 2.684249e-07, 2.684245e-07, 2.684247e-07, 2.684247e-07, 
    2.684249e-07, 2.684264e-07, 2.684262e-07, 2.684264e-07, 2.684264e-07, 
    2.684264e-07, 2.684266e-07, 2.684268e-07, 2.68427e-07, 2.68427e-07, 
    2.684268e-07, 2.684264e-07, 2.684265e-07, 2.684262e-07, 2.684262e-07, 
    2.684258e-07, 2.68426e-07, 2.684254e-07, 2.684256e-07, 2.684251e-07, 
    2.684252e-07, 2.684251e-07, 2.684251e-07, 2.684251e-07, 2.684252e-07, 
    2.684252e-07, 2.684253e-07, 2.68426e-07, 2.684258e-07, 2.684263e-07, 
    2.684267e-07, 2.684269e-07, 2.684271e-07, 2.68427e-07, 2.68427e-07, 
    2.684268e-07, 2.684266e-07, 2.684264e-07, 2.684263e-07, 2.684262e-07, 
    2.684259e-07, 2.684257e-07, 2.684253e-07, 2.684254e-07, 2.684253e-07, 
    2.684252e-07, 2.68425e-07, 2.68425e-07, 2.684249e-07, 2.684253e-07, 
    2.684251e-07, 2.684255e-07, 2.684253e-07, 2.684262e-07, 2.684265e-07, 
    2.684266e-07, 2.684267e-07, 2.68427e-07, 2.684268e-07, 2.684269e-07, 
    2.684267e-07, 2.684266e-07, 2.684267e-07, 2.684263e-07, 2.684264e-07, 
    2.684257e-07, 2.68426e-07, 2.684252e-07, 2.684254e-07, 2.684251e-07, 
    2.684253e-07, 2.684251e-07, 2.684253e-07, 2.684249e-07, 2.684249e-07, 
    2.684249e-07, 2.684247e-07, 2.684253e-07, 2.684251e-07, 2.684267e-07, 
    2.684266e-07, 2.684266e-07, 2.684268e-07, 2.684268e-07, 2.68427e-07, 
    2.684268e-07, 2.684268e-07, 2.684266e-07, 2.684265e-07, 2.684264e-07, 
    2.684262e-07, 2.684259e-07, 2.684256e-07, 2.684254e-07, 2.684252e-07, 
    2.684253e-07, 2.684252e-07, 2.684253e-07, 2.684254e-07, 2.684249e-07, 
    2.684252e-07, 2.684247e-07, 2.684248e-07, 2.684249e-07, 2.684248e-07, 
    2.684266e-07, 2.684267e-07, 2.684269e-07, 2.684267e-07, 2.68427e-07, 
    2.684269e-07, 2.684268e-07, 2.684264e-07, 2.684264e-07, 2.684263e-07, 
    2.684262e-07, 2.68426e-07, 2.684257e-07, 2.684254e-07, 2.684252e-07, 
    2.684252e-07, 2.684252e-07, 2.684251e-07, 2.684253e-07, 2.684251e-07, 
    2.684251e-07, 2.684252e-07, 2.684248e-07, 2.684249e-07, 2.684248e-07, 
    2.684248e-07, 2.684267e-07, 2.684266e-07, 2.684266e-07, 2.684266e-07, 
    2.684266e-07, 2.684263e-07, 2.684262e-07, 2.684258e-07, 2.68426e-07, 
    2.684257e-07, 2.68426e-07, 2.684259e-07, 2.684257e-07, 2.68426e-07, 
    2.684254e-07, 2.684258e-07, 2.684251e-07, 2.684255e-07, 2.684251e-07, 
    2.684252e-07, 2.684251e-07, 2.68425e-07, 2.684249e-07, 2.684246e-07, 
    2.684247e-07, 2.684245e-07, 2.684264e-07, 2.684263e-07, 2.684263e-07, 
    2.684262e-07, 2.684261e-07, 2.684259e-07, 2.684256e-07, 2.684257e-07, 
    2.684255e-07, 2.684255e-07, 2.684258e-07, 2.684256e-07, 2.684262e-07, 
    2.684261e-07, 2.684262e-07, 2.684264e-07, 2.684257e-07, 2.684261e-07, 
    2.684254e-07, 2.684256e-07, 2.68425e-07, 2.684253e-07, 2.684247e-07, 
    2.684245e-07, 2.684242e-07, 2.684239e-07, 2.684263e-07, 2.684264e-07, 
    2.684262e-07, 2.68426e-07, 2.684258e-07, 2.684256e-07, 2.684255e-07, 
    2.684255e-07, 2.684254e-07, 2.684253e-07, 2.684255e-07, 2.684253e-07, 
    2.684261e-07, 2.684257e-07, 2.684264e-07, 2.684262e-07, 2.68426e-07, 
    2.684261e-07, 2.684257e-07, 2.684257e-07, 2.684253e-07, 2.684255e-07, 
    2.684245e-07, 2.684249e-07, 2.684237e-07, 2.684241e-07, 2.684264e-07, 
    2.684263e-07, 2.684259e-07, 2.684261e-07, 2.684256e-07, 2.684254e-07, 
    2.684253e-07, 2.684252e-07, 2.684252e-07, 2.684251e-07, 2.684252e-07, 
    2.684251e-07, 2.684256e-07, 2.684254e-07, 2.684259e-07, 2.684258e-07, 
    2.684259e-07, 2.684259e-07, 2.684257e-07, 2.684255e-07, 2.684255e-07, 
    2.684254e-07, 2.684252e-07, 2.684256e-07, 2.684245e-07, 2.684251e-07, 
    2.684262e-07, 2.684259e-07, 2.684259e-07, 2.68426e-07, 2.684255e-07, 
    2.684257e-07, 2.684251e-07, 2.684253e-07, 2.68425e-07, 2.684251e-07, 
    2.684251e-07, 2.684253e-07, 2.684254e-07, 2.684256e-07, 2.684258e-07, 
    2.68426e-07, 2.684259e-07, 2.684258e-07, 2.684255e-07, 2.684252e-07, 
    2.684253e-07, 2.68425e-07, 2.684256e-07, 2.684254e-07, 2.684255e-07, 
    2.684252e-07, 2.684257e-07, 2.684253e-07, 2.684259e-07, 2.684258e-07, 
    2.684257e-07, 2.684253e-07, 2.684253e-07, 2.684252e-07, 2.684253e-07, 
    2.684255e-07, 2.684255e-07, 2.684257e-07, 2.684257e-07, 2.684258e-07, 
    2.684259e-07, 2.684258e-07, 2.684257e-07, 2.684255e-07, 2.684252e-07, 
    2.68425e-07, 2.684249e-07, 2.684246e-07, 2.684249e-07, 2.684245e-07, 
    2.684248e-07, 2.684242e-07, 2.684253e-07, 2.684248e-07, 2.684257e-07, 
    2.684255e-07, 2.684254e-07, 2.68425e-07, 2.684252e-07, 2.68425e-07, 
    2.684255e-07, 2.684258e-07, 2.684259e-07, 2.68426e-07, 2.684259e-07, 
    2.684259e-07, 2.684257e-07, 2.684258e-07, 2.684255e-07, 2.684256e-07, 
    2.684251e-07, 2.68425e-07, 2.684245e-07, 2.684242e-07, 2.684239e-07, 
    2.684238e-07, 2.684237e-07, 2.684237e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -3.921449e-26, 2.32836e-25, 1.56858e-25, 1.347998e-25, 1.715634e-26, 
    -5.391992e-26, 9.313441e-26, 6.862535e-26, 1.666616e-25, -1.078398e-25, 
    -1.740143e-25, -7.352717e-26, 1.911706e-25, 7.107626e-26, -3.063632e-25, 
    2.941087e-26, 2.450905e-26, 1.470543e-26, 1.495052e-25, -7.352717e-26, 
    2.573451e-25, 1.715634e-25, -9.803622e-26, -6.617445e-26, -1.397016e-25, 
    -2.450905e-26, 1.29898e-25, 2.132288e-25, 2.941087e-26, 4.41163e-26, 
    1.715634e-25, -2.450905e-26, -3.259704e-25, -4.41163e-26, -5.882173e-26, 
    3.186177e-26, 2.941087e-26, 1.127417e-25, 2.941087e-26, 7.352717e-27, 0, 
    -1.470543e-26, -2.671487e-25, -9.558531e-26, -6.127264e-26, 
    -3.431268e-26, 9.068351e-26, 3.357741e-25, 1.495052e-25, -1.470543e-26, 
    -1.715634e-26, 5.882173e-26, -3.186177e-26, -1.446034e-25, 1.764652e-25, 
    -9.803622e-27, -1.004871e-25, -7.842898e-26, -2.303851e-25, 2.695996e-26, 
    -2.205815e-25, 6.372354e-26, -2.622469e-25, -8.333079e-26, -1.593089e-25, 
    7.352717e-26, 2.401887e-25, 1.151926e-25, 1.29898e-25, -4.901811e-26, 
    2.499924e-25, -7.352717e-27, -3.186177e-26, -1.470543e-26, -1.715634e-26, 
    -6.372354e-26, 2.671487e-25, 1.617598e-25, 1.470543e-26, 5.882173e-26, 
    -1.200944e-25, -1.127417e-25, -2.818541e-25, 5.882173e-26, 1.274471e-25, 
    -6.127264e-26, -1.470543e-26, -2.156797e-25, -2.205815e-26, 
    -1.470543e-26, 2.843051e-25, 1.102908e-25, 2.450905e-26, 1.176435e-25, 
    4.901811e-27, 1.225453e-26, 9.803622e-26, -1.764652e-25, -4.901811e-27, 
    -8.82326e-26, -2.254833e-25, 1.715634e-26, 6.372354e-26, -2.279342e-25, 
    -4.166539e-26, -2.499924e-25, 2.205815e-26, 1.053889e-25, -1.02938e-25, 
    1.715634e-26, -1.985233e-25, -8.333079e-26, 2.058761e-25, 3.186177e-26, 
    -7.597807e-26, 9.558531e-26, 5.637083e-26, -4.901811e-26, -6.862535e-26, 
    -1.29898e-25, -5.146902e-26, -2.009742e-25, -6.372354e-26, 2.450905e-26, 
    1.495052e-25, -2.794032e-25, -1.127417e-25, -3.284213e-25, -7.107626e-26, 
    5.637083e-26, 1.470543e-26, -2.058761e-25, -5.146902e-26, -2.769523e-25, 
    8.333079e-26, 1.617598e-25, -8.578169e-26, -8.578169e-26, -4.901811e-26, 
    5.146902e-26, 2.377378e-25, -4.901811e-27, -1.274471e-25, 8.82326e-26, 
    -1.397016e-25, -7.352717e-27, 2.450906e-27, -7.597807e-26, 1.642107e-25, 
    -9.803622e-27, -2.671487e-25, 4.41163e-26, 2.181306e-25, 1.421525e-25, 
    8.82326e-26, -1.617598e-25, 3.186177e-26, -3.431268e-26, 1.347998e-25, 
    -2.450906e-27, -1.127417e-25, 3.431268e-26, -4.901811e-26, -1.397016e-25, 
    1.151926e-25, 2.450905e-26, -8.087988e-26, 7.842898e-26, 1.715634e-25, 
    -7.352717e-26, -6.862535e-26, 3.921449e-26, 4.41163e-26, -1.225453e-26, 
    2.695996e-26, -1.372507e-25, 7.352717e-26, 1.470543e-26, -1.102908e-25, 
    1.617598e-25, -6.372354e-26, 1.151926e-25, -2.941087e-26, 1.936215e-25, 
    1.519561e-25, 2.254833e-25, -3.186177e-26, -7.842898e-26, 1.936215e-25, 
    4.65672e-26, 8.333079e-26, -2.941087e-25, 1.666616e-25, -1.960724e-26, 
    9.068351e-26, -1.151926e-25, -2.695996e-26, -2.646978e-25, -2.034252e-25, 
    -7.597807e-26, 1.617598e-25, 2.08327e-25, 3.455777e-25, -3.431268e-26, 
    -1.200944e-25, -1.960724e-26, -3.921449e-26, 1.274471e-25, 2.843051e-25, 
    2.009742e-25, -3.186177e-26, -1.530638e-41, -3.186177e-26, -9.803622e-27, 
    3.676358e-26, -7.352717e-26, 1.715634e-26, -1.372507e-25, -3.063632e-25, 
    -3.431268e-26, -6.862535e-26, -4.901811e-26, -4.901811e-27, 
    -9.313441e-26, 1.200944e-25, 1.642107e-25, -1.666616e-25, -1.446034e-25, 
    -2.843051e-25, 2.377378e-25, 3.676358e-26, -9.313441e-26, -2.450906e-25, 
    -1.29898e-25, 2.230324e-25, -1.470543e-26, -2.058761e-25, 2.009742e-25, 
    2.132288e-25, -5.146902e-26, -2.695996e-26, -5.146902e-26, -1.495052e-25, 
    2.475414e-25, 2.009742e-25, -2.205815e-26, 3.186177e-26, -9.558531e-26, 
    -5.146902e-26, -3.676358e-26, -1.225453e-25, 2.548942e-25, -2.573451e-25, 
    -1.004871e-25, -2.034252e-25, 2.695996e-26, 4.901811e-27, -1.960724e-26, 
    8.82326e-26, -1.225453e-26, 7.597807e-26, -1.372507e-25, 7.842898e-26, 
    -9.803622e-27, -3.11265e-25, -6.372354e-26, -1.81367e-25, 8.578169e-26, 
    -2.32836e-25, -1.54407e-25, -3.186177e-26, 4.41163e-26, -8.087988e-26, 
    9.068351e-26, -3.676358e-26, -2.499924e-25, 1.691125e-25, 1.740143e-25, 
    1.960724e-26, -1.421525e-25, -1.911706e-25, -7.597807e-26, 1.593089e-25, 
    -7.597807e-26, 1.666616e-25, -7.842898e-26, 5.882173e-26, 7.107626e-26, 
    -3.676358e-26, -1.691125e-25, 1.642107e-25, -4.901811e-26, -1.470543e-26, 
    -3.431268e-26, -1.740143e-25, -4.166539e-26, 1.960724e-26, 2.843051e-25, 
    9.803622e-27, 1.053889e-25, -1.225453e-25, 1.470543e-25, -5.391992e-26, 
    -1.54407e-25, -5.882173e-26, -6.862535e-26, -1.004871e-25, 6.862535e-26, 
    -2.205815e-26, 6.372354e-26, 1.715634e-26, -2.941087e-26, 1.176435e-25, 
    -2.59796e-25, 2.450906e-25, 1.151926e-25, 7.352717e-27, 1.862688e-25, 
    -1.642107e-25, 5.391992e-26, -9.068351e-26, 6.372354e-26, -7.842898e-26, 
    1.078398e-25, -3.186177e-26, 2.450906e-27, 4.41163e-26, -3.431268e-25, 
    -2.450905e-26, -4.65672e-26, -2.034252e-25, 1.372507e-25, 4.166539e-26, 
    -1.421525e-25, 2.205815e-26, 2.156797e-25, -1.740143e-25, 1.960724e-26,
  2.676256e-32, 2.676253e-32, 2.676254e-32, 2.676252e-32, 2.676253e-32, 
    2.676251e-32, 2.676255e-32, 2.676253e-32, 2.676254e-32, 2.676256e-32, 
    2.676247e-32, 2.676252e-32, 2.676243e-32, 2.676245e-32, 2.676239e-32, 
    2.676243e-32, 2.676238e-32, 2.676239e-32, 2.676236e-32, 2.676237e-32, 
    2.676233e-32, 2.676235e-32, 2.676231e-32, 2.676233e-32, 2.676233e-32, 
    2.676235e-32, 2.676251e-32, 2.676248e-32, 2.676251e-32, 2.67625e-32, 
    2.676251e-32, 2.676253e-32, 2.676254e-32, 2.676256e-32, 2.676256e-32, 
    2.676254e-32, 2.67625e-32, 2.676252e-32, 2.676248e-32, 2.676248e-32, 
    2.676244e-32, 2.676246e-32, 2.67624e-32, 2.676242e-32, 2.676237e-32, 
    2.676238e-32, 2.676237e-32, 2.676237e-32, 2.676237e-32, 2.676239e-32, 
    2.676238e-32, 2.676239e-32, 2.676246e-32, 2.676244e-32, 2.67625e-32, 
    2.676253e-32, 2.676255e-32, 2.676257e-32, 2.676257e-32, 2.676256e-32, 
    2.676254e-32, 2.676252e-32, 2.67625e-32, 2.676249e-32, 2.676248e-32, 
    2.676245e-32, 2.676243e-32, 2.676239e-32, 2.67624e-32, 2.676239e-32, 
    2.676238e-32, 2.676236e-32, 2.676237e-32, 2.676236e-32, 2.676239e-32, 
    2.676237e-32, 2.676241e-32, 2.676239e-32, 2.676248e-32, 2.676251e-32, 
    2.676252e-32, 2.676254e-32, 2.676257e-32, 2.676254e-32, 2.676255e-32, 
    2.676254e-32, 2.676252e-32, 2.676253e-32, 2.676249e-32, 2.676251e-32, 
    2.676243e-32, 2.676247e-32, 2.676238e-32, 2.67624e-32, 2.676238e-32, 
    2.676239e-32, 2.676237e-32, 2.676239e-32, 2.676235e-32, 2.676235e-32, 
    2.676235e-32, 2.676233e-32, 2.676239e-32, 2.676237e-32, 2.676253e-32, 
    2.676253e-32, 2.676252e-32, 2.676254e-32, 2.676254e-32, 2.676256e-32, 
    2.676254e-32, 2.676254e-32, 2.676252e-32, 2.676251e-32, 2.67625e-32, 
    2.676248e-32, 2.676246e-32, 2.676242e-32, 2.67624e-32, 2.676238e-32, 
    2.676239e-32, 2.676239e-32, 2.676239e-32, 2.67624e-32, 2.676235e-32, 
    2.676238e-32, 2.676234e-32, 2.676234e-32, 2.676236e-32, 2.676234e-32, 
    2.676253e-32, 2.676253e-32, 2.676255e-32, 2.676254e-32, 2.676257e-32, 
    2.676255e-32, 2.676254e-32, 2.676251e-32, 2.67625e-32, 2.676249e-32, 
    2.676248e-32, 2.676246e-32, 2.676243e-32, 2.67624e-32, 2.676238e-32, 
    2.676238e-32, 2.676238e-32, 2.676237e-32, 2.676239e-32, 2.676237e-32, 
    2.676237e-32, 2.676238e-32, 2.676234e-32, 2.676235e-32, 2.676234e-32, 
    2.676234e-32, 2.676253e-32, 2.676252e-32, 2.676253e-32, 2.676252e-32, 
    2.676252e-32, 2.676249e-32, 2.676249e-32, 2.676244e-32, 2.676246e-32, 
    2.676243e-32, 2.676246e-32, 2.676245e-32, 2.676243e-32, 2.676246e-32, 
    2.676241e-32, 2.676244e-32, 2.676237e-32, 2.676241e-32, 2.676237e-32, 
    2.676238e-32, 2.676237e-32, 2.676236e-32, 2.676234e-32, 2.676232e-32, 
    2.676233e-32, 2.676231e-32, 2.676251e-32, 2.676249e-32, 2.67625e-32, 
    2.676248e-32, 2.676247e-32, 2.676245e-32, 2.676242e-32, 2.676244e-32, 
    2.676241e-32, 2.676241e-32, 2.676244e-32, 2.676242e-32, 2.676249e-32, 
    2.676248e-32, 2.676248e-32, 2.676251e-32, 2.676243e-32, 2.676247e-32, 
    2.67624e-32, 2.676242e-32, 2.676236e-32, 2.676239e-32, 2.676233e-32, 
    2.676231e-32, 2.676228e-32, 2.676225e-32, 2.676249e-32, 2.67625e-32, 
    2.676248e-32, 2.676246e-32, 2.676244e-32, 2.676242e-32, 2.676242e-32, 
    2.676241e-32, 2.67624e-32, 2.676239e-32, 2.676241e-32, 2.676239e-32, 
    2.676247e-32, 2.676243e-32, 2.67625e-32, 2.676248e-32, 2.676246e-32, 
    2.676247e-32, 2.676244e-32, 2.676243e-32, 2.676239e-32, 2.676241e-32, 
    2.676231e-32, 2.676236e-32, 2.676223e-32, 2.676227e-32, 2.67625e-32, 
    2.676249e-32, 2.676245e-32, 2.676247e-32, 2.676242e-32, 2.67624e-32, 
    2.676239e-32, 2.676238e-32, 2.676238e-32, 2.676237e-32, 2.676239e-32, 
    2.676237e-32, 2.676242e-32, 2.67624e-32, 2.676246e-32, 2.676244e-32, 
    2.676245e-32, 2.676245e-32, 2.676243e-32, 2.676241e-32, 2.676241e-32, 
    2.67624e-32, 2.676238e-32, 2.676242e-32, 2.676231e-32, 2.676237e-32, 
    2.676248e-32, 2.676246e-32, 2.676245e-32, 2.676246e-32, 2.676241e-32, 
    2.676243e-32, 2.676237e-32, 2.676239e-32, 2.676236e-32, 2.676237e-32, 
    2.676238e-32, 2.676239e-32, 2.67624e-32, 2.676242e-32, 2.676244e-32, 
    2.676246e-32, 2.676246e-32, 2.676244e-32, 2.676241e-32, 2.676238e-32, 
    2.676239e-32, 2.676237e-32, 2.676242e-32, 2.67624e-32, 2.676241e-32, 
    2.676238e-32, 2.676244e-32, 2.676239e-32, 2.676245e-32, 2.676244e-32, 
    2.676243e-32, 2.676239e-32, 2.676239e-32, 2.676238e-32, 2.676239e-32, 
    2.676241e-32, 2.676241e-32, 2.676243e-32, 2.676243e-32, 2.676244e-32, 
    2.676245e-32, 2.676244e-32, 2.676243e-32, 2.676241e-32, 2.676238e-32, 
    2.676236e-32, 2.676235e-32, 2.676232e-32, 2.676235e-32, 2.676231e-32, 
    2.676234e-32, 2.676228e-32, 2.676239e-32, 2.676234e-32, 2.676243e-32, 
    2.676242e-32, 2.67624e-32, 2.676236e-32, 2.676238e-32, 2.676236e-32, 
    2.676241e-32, 2.676244e-32, 2.676244e-32, 2.676246e-32, 2.676244e-32, 
    2.676245e-32, 2.676243e-32, 2.676244e-32, 2.676241e-32, 2.676242e-32, 
    2.676238e-32, 2.676236e-32, 2.676231e-32, 2.676228e-32, 2.676225e-32, 
    2.676224e-32, 2.676223e-32, 2.676223e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.321735e-15, 3.330745e-15, 3.328995e-15, 3.336256e-15, 3.33223e-15, 
    3.336982e-15, 3.323564e-15, 3.331102e-15, 3.326291e-15, 3.322548e-15, 
    3.350325e-15, 3.33658e-15, 3.364591e-15, 3.35584e-15, 3.377808e-15, 
    3.363228e-15, 3.380745e-15, 3.377391e-15, 3.38749e-15, 3.384598e-15, 
    3.397496e-15, 3.388824e-15, 3.404178e-15, 3.395427e-15, 3.396796e-15, 
    3.388538e-15, 3.33935e-15, 3.348615e-15, 3.338801e-15, 3.340122e-15, 
    3.33953e-15, 3.332312e-15, 3.328671e-15, 3.321048e-15, 3.322433e-15, 
    3.328032e-15, 3.340717e-15, 3.336415e-15, 3.347258e-15, 3.347014e-15, 
    3.359067e-15, 3.353635e-15, 3.37387e-15, 3.368125e-15, 3.384719e-15, 
    3.380549e-15, 3.384523e-15, 3.383318e-15, 3.384538e-15, 3.378421e-15, 
    3.381043e-15, 3.375659e-15, 3.354652e-15, 3.36083e-15, 3.342388e-15, 
    3.331276e-15, 3.323894e-15, 3.31865e-15, 3.319391e-15, 3.320805e-15, 
    3.328065e-15, 3.334888e-15, 3.340084e-15, 3.343557e-15, 3.346978e-15, 
    3.357318e-15, 3.362792e-15, 3.37503e-15, 3.372825e-15, 3.376562e-15, 
    3.380134e-15, 3.386123e-15, 3.385138e-15, 3.387775e-15, 3.376465e-15, 
    3.383983e-15, 3.371569e-15, 3.374966e-15, 3.347899e-15, 3.337576e-15, 
    3.333177e-15, 3.329331e-15, 3.319962e-15, 3.326433e-15, 3.323882e-15, 
    3.329951e-15, 3.333804e-15, 3.331899e-15, 3.343652e-15, 3.339084e-15, 
    3.363116e-15, 3.352773e-15, 3.379717e-15, 3.373278e-15, 3.38126e-15, 
    3.377189e-15, 3.384163e-15, 3.377887e-15, 3.388757e-15, 3.391121e-15, 
    3.389506e-15, 3.395713e-15, 3.377538e-15, 3.384522e-15, 3.331845e-15, 
    3.332155e-15, 3.333604e-15, 3.327236e-15, 3.326847e-15, 3.32101e-15, 
    3.326204e-15, 3.328415e-15, 3.334028e-15, 3.337344e-15, 3.340496e-15, 
    3.347423e-15, 3.35515e-15, 3.365947e-15, 3.373696e-15, 3.378885e-15, 
    3.375704e-15, 3.378513e-15, 3.375373e-15, 3.373901e-15, 3.390235e-15, 
    3.381066e-15, 3.394821e-15, 3.394061e-15, 3.387838e-15, 3.394146e-15, 
    3.332374e-15, 3.330586e-15, 3.324372e-15, 3.329235e-15, 3.320374e-15, 
    3.325334e-15, 3.328184e-15, 3.339178e-15, 3.341593e-15, 3.34383e-15, 
    3.348248e-15, 3.353913e-15, 3.363841e-15, 3.372471e-15, 3.380342e-15, 
    3.379765e-15, 3.379968e-15, 3.381725e-15, 3.377372e-15, 3.382439e-15, 
    3.383288e-15, 3.381066e-15, 3.393959e-15, 3.390278e-15, 3.394045e-15, 
    3.391648e-15, 3.331167e-15, 3.334176e-15, 3.33255e-15, 3.335607e-15, 
    3.333453e-15, 3.343024e-15, 3.345891e-15, 3.359298e-15, 3.353801e-15, 
    3.362551e-15, 3.354691e-15, 3.356083e-15, 3.362832e-15, 3.355116e-15, 
    3.371993e-15, 3.360551e-15, 3.381793e-15, 3.370378e-15, 3.382508e-15, 
    3.380308e-15, 3.383951e-15, 3.387211e-15, 3.391312e-15, 3.398872e-15, 
    3.397122e-15, 3.403441e-15, 3.33866e-15, 3.342558e-15, 3.342217e-15, 
    3.346296e-15, 3.349311e-15, 3.355844e-15, 3.366309e-15, 3.362375e-15, 
    3.369597e-15, 3.371045e-15, 3.360075e-15, 3.366811e-15, 3.345168e-15, 
    3.348666e-15, 3.346585e-15, 3.338967e-15, 3.36328e-15, 3.35081e-15, 
    3.373823e-15, 3.367079e-15, 3.386746e-15, 3.37697e-15, 3.396159e-15, 
    3.404343e-15, 3.412046e-15, 3.421029e-15, 3.344687e-15, 3.342039e-15, 
    3.346781e-15, 3.353335e-15, 3.359416e-15, 3.367491e-15, 3.368317e-15, 
    3.369828e-15, 3.373744e-15, 3.377033e-15, 3.370305e-15, 3.377858e-15, 
    3.349474e-15, 3.364362e-15, 3.341036e-15, 3.348065e-15, 3.352949e-15, 
    3.350809e-15, 3.361926e-15, 3.364544e-15, 3.375172e-15, 3.369681e-15, 
    3.402322e-15, 3.387897e-15, 3.427867e-15, 3.416717e-15, 3.341113e-15, 
    3.344679e-15, 3.357073e-15, 3.351178e-15, 3.36803e-15, 3.372172e-15, 
    3.375539e-15, 3.379838e-15, 3.380304e-15, 3.38285e-15, 3.378677e-15, 
    3.382686e-15, 3.367508e-15, 3.374294e-15, 3.35566e-15, 3.360198e-15, 
    3.358111e-15, 3.35582e-15, 3.362889e-15, 3.37041e-15, 3.370574e-15, 
    3.372983e-15, 3.379765e-15, 3.368099e-15, 3.404177e-15, 3.381911e-15, 
    3.348565e-15, 3.355421e-15, 3.356403e-15, 3.353748e-15, 3.371757e-15, 
    3.365236e-15, 3.382788e-15, 3.378049e-15, 3.385814e-15, 3.381956e-15, 
    3.381388e-15, 3.376431e-15, 3.373342e-15, 3.365534e-15, 3.359177e-15, 
    3.354133e-15, 3.355307e-15, 3.360846e-15, 3.370871e-15, 3.380345e-15, 
    3.37827e-15, 3.385224e-15, 3.36681e-15, 3.374535e-15, 3.371549e-15, 
    3.379333e-15, 3.36227e-15, 3.376794e-15, 3.358553e-15, 3.360155e-15, 
    3.365106e-15, 3.375057e-15, 3.377261e-15, 3.379608e-15, 3.37816e-15, 
    3.371125e-15, 3.369974e-15, 3.364987e-15, 3.363608e-15, 3.359806e-15, 
    3.356656e-15, 3.359533e-15, 3.362554e-15, 3.37113e-15, 3.378849e-15, 
    3.387257e-15, 3.389314e-15, 3.399118e-15, 3.391135e-15, 3.4043e-15, 
    3.393103e-15, 3.412479e-15, 3.377639e-15, 3.392779e-15, 3.365333e-15, 
    3.368294e-15, 3.373646e-15, 3.385913e-15, 3.379296e-15, 3.387036e-15, 
    3.369929e-15, 3.361035e-15, 3.358736e-15, 3.35444e-15, 3.358834e-15, 
    3.358477e-15, 3.362681e-15, 3.36133e-15, 3.371414e-15, 3.365999e-15, 
    3.381373e-15, 3.386975e-15, 3.402778e-15, 3.412448e-15, 3.422284e-15, 
    3.426621e-15, 3.42794e-15, 3.428492e-15 ;

 LITR2N_vr =
  1.532746e-05, 1.532744e-05, 1.532744e-05, 1.532743e-05, 1.532744e-05, 
    1.532743e-05, 1.532745e-05, 1.532744e-05, 1.532745e-05, 1.532746e-05, 
    1.532741e-05, 1.532743e-05, 1.532738e-05, 1.53274e-05, 1.532736e-05, 
    1.532738e-05, 1.532735e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 
    1.532732e-05, 1.532734e-05, 1.532731e-05, 1.532733e-05, 1.532733e-05, 
    1.532734e-05, 1.532743e-05, 1.532741e-05, 1.532743e-05, 1.532742e-05, 
    1.532743e-05, 1.532744e-05, 1.532744e-05, 1.532746e-05, 1.532746e-05, 
    1.532745e-05, 1.532742e-05, 1.532743e-05, 1.532741e-05, 1.532741e-05, 
    1.532739e-05, 1.53274e-05, 1.532737e-05, 1.532738e-05, 1.532735e-05, 
    1.532735e-05, 1.532735e-05, 1.532735e-05, 1.532735e-05, 1.532736e-05, 
    1.532735e-05, 1.532736e-05, 1.53274e-05, 1.532739e-05, 1.532742e-05, 
    1.532744e-05, 1.532745e-05, 1.532746e-05, 1.532746e-05, 1.532746e-05, 
    1.532745e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 1.532741e-05, 
    1.53274e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532734e-05, 1.532735e-05, 1.532734e-05, 1.532736e-05, 
    1.532735e-05, 1.532737e-05, 1.532736e-05, 1.532741e-05, 1.532743e-05, 
    1.532744e-05, 1.532744e-05, 1.532746e-05, 1.532745e-05, 1.532745e-05, 
    1.532744e-05, 1.532744e-05, 1.532744e-05, 1.532742e-05, 1.532743e-05, 
    1.532738e-05, 1.53274e-05, 1.532736e-05, 1.532737e-05, 1.532735e-05, 
    1.532736e-05, 1.532735e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532736e-05, 1.532735e-05, 1.532744e-05, 
    1.532744e-05, 1.532744e-05, 1.532745e-05, 1.532745e-05, 1.532746e-05, 
    1.532745e-05, 1.532744e-05, 1.532744e-05, 1.532743e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532738e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532736e-05, 1.532737e-05, 1.532734e-05, 
    1.532735e-05, 1.532733e-05, 1.532733e-05, 1.532734e-05, 1.532733e-05, 
    1.532744e-05, 1.532744e-05, 1.532745e-05, 1.532744e-05, 1.532746e-05, 
    1.532745e-05, 1.532745e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532738e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532736e-05, 1.532735e-05, 
    1.532735e-05, 1.532735e-05, 1.532733e-05, 1.532734e-05, 1.532733e-05, 
    1.532734e-05, 1.532744e-05, 1.532744e-05, 1.532744e-05, 1.532743e-05, 
    1.532744e-05, 1.532742e-05, 1.532742e-05, 1.532739e-05, 1.53274e-05, 
    1.532739e-05, 1.53274e-05, 1.53274e-05, 1.532738e-05, 1.53274e-05, 
    1.532737e-05, 1.532739e-05, 1.532735e-05, 1.532737e-05, 1.532735e-05, 
    1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532734e-05, 1.532732e-05, 
    1.532732e-05, 1.532731e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.53274e-05, 1.532738e-05, 1.532739e-05, 
    1.532737e-05, 1.532737e-05, 1.532739e-05, 1.532738e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.532743e-05, 1.532738e-05, 1.532741e-05, 
    1.532737e-05, 1.532738e-05, 1.532734e-05, 1.532736e-05, 1.532733e-05, 
    1.532731e-05, 1.53273e-05, 1.532728e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 1.532738e-05, 
    1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532737e-05, 1.532736e-05, 
    1.532741e-05, 1.532738e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 
    1.532741e-05, 1.532739e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532732e-05, 1.532734e-05, 1.532727e-05, 1.532729e-05, 1.532742e-05, 
    1.532742e-05, 1.53274e-05, 1.532741e-05, 1.532738e-05, 1.532737e-05, 
    1.532736e-05, 1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532736e-05, 
    1.532735e-05, 1.532738e-05, 1.532736e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.53274e-05, 1.532738e-05, 1.532737e-05, 1.532737e-05, 
    1.532737e-05, 1.532736e-05, 1.532738e-05, 1.532731e-05, 1.532735e-05, 
    1.532741e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 1.532737e-05, 
    1.532738e-05, 1.532735e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 
    1.532735e-05, 1.532736e-05, 1.532737e-05, 1.532738e-05, 1.532739e-05, 
    1.53274e-05, 1.53274e-05, 1.532739e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532735e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532736e-05, 1.532739e-05, 1.532736e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532736e-05, 1.532736e-05, 1.532736e-05, 1.532736e-05, 
    1.532737e-05, 1.532737e-05, 1.532738e-05, 1.532738e-05, 1.532739e-05, 
    1.53274e-05, 1.532739e-05, 1.532739e-05, 1.532737e-05, 1.532736e-05, 
    1.532734e-05, 1.532734e-05, 1.532732e-05, 1.532734e-05, 1.532731e-05, 
    1.532733e-05, 1.53273e-05, 1.532736e-05, 1.532733e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532734e-05, 1.532736e-05, 1.532734e-05, 
    1.532737e-05, 1.532739e-05, 1.532739e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.532739e-05, 1.532739e-05, 1.532737e-05, 1.532738e-05, 
    1.532735e-05, 1.532734e-05, 1.532732e-05, 1.53273e-05, 1.532728e-05, 
    1.532727e-05, 1.532727e-05, 1.532727e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.200113e-13, 1.203368e-13, 1.202736e-13, 1.205359e-13, 1.203904e-13, 
    1.205621e-13, 1.200773e-13, 1.203497e-13, 1.201759e-13, 1.200406e-13, 
    1.210442e-13, 1.205476e-13, 1.215596e-13, 1.212434e-13, 1.220371e-13, 
    1.215104e-13, 1.221432e-13, 1.22022e-13, 1.223869e-13, 1.222824e-13, 
    1.227484e-13, 1.224351e-13, 1.229898e-13, 1.226737e-13, 1.227231e-13, 
    1.224248e-13, 1.206477e-13, 1.209824e-13, 1.206278e-13, 1.206756e-13, 
    1.206542e-13, 1.203934e-13, 1.202618e-13, 1.199864e-13, 1.200365e-13, 
    1.202388e-13, 1.20697e-13, 1.205416e-13, 1.209334e-13, 1.209245e-13, 
    1.2136e-13, 1.211638e-13, 1.218949e-13, 1.216873e-13, 1.222868e-13, 
    1.221361e-13, 1.222797e-13, 1.222362e-13, 1.222803e-13, 1.220593e-13, 
    1.22154e-13, 1.219595e-13, 1.212005e-13, 1.214237e-13, 1.207574e-13, 
    1.20356e-13, 1.200893e-13, 1.198998e-13, 1.199266e-13, 1.199776e-13, 
    1.202399e-13, 1.204865e-13, 1.206742e-13, 1.207997e-13, 1.209233e-13, 
    1.212969e-13, 1.214946e-13, 1.219368e-13, 1.218571e-13, 1.219921e-13, 
    1.221211e-13, 1.223375e-13, 1.223019e-13, 1.223972e-13, 1.219886e-13, 
    1.222602e-13, 1.218117e-13, 1.219344e-13, 1.209565e-13, 1.205836e-13, 
    1.204246e-13, 1.202857e-13, 1.199472e-13, 1.20181e-13, 1.200888e-13, 
    1.203081e-13, 1.204473e-13, 1.203785e-13, 1.208031e-13, 1.206381e-13, 
    1.215063e-13, 1.211326e-13, 1.221061e-13, 1.218735e-13, 1.221618e-13, 
    1.220147e-13, 1.222667e-13, 1.2204e-13, 1.224327e-13, 1.225181e-13, 
    1.224597e-13, 1.22684e-13, 1.220274e-13, 1.222797e-13, 1.203765e-13, 
    1.203877e-13, 1.2044e-13, 1.2021e-13, 1.201959e-13, 1.19985e-13, 
    1.201727e-13, 1.202526e-13, 1.204554e-13, 1.205752e-13, 1.206891e-13, 
    1.209393e-13, 1.212185e-13, 1.216086e-13, 1.218885e-13, 1.22076e-13, 
    1.219611e-13, 1.220626e-13, 1.219491e-13, 1.21896e-13, 1.224861e-13, 
    1.221548e-13, 1.226518e-13, 1.226243e-13, 1.223995e-13, 1.226274e-13, 
    1.203956e-13, 1.20331e-13, 1.201065e-13, 1.202822e-13, 1.199621e-13, 
    1.201413e-13, 1.202443e-13, 1.206414e-13, 1.207287e-13, 1.208095e-13, 
    1.209691e-13, 1.211738e-13, 1.215325e-13, 1.218443e-13, 1.221287e-13, 
    1.221078e-13, 1.221152e-13, 1.221786e-13, 1.220214e-13, 1.222044e-13, 
    1.222351e-13, 1.221548e-13, 1.226206e-13, 1.224876e-13, 1.226237e-13, 
    1.225372e-13, 1.20352e-13, 1.204607e-13, 1.20402e-13, 1.205124e-13, 
    1.204346e-13, 1.207804e-13, 1.20884e-13, 1.213684e-13, 1.211698e-13, 
    1.214859e-13, 1.212019e-13, 1.212522e-13, 1.21496e-13, 1.212173e-13, 
    1.21827e-13, 1.214136e-13, 1.221811e-13, 1.217687e-13, 1.222069e-13, 
    1.221274e-13, 1.22259e-13, 1.223768e-13, 1.22525e-13, 1.227981e-13, 
    1.227349e-13, 1.229632e-13, 1.206227e-13, 1.207636e-13, 1.207512e-13, 
    1.208986e-13, 1.210075e-13, 1.212436e-13, 1.216217e-13, 1.214796e-13, 
    1.217405e-13, 1.217928e-13, 1.213964e-13, 1.216398e-13, 1.208578e-13, 
    1.209843e-13, 1.20909e-13, 1.206338e-13, 1.215122e-13, 1.210617e-13, 
    1.218932e-13, 1.216495e-13, 1.2236e-13, 1.220068e-13, 1.227001e-13, 
    1.229958e-13, 1.232741e-13, 1.235986e-13, 1.208405e-13, 1.207448e-13, 
    1.209161e-13, 1.211529e-13, 1.213726e-13, 1.216644e-13, 1.216942e-13, 
    1.217488e-13, 1.218903e-13, 1.220091e-13, 1.21766e-13, 1.220389e-13, 
    1.210134e-13, 1.215513e-13, 1.207086e-13, 1.209625e-13, 1.21139e-13, 
    1.210616e-13, 1.214633e-13, 1.215579e-13, 1.219419e-13, 1.217435e-13, 
    1.229228e-13, 1.224016e-13, 1.238457e-13, 1.234429e-13, 1.207114e-13, 
    1.208402e-13, 1.21288e-13, 1.21075e-13, 1.216839e-13, 1.218335e-13, 
    1.219552e-13, 1.221105e-13, 1.221273e-13, 1.222193e-13, 1.220685e-13, 
    1.222134e-13, 1.21665e-13, 1.219102e-13, 1.212369e-13, 1.214009e-13, 
    1.213255e-13, 1.212427e-13, 1.214981e-13, 1.217698e-13, 1.217757e-13, 
    1.218628e-13, 1.221078e-13, 1.216863e-13, 1.229898e-13, 1.221853e-13, 
    1.209806e-13, 1.212283e-13, 1.212638e-13, 1.211678e-13, 1.218185e-13, 
    1.215829e-13, 1.222171e-13, 1.220458e-13, 1.223264e-13, 1.22187e-13, 
    1.221665e-13, 1.219874e-13, 1.218758e-13, 1.215937e-13, 1.21364e-13, 
    1.211818e-13, 1.212242e-13, 1.214243e-13, 1.217865e-13, 1.221288e-13, 
    1.220538e-13, 1.223051e-13, 1.216398e-13, 1.219189e-13, 1.21811e-13, 
    1.220922e-13, 1.214758e-13, 1.220005e-13, 1.213415e-13, 1.213993e-13, 
    1.215782e-13, 1.219377e-13, 1.220173e-13, 1.221021e-13, 1.220498e-13, 
    1.217957e-13, 1.217541e-13, 1.215739e-13, 1.215241e-13, 1.213867e-13, 
    1.212729e-13, 1.213769e-13, 1.21486e-13, 1.217958e-13, 1.220747e-13, 
    1.223785e-13, 1.224528e-13, 1.22807e-13, 1.225186e-13, 1.229943e-13, 
    1.225897e-13, 1.232898e-13, 1.22031e-13, 1.22578e-13, 1.215864e-13, 
    1.216934e-13, 1.218868e-13, 1.2233e-13, 1.220909e-13, 1.223705e-13, 
    1.217524e-13, 1.214311e-13, 1.213481e-13, 1.211928e-13, 1.213516e-13, 
    1.213387e-13, 1.214906e-13, 1.214418e-13, 1.218061e-13, 1.216105e-13, 
    1.221659e-13, 1.223683e-13, 1.229393e-13, 1.232886e-13, 1.23644e-13, 
    1.238007e-13, 1.238483e-13, 1.238683e-13 ;

 LITR3C =
  9.698018e-06, 9.698008e-06, 9.69801e-06, 9.698002e-06, 9.698007e-06, 
    9.698002e-06, 9.698017e-06, 9.698008e-06, 9.698014e-06, 9.698017e-06, 
    9.697987e-06, 9.698002e-06, 9.697971e-06, 9.697981e-06, 9.697957e-06, 
    9.697973e-06, 9.697953e-06, 9.697957e-06, 9.697946e-06, 9.697949e-06, 
    9.697935e-06, 9.697945e-06, 9.697927e-06, 9.697937e-06, 9.697936e-06, 
    9.697945e-06, 9.697999e-06, 9.697988e-06, 9.697999e-06, 9.697998e-06, 
    9.697999e-06, 9.698007e-06, 9.698011e-06, 9.698019e-06, 9.698017e-06, 
    9.698011e-06, 9.697997e-06, 9.698002e-06, 9.69799e-06, 9.69799e-06, 
    9.697977e-06, 9.697983e-06, 9.697961e-06, 9.697967e-06, 9.697949e-06, 
    9.697954e-06, 9.697949e-06, 9.69795e-06, 9.697949e-06, 9.697956e-06, 
    9.697953e-06, 9.697959e-06, 9.697982e-06, 9.697976e-06, 9.697996e-06, 
    9.698008e-06, 9.698016e-06, 9.698022e-06, 9.698021e-06, 9.698019e-06, 
    9.698011e-06, 9.698004e-06, 9.697998e-06, 9.697995e-06, 9.69799e-06, 
    9.697979e-06, 9.697973e-06, 9.697959e-06, 9.697962e-06, 9.697958e-06, 
    9.697954e-06, 9.697947e-06, 9.697948e-06, 9.697946e-06, 9.697958e-06, 
    9.69795e-06, 9.697964e-06, 9.69796e-06, 9.697989e-06, 9.698001e-06, 
    9.698006e-06, 9.69801e-06, 9.69802e-06, 9.698013e-06, 9.698017e-06, 
    9.698009e-06, 9.698005e-06, 9.698007e-06, 9.697995e-06, 9.697999e-06, 
    9.697973e-06, 9.697984e-06, 9.697955e-06, 9.697962e-06, 9.697953e-06, 
    9.697957e-06, 9.697949e-06, 9.697957e-06, 9.697945e-06, 9.697942e-06, 
    9.697944e-06, 9.697937e-06, 9.697957e-06, 9.697949e-06, 9.698007e-06, 
    9.698007e-06, 9.698006e-06, 9.698012e-06, 9.698013e-06, 9.698019e-06, 
    9.698014e-06, 9.698011e-06, 9.698005e-06, 9.698001e-06, 9.697997e-06, 
    9.69799e-06, 9.697982e-06, 9.697969e-06, 9.697961e-06, 9.697956e-06, 
    9.697959e-06, 9.697956e-06, 9.697959e-06, 9.697961e-06, 9.697943e-06, 
    9.697953e-06, 9.697937e-06, 9.697938e-06, 9.697946e-06, 9.697938e-06, 
    9.698007e-06, 9.698008e-06, 9.698016e-06, 9.69801e-06, 9.69802e-06, 
    9.698015e-06, 9.698011e-06, 9.697999e-06, 9.697997e-06, 9.697994e-06, 
    9.697989e-06, 9.697983e-06, 9.697972e-06, 9.697963e-06, 9.697954e-06, 
    9.697955e-06, 9.697954e-06, 9.697952e-06, 9.697957e-06, 9.697951e-06, 
    9.69795e-06, 9.697953e-06, 9.697938e-06, 9.697943e-06, 9.697938e-06, 
    9.697941e-06, 9.698008e-06, 9.698005e-06, 9.698007e-06, 9.698003e-06, 
    9.698006e-06, 9.697995e-06, 9.697992e-06, 9.697977e-06, 9.697983e-06, 
    9.697974e-06, 9.697982e-06, 9.69798e-06, 9.697973e-06, 9.697982e-06, 
    9.697963e-06, 9.697976e-06, 9.697952e-06, 9.697965e-06, 9.697951e-06, 
    9.697954e-06, 9.69795e-06, 9.697947e-06, 9.697942e-06, 9.697933e-06, 
    9.697936e-06, 9.697928e-06, 9.698e-06, 9.697996e-06, 9.697996e-06, 
    9.697991e-06, 9.697988e-06, 9.697981e-06, 9.697969e-06, 9.697974e-06, 
    9.697966e-06, 9.697964e-06, 9.697977e-06, 9.697968e-06, 9.697993e-06, 
    9.697988e-06, 9.697991e-06, 9.697999e-06, 9.697973e-06, 9.697987e-06, 
    9.697961e-06, 9.697968e-06, 9.697947e-06, 9.697957e-06, 9.697937e-06, 
    9.697927e-06, 9.697918e-06, 9.697909e-06, 9.697993e-06, 9.697996e-06, 
    9.697991e-06, 9.697984e-06, 9.697977e-06, 9.697968e-06, 9.697967e-06, 
    9.697966e-06, 9.697961e-06, 9.697957e-06, 9.697965e-06, 9.697957e-06, 
    9.697987e-06, 9.697971e-06, 9.697997e-06, 9.697989e-06, 9.697984e-06, 
    9.697987e-06, 9.697974e-06, 9.697971e-06, 9.697959e-06, 9.697966e-06, 
    9.697929e-06, 9.697946e-06, 9.697901e-06, 9.697914e-06, 9.697997e-06, 
    9.697993e-06, 9.697979e-06, 9.697986e-06, 9.697967e-06, 9.697963e-06, 
    9.697959e-06, 9.697955e-06, 9.697954e-06, 9.697951e-06, 9.697956e-06, 
    9.697951e-06, 9.697968e-06, 9.69796e-06, 9.697981e-06, 9.697976e-06, 
    9.697978e-06, 9.697981e-06, 9.697973e-06, 9.697965e-06, 9.697965e-06, 
    9.697962e-06, 9.697955e-06, 9.697967e-06, 9.697927e-06, 9.697952e-06, 
    9.697989e-06, 9.697981e-06, 9.69798e-06, 9.697983e-06, 9.697963e-06, 
    9.69797e-06, 9.697951e-06, 9.697957e-06, 9.697947e-06, 9.697952e-06, 
    9.697953e-06, 9.697958e-06, 9.697961e-06, 9.69797e-06, 9.697977e-06, 
    9.697983e-06, 9.697981e-06, 9.697976e-06, 9.697964e-06, 9.697954e-06, 
    9.697956e-06, 9.697948e-06, 9.697968e-06, 9.69796e-06, 9.697964e-06, 
    9.697955e-06, 9.697974e-06, 9.697957e-06, 9.697977e-06, 9.697976e-06, 
    9.69797e-06, 9.697959e-06, 9.697957e-06, 9.697955e-06, 9.697957e-06, 
    9.697964e-06, 9.697966e-06, 9.697971e-06, 9.697972e-06, 9.697977e-06, 
    9.69798e-06, 9.697977e-06, 9.697974e-06, 9.697964e-06, 9.697956e-06, 
    9.697947e-06, 9.697944e-06, 9.697933e-06, 9.697942e-06, 9.697927e-06, 
    9.697939e-06, 9.697918e-06, 9.697957e-06, 9.69794e-06, 9.69797e-06, 
    9.697967e-06, 9.697961e-06, 9.697947e-06, 9.697955e-06, 9.697947e-06, 
    9.697966e-06, 9.697975e-06, 9.697977e-06, 9.697982e-06, 9.697977e-06, 
    9.697978e-06, 9.697973e-06, 9.697975e-06, 9.697964e-06, 9.697969e-06, 
    9.697953e-06, 9.697947e-06, 9.697929e-06, 9.697918e-06, 9.697907e-06, 
    9.697903e-06, 9.697901e-06, 9.697901e-06 ;

 LITR3C_TO_SOIL2C =
  6.000561e-14, 6.016838e-14, 6.013676e-14, 6.026792e-14, 6.01952e-14, 
    6.028104e-14, 6.003864e-14, 6.017481e-14, 6.008791e-14, 6.00203e-14, 
    6.052208e-14, 6.027377e-14, 6.077978e-14, 6.06217e-14, 6.101855e-14, 
    6.075516e-14, 6.10716e-14, 6.1011e-14, 6.119344e-14, 6.11412e-14, 
    6.13742e-14, 6.121755e-14, 6.14949e-14, 6.133683e-14, 6.136155e-14, 
    6.121237e-14, 6.032382e-14, 6.049118e-14, 6.031389e-14, 6.033777e-14, 
    6.032706e-14, 6.019668e-14, 6.01309e-14, 5.99932e-14, 6.001821e-14, 
    6.011937e-14, 6.034851e-14, 6.027079e-14, 6.046667e-14, 6.046226e-14, 
    6.068e-14, 6.058186e-14, 6.094741e-14, 6.084362e-14, 6.114339e-14, 
    6.106805e-14, 6.113984e-14, 6.111808e-14, 6.114013e-14, 6.102962e-14, 
    6.107697e-14, 6.097971e-14, 6.060023e-14, 6.071185e-14, 6.03787e-14, 
    6.017796e-14, 6.004461e-14, 5.994987e-14, 5.996327e-14, 5.99888e-14, 
    6.011996e-14, 6.024322e-14, 6.033707e-14, 6.039982e-14, 6.046162e-14, 
    6.064841e-14, 6.074729e-14, 6.096836e-14, 6.092854e-14, 6.099604e-14, 
    6.106055e-14, 6.116875e-14, 6.115095e-14, 6.119859e-14, 6.099429e-14, 
    6.113009e-14, 6.090583e-14, 6.09672e-14, 6.047825e-14, 6.029177e-14, 
    6.02123e-14, 6.014283e-14, 5.997357e-14, 6.009047e-14, 6.004439e-14, 
    6.015402e-14, 6.022362e-14, 6.018921e-14, 6.040153e-14, 6.031901e-14, 
    6.075314e-14, 6.05663e-14, 6.105303e-14, 6.093672e-14, 6.10809e-14, 
    6.100735e-14, 6.113334e-14, 6.101996e-14, 6.121633e-14, 6.125904e-14, 
    6.122986e-14, 6.134199e-14, 6.101367e-14, 6.113982e-14, 6.018824e-14, 
    6.019385e-14, 6.022001e-14, 6.010498e-14, 6.009795e-14, 5.99925e-14, 
    6.008635e-14, 6.012627e-14, 6.022767e-14, 6.028758e-14, 6.034452e-14, 
    6.046965e-14, 6.060924e-14, 6.080427e-14, 6.094425e-14, 6.1038e-14, 
    6.098054e-14, 6.103127e-14, 6.097455e-14, 6.094796e-14, 6.124303e-14, 
    6.10774e-14, 6.132587e-14, 6.131214e-14, 6.119972e-14, 6.131369e-14, 
    6.019779e-14, 6.016549e-14, 6.005324e-14, 6.014109e-14, 5.998102e-14, 
    6.007062e-14, 6.012211e-14, 6.03207e-14, 6.036434e-14, 6.040475e-14, 
    6.048455e-14, 6.058688e-14, 6.076623e-14, 6.092212e-14, 6.106431e-14, 
    6.10539e-14, 6.105756e-14, 6.10893e-14, 6.101067e-14, 6.110221e-14, 
    6.111755e-14, 6.10774e-14, 6.13103e-14, 6.12438e-14, 6.131184e-14, 
    6.126856e-14, 6.0176e-14, 6.023034e-14, 6.020098e-14, 6.025619e-14, 
    6.021728e-14, 6.039018e-14, 6.044198e-14, 6.068416e-14, 6.058486e-14, 
    6.074292e-14, 6.060094e-14, 6.06261e-14, 6.074801e-14, 6.060862e-14, 
    6.09135e-14, 6.070681e-14, 6.109053e-14, 6.088431e-14, 6.110344e-14, 
    6.10637e-14, 6.112951e-14, 6.11884e-14, 6.126249e-14, 6.139905e-14, 
    6.136744e-14, 6.14816e-14, 6.031135e-14, 6.038177e-14, 6.03756e-14, 
    6.044929e-14, 6.050375e-14, 6.062176e-14, 6.081082e-14, 6.073976e-14, 
    6.087021e-14, 6.089638e-14, 6.06982e-14, 6.081988e-14, 6.04289e-14, 
    6.049211e-14, 6.04545e-14, 6.031689e-14, 6.075609e-14, 6.053084e-14, 
    6.094656e-14, 6.082474e-14, 6.118e-14, 6.10034e-14, 6.135003e-14, 
    6.149789e-14, 6.163704e-14, 6.17993e-14, 6.042022e-14, 6.037239e-14, 
    6.045805e-14, 6.057644e-14, 6.068629e-14, 6.083216e-14, 6.08471e-14, 
    6.087439e-14, 6.094512e-14, 6.100455e-14, 6.088299e-14, 6.101944e-14, 
    6.05067e-14, 6.077565e-14, 6.035427e-14, 6.048124e-14, 6.056948e-14, 
    6.053081e-14, 6.073165e-14, 6.077894e-14, 6.097092e-14, 6.087172e-14, 
    6.146138e-14, 6.120079e-14, 6.192283e-14, 6.172141e-14, 6.035566e-14, 
    6.042007e-14, 6.064398e-14, 6.053749e-14, 6.084191e-14, 6.091673e-14, 
    6.097756e-14, 6.105523e-14, 6.106363e-14, 6.110963e-14, 6.103424e-14, 
    6.110666e-14, 6.083248e-14, 6.095507e-14, 6.061844e-14, 6.070042e-14, 
    6.066272e-14, 6.062133e-14, 6.074903e-14, 6.08849e-14, 6.088785e-14, 
    6.093138e-14, 6.105389e-14, 6.084315e-14, 6.149488e-14, 6.109265e-14, 
    6.049028e-14, 6.061413e-14, 6.063187e-14, 6.05839e-14, 6.090923e-14, 
    6.079143e-14, 6.110851e-14, 6.10229e-14, 6.116316e-14, 6.109347e-14, 
    6.108321e-14, 6.099366e-14, 6.093787e-14, 6.079683e-14, 6.068198e-14, 
    6.059087e-14, 6.061206e-14, 6.071212e-14, 6.089322e-14, 6.106437e-14, 
    6.102689e-14, 6.115251e-14, 6.081986e-14, 6.095941e-14, 6.090548e-14, 
    6.104608e-14, 6.073786e-14, 6.100022e-14, 6.067071e-14, 6.069964e-14, 
    6.078909e-14, 6.096884e-14, 6.100865e-14, 6.105106e-14, 6.10249e-14, 
    6.089783e-14, 6.087702e-14, 6.078693e-14, 6.076202e-14, 6.069335e-14, 
    6.063644e-14, 6.068842e-14, 6.074298e-14, 6.08979e-14, 6.103734e-14, 
    6.118923e-14, 6.12264e-14, 6.140349e-14, 6.125928e-14, 6.149711e-14, 
    6.129483e-14, 6.164486e-14, 6.101548e-14, 6.128898e-14, 6.079318e-14, 
    6.084669e-14, 6.094336e-14, 6.116496e-14, 6.104542e-14, 6.118524e-14, 
    6.08762e-14, 6.071555e-14, 6.067402e-14, 6.05964e-14, 6.06758e-14, 
    6.066934e-14, 6.074527e-14, 6.072088e-14, 6.090304e-14, 6.080522e-14, 
    6.108295e-14, 6.118414e-14, 6.146962e-14, 6.164431e-14, 6.182198e-14, 
    6.190031e-14, 6.192415e-14, 6.193412e-14 ;

 LITR3C_vr =
  0.0005537669, 0.0005537663, 0.0005537664, 0.000553766, 0.0005537662, 
    0.0005537659, 0.0005537668, 0.0005537663, 0.0005537666, 0.0005537668, 
    0.0005537651, 0.0005537659, 0.0005537642, 0.0005537648, 0.0005537634, 
    0.0005537643, 0.0005537632, 0.0005537634, 0.0005537627, 0.0005537629, 
    0.0005537621, 0.0005537627, 0.0005537617, 0.0005537622, 0.0005537621, 
    0.0005537627, 0.0005537657, 0.0005537652, 0.0005537658, 0.0005537657, 
    0.0005537657, 0.0005537662, 0.0005537664, 0.0005537669, 0.0005537668, 
    0.0005537665, 0.0005537657, 0.000553766, 0.0005537653, 0.0005537653, 
    0.0005537645, 0.0005537649, 0.0005537636, 0.0005537639, 0.0005537629, 
    0.0005537632, 0.0005537629, 0.000553763, 0.0005537629, 0.0005537633, 
    0.0005537631, 0.0005537635, 0.0005537648, 0.0005537644, 0.0005537656, 
    0.0005537663, 0.0005537667, 0.0005537671, 0.000553767, 0.000553767, 
    0.0005537665, 0.000553766, 0.0005537657, 0.0005537655, 0.0005537653, 
    0.0005537646, 0.0005537643, 0.0005537635, 0.0005537636, 0.0005537634, 
    0.0005537632, 0.0005537628, 0.0005537629, 0.0005537627, 0.0005537634, 
    0.0005537629, 0.0005537638, 0.0005537635, 0.0005537652, 0.0005537659, 
    0.0005537661, 0.0005537664, 0.000553767, 0.0005537666, 0.0005537667, 
    0.0005537664, 0.0005537661, 0.0005537663, 0.0005537655, 0.0005537658, 
    0.0005537643, 0.0005537649, 0.0005537632, 0.0005537636, 0.0005537631, 
    0.0005537634, 0.0005537629, 0.0005537634, 0.0005537627, 0.0005537625, 
    0.0005537626, 0.0005537622, 0.0005537634, 0.0005537629, 0.0005537663, 
    0.0005537662, 0.0005537661, 0.0005537666, 0.0005537666, 0.0005537669, 
    0.0005537666, 0.0005537664, 0.0005537661, 0.0005537659, 0.0005537657, 
    0.0005537653, 0.0005537648, 0.0005537641, 0.0005537636, 0.0005537633, 
    0.0005537635, 0.0005537633, 0.0005537635, 0.0005537636, 0.0005537625, 
    0.0005537631, 0.0005537622, 0.0005537623, 0.0005537627, 0.0005537623, 
    0.0005537662, 0.0005537663, 0.0005537667, 0.0005537664, 0.000553767, 
    0.0005537667, 0.0005537665, 0.0005537658, 0.0005537656, 0.0005537655, 
    0.0005537652, 0.0005537649, 0.0005537642, 0.0005537637, 0.0005537632, 
    0.0005537632, 0.0005537632, 0.0005537631, 0.0005537634, 0.0005537631, 
    0.000553763, 0.0005537631, 0.0005537623, 0.0005537625, 0.0005537623, 
    0.0005537625, 0.0005537663, 0.0005537661, 0.0005537662, 0.000553766, 
    0.0005537661, 0.0005537655, 0.0005537653, 0.0005537645, 0.0005537649, 
    0.0005537643, 0.0005537648, 0.0005537647, 0.0005537643, 0.0005537648, 
    0.0005537637, 0.0005537644, 0.0005537631, 0.0005537638, 0.0005537631, 
    0.0005537632, 0.0005537629, 0.0005537628, 0.0005537625, 0.000553762, 
    0.0005537621, 0.0005537617, 0.0005537658, 0.0005537656, 0.0005537656, 
    0.0005537653, 0.0005537652, 0.0005537648, 0.0005537641, 0.0005537643, 
    0.0005537639, 0.0005537638, 0.0005537645, 0.0005537641, 0.0005537654, 
    0.0005537652, 0.0005537653, 0.0005537658, 0.0005537643, 0.000553765, 
    0.0005537636, 0.000553764, 0.0005537628, 0.0005537634, 0.0005537622, 
    0.0005537617, 0.0005537612, 0.0005537606, 0.0005537655, 0.0005537656, 
    0.0005537653, 0.0005537649, 0.0005537645, 0.000553764, 0.0005537639, 
    0.0005537638, 0.0005537636, 0.0005537634, 0.0005537638, 0.0005537634, 
    0.0005537651, 0.0005537642, 0.0005537657, 0.0005537652, 0.0005537649, 
    0.000553765, 0.0005537643, 0.0005537642, 0.0005537635, 0.0005537639, 
    0.0005537618, 0.0005537627, 0.0005537602, 0.0005537609, 0.0005537657, 
    0.0005537655, 0.0005537646, 0.000553765, 0.0005537639, 0.0005537637, 
    0.0005537635, 0.0005537632, 0.0005537632, 0.000553763, 0.0005537633, 
    0.0005537631, 0.000553764, 0.0005537636, 0.0005537648, 0.0005537645, 
    0.0005537646, 0.0005537648, 0.0005537643, 0.0005537638, 0.0005537638, 
    0.0005537636, 0.0005537632, 0.0005537639, 0.0005537617, 0.0005537631, 
    0.0005537652, 0.0005537648, 0.0005537647, 0.0005537649, 0.0005537637, 
    0.0005537641, 0.000553763, 0.0005537634, 0.0005537628, 0.0005537631, 
    0.0005537631, 0.0005537634, 0.0005537636, 0.0005537641, 0.0005537645, 
    0.0005537648, 0.0005537648, 0.0005537644, 0.0005537638, 0.0005537632, 
    0.0005537633, 0.0005537629, 0.0005537641, 0.0005537635, 0.0005537638, 
    0.0005537632, 0.0005537643, 0.0005537634, 0.0005537646, 0.0005537645, 
    0.0005537642, 0.0005537635, 0.0005537634, 0.0005537632, 0.0005537633, 
    0.0005537638, 0.0005537638, 0.0005537642, 0.0005537642, 0.0005537645, 
    0.0005537647, 0.0005537645, 0.0005537643, 0.0005537638, 0.0005537633, 
    0.0005537628, 0.0005537626, 0.000553762, 0.0005537625, 0.0005537617, 
    0.0005537624, 0.0005537611, 0.0005537634, 0.0005537624, 0.0005537641, 
    0.0005537639, 0.0005537636, 0.0005537628, 0.0005537632, 0.0005537628, 
    0.0005537638, 0.0005537644, 0.0005537645, 0.0005537648, 0.0005537645, 
    0.0005537646, 0.0005537643, 0.0005537644, 0.0005537638, 0.0005537641, 
    0.0005537631, 0.0005537628, 0.0005537618, 0.0005537611, 0.0005537606, 
    0.0005537603, 0.0005537602, 0.0005537602,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342135e-07, 1.342133e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342133e-07, 1.342135e-07, 1.342133e-07, 1.342134e-07, 1.342135e-07, 
    1.34213e-07, 1.342133e-07, 1.342128e-07, 1.34213e-07, 1.342126e-07, 
    1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342125e-07, 1.342125e-07, 
    1.342123e-07, 1.342125e-07, 1.342122e-07, 1.342124e-07, 1.342123e-07, 
    1.342125e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342132e-07, 1.342133e-07, 1.342134e-07, 1.342135e-07, 1.342135e-07, 
    1.342134e-07, 1.342132e-07, 1.342133e-07, 1.342131e-07, 1.342131e-07, 
    1.342129e-07, 1.34213e-07, 1.342127e-07, 1.342128e-07, 1.342125e-07, 
    1.342126e-07, 1.342125e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 
    1.342126e-07, 1.342127e-07, 1.34213e-07, 1.342129e-07, 1.342132e-07, 
    1.342133e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 1.342135e-07, 
    1.342134e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 
    1.342129e-07, 1.342129e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342125e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 
    1.342125e-07, 1.342127e-07, 1.342127e-07, 1.342131e-07, 1.342132e-07, 
    1.342133e-07, 1.342134e-07, 1.342135e-07, 1.342134e-07, 1.342135e-07, 
    1.342134e-07, 1.342133e-07, 1.342133e-07, 1.342131e-07, 1.342132e-07, 
    1.342129e-07, 1.34213e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342125e-07, 1.342126e-07, 1.342125e-07, 1.342124e-07, 
    1.342124e-07, 1.342123e-07, 1.342126e-07, 1.342125e-07, 1.342133e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 1.342135e-07, 
    1.342134e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 
    1.342127e-07, 1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342124e-07, 
    1.342126e-07, 1.342124e-07, 1.342124e-07, 1.342125e-07, 1.342124e-07, 
    1.342133e-07, 1.342134e-07, 1.342134e-07, 1.342134e-07, 1.342135e-07, 
    1.342134e-07, 1.342134e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.34213e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 
    1.342125e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 1.342124e-07, 
    1.342124e-07, 1.342133e-07, 1.342133e-07, 1.342133e-07, 1.342133e-07, 
    1.342133e-07, 1.342132e-07, 1.342131e-07, 1.342129e-07, 1.34213e-07, 
    1.342129e-07, 1.34213e-07, 1.34213e-07, 1.342129e-07, 1.34213e-07, 
    1.342127e-07, 1.342129e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342125e-07, 1.342125e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342132e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342128e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342129e-07, 1.342128e-07, 1.342131e-07, 
    1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342128e-07, 1.34213e-07, 
    1.342127e-07, 1.342128e-07, 1.342125e-07, 1.342126e-07, 1.342123e-07, 
    1.342122e-07, 1.342121e-07, 1.34212e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342131e-07, 1.342128e-07, 1.342132e-07, 1.342131e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342127e-07, 
    1.342122e-07, 1.342125e-07, 1.342119e-07, 1.34212e-07, 1.342132e-07, 
    1.342131e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 
    1.342125e-07, 1.342128e-07, 1.342127e-07, 1.34213e-07, 1.342129e-07, 
    1.342129e-07, 1.34213e-07, 1.342129e-07, 1.342127e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342128e-07, 1.342122e-07, 1.342126e-07, 
    1.342131e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 1.342127e-07, 
    1.342128e-07, 1.342125e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342127e-07, 1.342128e-07, 1.342129e-07, 
    1.34213e-07, 1.34213e-07, 1.342129e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342125e-07, 1.342128e-07, 1.342127e-07, 1.342127e-07, 
    1.342126e-07, 1.342129e-07, 1.342126e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342128e-07, 1.342128e-07, 1.342129e-07, 
    1.342129e-07, 1.342129e-07, 1.342129e-07, 1.342127e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 
    1.342124e-07, 1.342121e-07, 1.342126e-07, 1.342124e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342126e-07, 1.342125e-07, 
    1.342127e-07, 1.342129e-07, 1.342129e-07, 1.34213e-07, 1.342129e-07, 
    1.342129e-07, 1.342129e-07, 1.342129e-07, 1.342127e-07, 1.342128e-07, 
    1.342126e-07, 1.342125e-07, 1.342122e-07, 1.342121e-07, 1.342119e-07, 
    1.342119e-07, 1.342119e-07, 1.342118e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  6.4949e-26, 9.068351e-26, 8.700715e-26, 9.435986e-26, -5.637083e-26, 
    3.921449e-26, -3.798904e-26, -4.901811e-27, -4.901811e-26, 2.450906e-27, 
    3.676358e-26, -8.700715e-26, -9.558531e-26, 9.558531e-26, 2.818541e-26, 
    3.921449e-26, -9.803622e-27, -2.818541e-26, -4.166539e-26, 9.803622e-27, 
    1.02938e-25, -1.286725e-25, 3.553813e-26, -9.803622e-26, 5.759628e-26, 
    -5.391992e-26, 1.102908e-26, 9.190896e-26, -2.818541e-26, -1.102908e-26, 
    7.230172e-26, -1.580834e-25, -2.941087e-26, -2.32836e-26, -2.08327e-26, 
    -2.08327e-26, -2.941087e-26, -1.446034e-25, 1.838179e-26, 1.249962e-25, 
    4.901811e-26, -2.205815e-26, 1.715634e-26, 4.289085e-26, 8.455624e-26, 
    2.941087e-26, -5.514538e-26, -1.102908e-26, 3.798904e-26, 3.308722e-26, 
    9.803622e-27, 2.450905e-26, -3.308722e-26, -8.087988e-26, -4.41163e-26, 
    1.225453e-27, -1.225453e-27, -4.779266e-26, 7.597807e-26, -8.82326e-26, 
    -5.637083e-26, -7.352717e-27, 3.553813e-26, 7.230172e-26, 2.205815e-26, 
    -9.190896e-26, -6.862535e-26, -7.352717e-26, 1.715634e-26, -1.593089e-26, 
    -4.534175e-26, -1.16418e-25, 5.514538e-26, -5.146902e-26, 2.32836e-26, 
    -4.779266e-26, -4.043994e-26, 2.450906e-27, -3.063632e-26, 2.450906e-27, 
    -1.347998e-26, -7.230172e-26, -2.205815e-26, 5.391992e-26, -8.210533e-26, 
    7.597807e-26, 1.139671e-25, -1.470543e-26, 3.431268e-26, 1.102908e-26, 
    8.945805e-26, -2.573451e-26, -6.004719e-26, -1.225453e-27, 1.470543e-26, 
    -5.269447e-26, -1.102908e-25, 1.470543e-26, -6.617445e-26, 4.901811e-27, 
    5.882173e-26, -1.801416e-25, 2.32836e-26, -1.078398e-25, -1.629852e-25, 
    -5.637083e-26, -6.73999e-26, 4.534175e-26, 8.210533e-26, -2.941087e-26, 
    -2.450905e-26, 4.779266e-26, -7.107626e-26, 9.926167e-26, -1.225453e-26, 
    9.435986e-26, -7.720352e-26, -5.882173e-26, -2.573451e-26, 7.352717e-27, 
    1.102908e-26, -1.470543e-26, -7.352717e-27, -9.803622e-27, -8.578169e-26, 
    -5.637083e-26, 2.818541e-26, 7.597807e-26, -9.190896e-26, -3.186177e-26, 
    -1.715634e-26, 1.960724e-26, 2.695996e-26, 7.107626e-26, 1.593089e-26, 
    4.166539e-26, -1.102908e-26, -1.347998e-26, -7.230172e-26, 3.308722e-26, 
    1.56858e-25, 4.043994e-26, -2.450906e-27, 2.450905e-26, 1.715634e-26, 
    4.901811e-27, 1.960724e-26, -5.269447e-26, -6.4949e-26, -4.779266e-26, 
    -7.352717e-27, -6.249809e-26, 5.146902e-26, -9.190896e-26, 1.16418e-25, 
    -6.862535e-26, 4.41163e-26, 3.431268e-26, -6.127264e-27, 5.391992e-26, 
    -4.65672e-26, -2.450905e-26, 1.874943e-25, 1.004871e-25, 7.652491e-42, 
    1.225453e-27, -2.205815e-26, 4.65672e-26, -3.921449e-26, -3.676358e-27, 
    1.225453e-27, -7.352717e-27, 2.818541e-26, 2.818541e-26, 4.289085e-26, 
    7.107626e-26, -1.960724e-26, -3.063632e-26, 9.435986e-26, -7.107626e-26, 
    6.862535e-26, 4.534175e-26, 8.700715e-26, 6.73999e-26, -2.818541e-26, 
    -6.127264e-27, 1.225453e-26, -4.65672e-26, -6.862535e-26, 1.02938e-25, 
    6.372354e-26, 1.593089e-26, -3.308722e-26, -3.431268e-26, -2.941087e-26, 
    2.450905e-26, 1.470543e-26, 1.519561e-25, -1.960724e-26, -6.127264e-27, 
    -8.700715e-26, 3.431268e-26, 2.695996e-26, -7.842898e-26, 1.004871e-25, 
    -7.720352e-26, 7.475262e-26, -1.960724e-26, -1.495052e-25, -1.237707e-25, 
    -1.225453e-27, -5.024356e-26, -1.127417e-25, -3.063632e-26, 
    -4.166539e-26, -8.82326e-26, -2.32836e-26, 1.02938e-25, -1.102908e-25, 
    1.593089e-26, 5.637083e-26, 9.803622e-27, -2.475414e-25, -2.08327e-26, 
    -9.803622e-27, -8.945805e-26, 1.347998e-26, -1.041635e-25, -4.289085e-26, 
    6.127264e-27, -2.32836e-26, 7.720352e-26, -3.431268e-26, 1.715634e-26, 
    1.139671e-25, 1.960724e-26, -1.960724e-26, 2.818541e-26, -9.435986e-26, 
    -6.862535e-26, -1.507307e-25, 0, 3.676358e-26, 3.921449e-26, 
    -8.578169e-27, -4.166539e-26, -1.102908e-25, -1.311234e-25, 
    -1.593089e-26, -1.715634e-26, 2.941087e-26, 8.82326e-26, -8.945805e-26, 
    1.715634e-26, 7.597807e-26, 6.372354e-26, -2.818541e-26, -1.066144e-25, 
    -3.063632e-26, -7.230172e-26, -1.225453e-27, -9.435986e-26, 8.087988e-26, 
    -2.941087e-26, -1.16418e-25, -4.289085e-26, 2.450906e-27, -2.695996e-26, 
    2.32836e-26, 1.02938e-25, 2.205815e-26, -1.004871e-25, -3.798904e-26, 
    1.02938e-25, -3.798904e-26, -4.901811e-26, 8.578169e-27, 4.41163e-26, 
    3.308722e-26, 7.352717e-27, 1.838179e-26, 6.127264e-27, 1.225453e-27, 
    -1.200944e-25, 1.078398e-25, 4.166539e-26, -6.4949e-26, -8.578169e-26, 
    3.676358e-27, -2.034252e-25, 4.901811e-26, -8.455624e-26, 3.921449e-26, 
    -6.617445e-26, -5.391992e-26, 4.534175e-26, -2.08327e-26, 1.115162e-25, 
    1.225453e-27, 1.715634e-26, 5.146902e-26, -1.151926e-25, 6.127264e-27, 
    -3.676358e-27, -1.838179e-26, -1.225453e-27, -3.676358e-27, 2.818541e-26, 
    -1.470543e-26, 4.779266e-26, 2.32836e-26, 8.700715e-26, -1.225453e-27, 
    -1.249962e-25, -1.16418e-25, -4.289085e-26, -3.553813e-26, -1.593089e-26, 
    2.32836e-26, 4.534175e-26, -1.789161e-25, -5.637083e-26, 6.98508e-26, 
    -1.225453e-27, 1.838179e-26, 2.32836e-26, -2.450906e-27, -2.941087e-26, 
    1.347998e-26, 8.210533e-26, -2.695996e-26, -2.818541e-26, -6.4949e-26, 
    9.190896e-26, 1.470543e-26, -1.347998e-26, -7.352717e-27, -9.681077e-26,
  1.338128e-32, 1.338126e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338126e-32, 1.338128e-32, 1.338126e-32, 1.338127e-32, 1.338128e-32, 
    1.338124e-32, 1.338126e-32, 1.338121e-32, 1.338123e-32, 1.338119e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338118e-32, 1.338118e-32, 
    1.338116e-32, 1.338118e-32, 1.338115e-32, 1.338117e-32, 1.338116e-32, 
    1.338118e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338125e-32, 1.338126e-32, 1.338127e-32, 1.338128e-32, 1.338128e-32, 
    1.338127e-32, 1.338125e-32, 1.338126e-32, 1.338124e-32, 1.338124e-32, 
    1.338122e-32, 1.338123e-32, 1.33812e-32, 1.338121e-32, 1.338118e-32, 
    1.338119e-32, 1.338118e-32, 1.338118e-32, 1.338118e-32, 1.338119e-32, 
    1.338119e-32, 1.33812e-32, 1.338123e-32, 1.338122e-32, 1.338125e-32, 
    1.338126e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 1.338128e-32, 
    1.338127e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 
    1.338123e-32, 1.338122e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338118e-32, 1.338118e-32, 1.338118e-32, 1.338119e-32, 
    1.338118e-32, 1.33812e-32, 1.33812e-32, 1.338124e-32, 1.338125e-32, 
    1.338126e-32, 1.338127e-32, 1.338128e-32, 1.338127e-32, 1.338128e-32, 
    1.338127e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 
    1.338121e-32, 1.338123e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338118e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338118e-32, 1.338117e-32, 1.338119e-32, 1.338118e-32, 1.338126e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 1.338128e-32, 
    1.338127e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 
    1.33812e-32, 1.338119e-32, 1.33812e-32, 1.33812e-32, 1.338117e-32, 
    1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338117e-32, 
    1.338126e-32, 1.338126e-32, 1.338128e-32, 1.338127e-32, 1.338128e-32, 
    1.338127e-32, 1.338127e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 
    1.338118e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 
    1.338117e-32, 1.338126e-32, 1.338126e-32, 1.338126e-32, 1.338126e-32, 
    1.338126e-32, 1.338125e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 
    1.338122e-32, 1.338123e-32, 1.338123e-32, 1.338122e-32, 1.338123e-32, 
    1.33812e-32, 1.338122e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338118e-32, 1.338118e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338121e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338122e-32, 1.338121e-32, 1.338124e-32, 
    1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338121e-32, 1.338123e-32, 
    1.33812e-32, 1.338121e-32, 1.338118e-32, 1.338119e-32, 1.338117e-32, 
    1.338115e-32, 1.338114e-32, 1.338113e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338124e-32, 1.338121e-32, 1.338125e-32, 1.338124e-32, 1.338123e-32, 
    1.338123e-32, 1.338122e-32, 1.338121e-32, 1.33812e-32, 1.338121e-32, 
    1.338115e-32, 1.338118e-32, 1.338112e-32, 1.338113e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338121e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 
    1.338119e-32, 1.338121e-32, 1.33812e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338123e-32, 1.338122e-32, 1.33812e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338121e-32, 1.338115e-32, 1.338119e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 1.33812e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338118e-32, 1.338119e-32, 
    1.338119e-32, 1.33812e-32, 1.33812e-32, 1.338121e-32, 1.338122e-32, 
    1.338123e-32, 1.338123e-32, 1.338122e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338118e-32, 1.338121e-32, 1.33812e-32, 1.33812e-32, 
    1.338119e-32, 1.338122e-32, 1.338119e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338119e-32, 1.338119e-32, 
    1.33812e-32, 1.33812e-32, 1.338121e-32, 1.338121e-32, 1.338122e-32, 
    1.338123e-32, 1.338122e-32, 1.338122e-32, 1.33812e-32, 1.338119e-32, 
    1.338118e-32, 1.338118e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 
    1.338117e-32, 1.338114e-32, 1.338119e-32, 1.338117e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338119e-32, 1.338118e-32, 
    1.33812e-32, 1.338122e-32, 1.338122e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338122e-32, 1.338122e-32, 1.33812e-32, 1.338121e-32, 
    1.338119e-32, 1.338118e-32, 1.338115e-32, 1.338114e-32, 1.338113e-32, 
    1.338112e-32, 1.338112e-32, 1.338112e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.660867e-15, 1.665373e-15, 1.664498e-15, 1.668128e-15, 1.666115e-15, 
    1.668491e-15, 1.661782e-15, 1.665551e-15, 1.663145e-15, 1.661274e-15, 
    1.675163e-15, 1.66829e-15, 1.682295e-15, 1.67792e-15, 1.688904e-15, 
    1.681614e-15, 1.690373e-15, 1.688695e-15, 1.693745e-15, 1.692299e-15, 
    1.698748e-15, 1.694412e-15, 1.702089e-15, 1.697714e-15, 1.698398e-15, 
    1.694269e-15, 1.669675e-15, 1.674307e-15, 1.6694e-15, 1.670061e-15, 
    1.669765e-15, 1.666156e-15, 1.664335e-15, 1.660524e-15, 1.661216e-15, 
    1.664016e-15, 1.670358e-15, 1.668207e-15, 1.673629e-15, 1.673507e-15, 
    1.679534e-15, 1.676817e-15, 1.686935e-15, 1.684062e-15, 1.692359e-15, 
    1.690274e-15, 1.692261e-15, 1.691659e-15, 1.692269e-15, 1.689211e-15, 
    1.690521e-15, 1.687829e-15, 1.677326e-15, 1.680415e-15, 1.671194e-15, 
    1.665638e-15, 1.661947e-15, 1.659325e-15, 1.659696e-15, 1.660402e-15, 
    1.664032e-15, 1.667444e-15, 1.670042e-15, 1.671779e-15, 1.673489e-15, 
    1.678659e-15, 1.681396e-15, 1.687515e-15, 1.686413e-15, 1.688281e-15, 
    1.690067e-15, 1.693062e-15, 1.692569e-15, 1.693888e-15, 1.688233e-15, 
    1.691991e-15, 1.685784e-15, 1.687483e-15, 1.673949e-15, 1.668788e-15, 
    1.666588e-15, 1.664666e-15, 1.659981e-15, 1.663216e-15, 1.661941e-15, 
    1.664975e-15, 1.666902e-15, 1.665949e-15, 1.671826e-15, 1.669542e-15, 
    1.681558e-15, 1.676387e-15, 1.689858e-15, 1.686639e-15, 1.69063e-15, 
    1.688594e-15, 1.692081e-15, 1.688943e-15, 1.694379e-15, 1.695561e-15, 
    1.694753e-15, 1.697857e-15, 1.688769e-15, 1.692261e-15, 1.665922e-15, 
    1.666078e-15, 1.666802e-15, 1.663618e-15, 1.663423e-15, 1.660505e-15, 
    1.663102e-15, 1.664207e-15, 1.667014e-15, 1.668672e-15, 1.670248e-15, 
    1.673711e-15, 1.677575e-15, 1.682973e-15, 1.686848e-15, 1.689443e-15, 
    1.687852e-15, 1.689256e-15, 1.687686e-15, 1.68695e-15, 1.695117e-15, 
    1.690533e-15, 1.69741e-15, 1.69703e-15, 1.693919e-15, 1.697073e-15, 
    1.666187e-15, 1.665293e-15, 1.662186e-15, 1.664618e-15, 1.660187e-15, 
    1.662667e-15, 1.664092e-15, 1.669589e-15, 1.670797e-15, 1.671915e-15, 
    1.674124e-15, 1.676956e-15, 1.68192e-15, 1.686235e-15, 1.690171e-15, 
    1.689883e-15, 1.689984e-15, 1.690862e-15, 1.688686e-15, 1.69122e-15, 
    1.691644e-15, 1.690533e-15, 1.696979e-15, 1.695139e-15, 1.697022e-15, 
    1.695824e-15, 1.665584e-15, 1.667088e-15, 1.666275e-15, 1.667803e-15, 
    1.666726e-15, 1.671512e-15, 1.672946e-15, 1.679649e-15, 1.6769e-15, 
    1.681275e-15, 1.677345e-15, 1.678042e-15, 1.681416e-15, 1.677558e-15, 
    1.685997e-15, 1.680276e-15, 1.690896e-15, 1.685189e-15, 1.691254e-15, 
    1.690154e-15, 1.691975e-15, 1.693605e-15, 1.695656e-15, 1.699436e-15, 
    1.698561e-15, 1.701721e-15, 1.66933e-15, 1.671279e-15, 1.671108e-15, 
    1.673148e-15, 1.674655e-15, 1.677922e-15, 1.683154e-15, 1.681188e-15, 
    1.684799e-15, 1.685523e-15, 1.680037e-15, 1.683405e-15, 1.672584e-15, 
    1.674333e-15, 1.673292e-15, 1.669483e-15, 1.68164e-15, 1.675405e-15, 
    1.686912e-15, 1.68354e-15, 1.693373e-15, 1.688485e-15, 1.698079e-15, 
    1.702171e-15, 1.706023e-15, 1.710514e-15, 1.672343e-15, 1.671019e-15, 
    1.673391e-15, 1.676667e-15, 1.679708e-15, 1.683745e-15, 1.684159e-15, 
    1.684914e-15, 1.686872e-15, 1.688517e-15, 1.685152e-15, 1.688929e-15, 
    1.674737e-15, 1.682181e-15, 1.670518e-15, 1.674032e-15, 1.676475e-15, 
    1.675404e-15, 1.680963e-15, 1.682272e-15, 1.687586e-15, 1.68484e-15, 
    1.701161e-15, 1.693948e-15, 1.713933e-15, 1.708358e-15, 1.670556e-15, 
    1.672339e-15, 1.678537e-15, 1.675589e-15, 1.684015e-15, 1.686086e-15, 
    1.68777e-15, 1.689919e-15, 1.690152e-15, 1.691425e-15, 1.689338e-15, 
    1.691343e-15, 1.683754e-15, 1.687147e-15, 1.67783e-15, 1.680099e-15, 
    1.679055e-15, 1.67791e-15, 1.681444e-15, 1.685205e-15, 1.685287e-15, 
    1.686492e-15, 1.689882e-15, 1.684049e-15, 1.702088e-15, 1.690955e-15, 
    1.674282e-15, 1.67771e-15, 1.678202e-15, 1.676874e-15, 1.685878e-15, 
    1.682618e-15, 1.691394e-15, 1.689024e-15, 1.692907e-15, 1.690978e-15, 
    1.690694e-15, 1.688215e-15, 1.686671e-15, 1.682767e-15, 1.679588e-15, 
    1.677067e-15, 1.677653e-15, 1.680423e-15, 1.685435e-15, 1.690172e-15, 
    1.689135e-15, 1.692612e-15, 1.683405e-15, 1.687267e-15, 1.685774e-15, 
    1.689666e-15, 1.681135e-15, 1.688397e-15, 1.679276e-15, 1.680077e-15, 
    1.682553e-15, 1.687528e-15, 1.68863e-15, 1.689804e-15, 1.68908e-15, 
    1.685563e-15, 1.684987e-15, 1.682493e-15, 1.681804e-15, 1.679903e-15, 
    1.678328e-15, 1.679767e-15, 1.681277e-15, 1.685565e-15, 1.689424e-15, 
    1.693628e-15, 1.694657e-15, 1.699559e-15, 1.695567e-15, 1.70215e-15, 
    1.696551e-15, 1.70624e-15, 1.688819e-15, 1.696389e-15, 1.682666e-15, 
    1.684147e-15, 1.686823e-15, 1.692957e-15, 1.689648e-15, 1.693518e-15, 
    1.684964e-15, 1.680518e-15, 1.679368e-15, 1.67722e-15, 1.679417e-15, 
    1.679239e-15, 1.68134e-15, 1.680665e-15, 1.685707e-15, 1.683e-15, 
    1.690687e-15, 1.693488e-15, 1.701389e-15, 1.706224e-15, 1.711142e-15, 
    1.71331e-15, 1.71397e-15, 1.714246e-15 ;

 LITR3N_vr =
  7.663728e-06, 7.663721e-06, 7.663722e-06, 7.663716e-06, 7.663719e-06, 
    7.663715e-06, 7.663727e-06, 7.663721e-06, 7.663724e-06, 7.663728e-06, 
    7.663703e-06, 7.663715e-06, 7.663691e-06, 7.663699e-06, 7.66368e-06, 
    7.663692e-06, 7.663677e-06, 7.66368e-06, 7.663671e-06, 7.663673e-06, 
    7.663662e-06, 7.66367e-06, 7.663656e-06, 7.663664e-06, 7.663662e-06, 
    7.66367e-06, 7.663713e-06, 7.663705e-06, 7.663713e-06, 7.663712e-06, 
    7.663712e-06, 7.663719e-06, 7.663722e-06, 7.663729e-06, 7.663728e-06, 
    7.663722e-06, 7.663712e-06, 7.663715e-06, 7.663706e-06, 7.663706e-06, 
    7.663696e-06, 7.663701e-06, 7.663682e-06, 7.663688e-06, 7.663673e-06, 
    7.663677e-06, 7.663673e-06, 7.663674e-06, 7.663673e-06, 7.663679e-06, 
    7.663677e-06, 7.663682e-06, 7.6637e-06, 7.663694e-06, 7.663711e-06, 
    7.66372e-06, 7.663726e-06, 7.663731e-06, 7.663731e-06, 7.663729e-06, 
    7.663722e-06, 7.663717e-06, 7.663712e-06, 7.66371e-06, 7.663706e-06, 
    7.663697e-06, 7.663692e-06, 7.663682e-06, 7.663683e-06, 7.663681e-06, 
    7.663677e-06, 7.663672e-06, 7.663673e-06, 7.663671e-06, 7.663681e-06, 
    7.663674e-06, 7.663685e-06, 7.663682e-06, 7.663705e-06, 7.663714e-06, 
    7.663719e-06, 7.663722e-06, 7.66373e-06, 7.663724e-06, 7.663726e-06, 
    7.663722e-06, 7.663718e-06, 7.66372e-06, 7.663709e-06, 7.663713e-06, 
    7.663692e-06, 7.663702e-06, 7.663678e-06, 7.663683e-06, 7.663676e-06, 
    7.66368e-06, 7.663674e-06, 7.66368e-06, 7.66367e-06, 7.663668e-06, 
    7.663669e-06, 7.663663e-06, 7.66368e-06, 7.663673e-06, 7.66372e-06, 
    7.663719e-06, 7.663718e-06, 7.663723e-06, 7.663724e-06, 7.663729e-06, 
    7.663724e-06, 7.663722e-06, 7.663718e-06, 7.663715e-06, 7.663712e-06, 
    7.663706e-06, 7.663699e-06, 7.66369e-06, 7.663683e-06, 7.663679e-06, 
    7.663682e-06, 7.663679e-06, 7.663682e-06, 7.663682e-06, 7.663669e-06, 
    7.663677e-06, 7.663664e-06, 7.663665e-06, 7.663671e-06, 7.663665e-06, 
    7.663719e-06, 7.663721e-06, 7.663726e-06, 7.663722e-06, 7.66373e-06, 
    7.663725e-06, 7.663722e-06, 7.663713e-06, 7.663711e-06, 7.663709e-06, 
    7.663705e-06, 7.663701e-06, 7.663692e-06, 7.663684e-06, 7.663677e-06, 
    7.663678e-06, 7.663678e-06, 7.663676e-06, 7.66368e-06, 7.663675e-06, 
    7.663674e-06, 7.663677e-06, 7.663665e-06, 7.663669e-06, 7.663665e-06, 
    7.663667e-06, 7.66372e-06, 7.663718e-06, 7.663719e-06, 7.663716e-06, 
    7.663718e-06, 7.66371e-06, 7.663707e-06, 7.663695e-06, 7.663701e-06, 
    7.663692e-06, 7.6637e-06, 7.663699e-06, 7.663692e-06, 7.663699e-06, 
    7.663684e-06, 7.663694e-06, 7.663676e-06, 7.663686e-06, 7.663675e-06, 
    7.663677e-06, 7.663674e-06, 7.663672e-06, 7.663668e-06, 7.663661e-06, 
    7.663662e-06, 7.663657e-06, 7.663713e-06, 7.663711e-06, 7.663711e-06, 
    7.663707e-06, 7.663704e-06, 7.663699e-06, 7.66369e-06, 7.663692e-06, 
    7.663687e-06, 7.663685e-06, 7.663695e-06, 7.663689e-06, 7.663708e-06, 
    7.663705e-06, 7.663707e-06, 7.663713e-06, 7.663692e-06, 7.663703e-06, 
    7.663682e-06, 7.663689e-06, 7.663672e-06, 7.66368e-06, 7.663663e-06, 
    7.663656e-06, 7.66365e-06, 7.663642e-06, 7.663708e-06, 7.663711e-06, 
    7.663706e-06, 7.663701e-06, 7.663695e-06, 7.663689e-06, 7.663688e-06, 
    7.663686e-06, 7.663683e-06, 7.66368e-06, 7.663686e-06, 7.66368e-06, 
    7.663704e-06, 7.663692e-06, 7.663712e-06, 7.663705e-06, 7.663702e-06, 
    7.663703e-06, 7.663693e-06, 7.663691e-06, 7.663682e-06, 7.663686e-06, 
    7.663658e-06, 7.663671e-06, 7.663636e-06, 7.663645e-06, 7.663712e-06, 
    7.663708e-06, 7.663698e-06, 7.663702e-06, 7.663688e-06, 7.663684e-06, 
    7.663682e-06, 7.663678e-06, 7.663677e-06, 7.663675e-06, 7.663679e-06, 
    7.663675e-06, 7.663689e-06, 7.663682e-06, 7.663699e-06, 7.663695e-06, 
    7.663697e-06, 7.663699e-06, 7.663692e-06, 7.663686e-06, 7.663686e-06, 
    7.663683e-06, 7.663678e-06, 7.663688e-06, 7.663656e-06, 7.663676e-06, 
    7.663705e-06, 7.663699e-06, 7.663698e-06, 7.663701e-06, 7.663684e-06, 
    7.663691e-06, 7.663675e-06, 7.663679e-06, 7.663672e-06, 7.663676e-06, 
    7.663676e-06, 7.663681e-06, 7.663683e-06, 7.66369e-06, 7.663696e-06, 
    7.6637e-06, 7.663699e-06, 7.663694e-06, 7.663685e-06, 7.663677e-06, 
    7.663679e-06, 7.663673e-06, 7.663689e-06, 7.663682e-06, 7.663685e-06, 
    7.663678e-06, 7.663693e-06, 7.663681e-06, 7.663696e-06, 7.663695e-06, 
    7.663691e-06, 7.663682e-06, 7.66368e-06, 7.663678e-06, 7.663679e-06, 
    7.663685e-06, 7.663686e-06, 7.663691e-06, 7.663692e-06, 7.663695e-06, 
    7.663698e-06, 7.663695e-06, 7.663692e-06, 7.663685e-06, 7.663679e-06, 
    7.663672e-06, 7.66367e-06, 7.663661e-06, 7.663668e-06, 7.663656e-06, 
    7.663666e-06, 7.663649e-06, 7.66368e-06, 7.663666e-06, 7.663691e-06, 
    7.663688e-06, 7.663683e-06, 7.663672e-06, 7.663678e-06, 7.663672e-06, 
    7.663686e-06, 7.663694e-06, 7.663696e-06, 7.6637e-06, 7.663696e-06, 
    7.663696e-06, 7.663692e-06, 7.663693e-06, 7.663685e-06, 7.66369e-06, 
    7.663676e-06, 7.663672e-06, 7.663658e-06, 7.663649e-06, 7.663641e-06, 
    7.663637e-06, 7.663636e-06, 7.663635e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  6.000561e-14, 6.016838e-14, 6.013676e-14, 6.026792e-14, 6.01952e-14, 
    6.028104e-14, 6.003864e-14, 6.017481e-14, 6.008791e-14, 6.00203e-14, 
    6.052208e-14, 6.027377e-14, 6.077978e-14, 6.06217e-14, 6.101855e-14, 
    6.075516e-14, 6.10716e-14, 6.1011e-14, 6.119344e-14, 6.11412e-14, 
    6.13742e-14, 6.121755e-14, 6.14949e-14, 6.133683e-14, 6.136155e-14, 
    6.121237e-14, 6.032382e-14, 6.049118e-14, 6.031389e-14, 6.033777e-14, 
    6.032706e-14, 6.019668e-14, 6.01309e-14, 5.99932e-14, 6.001821e-14, 
    6.011937e-14, 6.034851e-14, 6.027079e-14, 6.046667e-14, 6.046226e-14, 
    6.068e-14, 6.058186e-14, 6.094741e-14, 6.084362e-14, 6.114339e-14, 
    6.106805e-14, 6.113984e-14, 6.111808e-14, 6.114013e-14, 6.102962e-14, 
    6.107697e-14, 6.097971e-14, 6.060023e-14, 6.071185e-14, 6.03787e-14, 
    6.017796e-14, 6.004461e-14, 5.994987e-14, 5.996327e-14, 5.99888e-14, 
    6.011996e-14, 6.024322e-14, 6.033707e-14, 6.039982e-14, 6.046162e-14, 
    6.064841e-14, 6.074729e-14, 6.096836e-14, 6.092854e-14, 6.099604e-14, 
    6.106055e-14, 6.116875e-14, 6.115095e-14, 6.119859e-14, 6.099429e-14, 
    6.113009e-14, 6.090583e-14, 6.09672e-14, 6.047825e-14, 6.029177e-14, 
    6.02123e-14, 6.014283e-14, 5.997357e-14, 6.009047e-14, 6.004439e-14, 
    6.015402e-14, 6.022362e-14, 6.018921e-14, 6.040153e-14, 6.031901e-14, 
    6.075314e-14, 6.05663e-14, 6.105303e-14, 6.093672e-14, 6.10809e-14, 
    6.100735e-14, 6.113334e-14, 6.101996e-14, 6.121633e-14, 6.125904e-14, 
    6.122986e-14, 6.134199e-14, 6.101367e-14, 6.113982e-14, 6.018824e-14, 
    6.019385e-14, 6.022001e-14, 6.010498e-14, 6.009795e-14, 5.99925e-14, 
    6.008635e-14, 6.012627e-14, 6.022767e-14, 6.028758e-14, 6.034452e-14, 
    6.046965e-14, 6.060924e-14, 6.080427e-14, 6.094425e-14, 6.1038e-14, 
    6.098054e-14, 6.103127e-14, 6.097455e-14, 6.094796e-14, 6.124303e-14, 
    6.10774e-14, 6.132587e-14, 6.131214e-14, 6.119972e-14, 6.131369e-14, 
    6.019779e-14, 6.016549e-14, 6.005324e-14, 6.014109e-14, 5.998102e-14, 
    6.007062e-14, 6.012211e-14, 6.03207e-14, 6.036434e-14, 6.040475e-14, 
    6.048455e-14, 6.058688e-14, 6.076623e-14, 6.092212e-14, 6.106431e-14, 
    6.10539e-14, 6.105756e-14, 6.10893e-14, 6.101067e-14, 6.110221e-14, 
    6.111755e-14, 6.10774e-14, 6.13103e-14, 6.12438e-14, 6.131184e-14, 
    6.126856e-14, 6.0176e-14, 6.023034e-14, 6.020098e-14, 6.025619e-14, 
    6.021728e-14, 6.039018e-14, 6.044198e-14, 6.068416e-14, 6.058486e-14, 
    6.074292e-14, 6.060094e-14, 6.06261e-14, 6.074801e-14, 6.060862e-14, 
    6.09135e-14, 6.070681e-14, 6.109053e-14, 6.088431e-14, 6.110344e-14, 
    6.10637e-14, 6.112951e-14, 6.11884e-14, 6.126249e-14, 6.139905e-14, 
    6.136744e-14, 6.14816e-14, 6.031135e-14, 6.038177e-14, 6.03756e-14, 
    6.044929e-14, 6.050375e-14, 6.062176e-14, 6.081082e-14, 6.073976e-14, 
    6.087021e-14, 6.089638e-14, 6.06982e-14, 6.081988e-14, 6.04289e-14, 
    6.049211e-14, 6.04545e-14, 6.031689e-14, 6.075609e-14, 6.053084e-14, 
    6.094656e-14, 6.082474e-14, 6.118e-14, 6.10034e-14, 6.135003e-14, 
    6.149789e-14, 6.163704e-14, 6.17993e-14, 6.042022e-14, 6.037239e-14, 
    6.045805e-14, 6.057644e-14, 6.068629e-14, 6.083216e-14, 6.08471e-14, 
    6.087439e-14, 6.094512e-14, 6.100455e-14, 6.088299e-14, 6.101944e-14, 
    6.05067e-14, 6.077565e-14, 6.035427e-14, 6.048124e-14, 6.056948e-14, 
    6.053081e-14, 6.073165e-14, 6.077894e-14, 6.097092e-14, 6.087172e-14, 
    6.146138e-14, 6.120079e-14, 6.192283e-14, 6.172141e-14, 6.035566e-14, 
    6.042007e-14, 6.064398e-14, 6.053749e-14, 6.084191e-14, 6.091673e-14, 
    6.097756e-14, 6.105523e-14, 6.106363e-14, 6.110963e-14, 6.103424e-14, 
    6.110666e-14, 6.083248e-14, 6.095507e-14, 6.061844e-14, 6.070042e-14, 
    6.066272e-14, 6.062133e-14, 6.074903e-14, 6.08849e-14, 6.088785e-14, 
    6.093138e-14, 6.105389e-14, 6.084315e-14, 6.149488e-14, 6.109265e-14, 
    6.049028e-14, 6.061413e-14, 6.063187e-14, 6.05839e-14, 6.090923e-14, 
    6.079143e-14, 6.110851e-14, 6.10229e-14, 6.116316e-14, 6.109347e-14, 
    6.108321e-14, 6.099366e-14, 6.093787e-14, 6.079683e-14, 6.068198e-14, 
    6.059087e-14, 6.061206e-14, 6.071212e-14, 6.089322e-14, 6.106437e-14, 
    6.102689e-14, 6.115251e-14, 6.081986e-14, 6.095941e-14, 6.090548e-14, 
    6.104608e-14, 6.073786e-14, 6.100022e-14, 6.067071e-14, 6.069964e-14, 
    6.078909e-14, 6.096884e-14, 6.100865e-14, 6.105106e-14, 6.10249e-14, 
    6.089783e-14, 6.087702e-14, 6.078693e-14, 6.076202e-14, 6.069335e-14, 
    6.063644e-14, 6.068842e-14, 6.074298e-14, 6.08979e-14, 6.103734e-14, 
    6.118923e-14, 6.12264e-14, 6.140349e-14, 6.125928e-14, 6.149711e-14, 
    6.129483e-14, 6.164486e-14, 6.101548e-14, 6.128898e-14, 6.079318e-14, 
    6.084669e-14, 6.094336e-14, 6.116496e-14, 6.104542e-14, 6.118524e-14, 
    6.08762e-14, 6.071555e-14, 6.067402e-14, 6.05964e-14, 6.06758e-14, 
    6.066934e-14, 6.074527e-14, 6.072088e-14, 6.090304e-14, 6.080522e-14, 
    6.108295e-14, 6.118414e-14, 6.146962e-14, 6.164431e-14, 6.182198e-14, 
    6.190031e-14, 6.192415e-14, 6.193412e-14 ;

 LITTERC =
  5.976235e-05, 5.97622e-05, 5.976223e-05, 5.976211e-05, 5.976218e-05, 
    5.97621e-05, 5.976232e-05, 5.97622e-05, 5.976228e-05, 5.976234e-05, 
    5.976188e-05, 5.976211e-05, 5.976165e-05, 5.976179e-05, 5.976143e-05, 
    5.976167e-05, 5.976138e-05, 5.976143e-05, 5.976127e-05, 5.976131e-05, 
    5.97611e-05, 5.976125e-05, 5.976099e-05, 5.976114e-05, 5.976111e-05, 
    5.976125e-05, 5.976206e-05, 5.976191e-05, 5.976207e-05, 5.976205e-05, 
    5.976206e-05, 5.976218e-05, 5.976224e-05, 5.976236e-05, 5.976234e-05, 
    5.976225e-05, 5.976204e-05, 5.976211e-05, 5.976193e-05, 5.976194e-05, 
    5.976174e-05, 5.976183e-05, 5.976149e-05, 5.976159e-05, 5.976131e-05, 
    5.976138e-05, 5.976131e-05, 5.976134e-05, 5.976131e-05, 5.976142e-05, 
    5.976137e-05, 5.976146e-05, 5.976181e-05, 5.976171e-05, 5.976201e-05, 
    5.976219e-05, 5.976231e-05, 5.97624e-05, 5.976239e-05, 5.976237e-05, 
    5.976225e-05, 5.976214e-05, 5.976205e-05, 5.976199e-05, 5.976194e-05, 
    5.976177e-05, 5.976167e-05, 5.976147e-05, 5.976151e-05, 5.976145e-05, 
    5.976139e-05, 5.976129e-05, 5.976131e-05, 5.976126e-05, 5.976145e-05, 
    5.976133e-05, 5.976153e-05, 5.976147e-05, 5.976192e-05, 5.976209e-05, 
    5.976216e-05, 5.976223e-05, 5.976238e-05, 5.976227e-05, 5.976231e-05, 
    5.976222e-05, 5.976215e-05, 5.976218e-05, 5.976199e-05, 5.976207e-05, 
    5.976167e-05, 5.976184e-05, 5.976139e-05, 5.97615e-05, 5.976137e-05, 
    5.976144e-05, 5.976132e-05, 5.976143e-05, 5.976125e-05, 5.976121e-05, 
    5.976123e-05, 5.976113e-05, 5.976143e-05, 5.976131e-05, 5.976218e-05, 
    5.976218e-05, 5.976215e-05, 5.976226e-05, 5.976227e-05, 5.976237e-05, 
    5.976228e-05, 5.976224e-05, 5.976215e-05, 5.976209e-05, 5.976204e-05, 
    5.976193e-05, 5.97618e-05, 5.976162e-05, 5.97615e-05, 5.976141e-05, 
    5.976146e-05, 5.976142e-05, 5.976147e-05, 5.976149e-05, 5.976122e-05, 
    5.976137e-05, 5.976115e-05, 5.976116e-05, 5.976126e-05, 5.976116e-05, 
    5.976218e-05, 5.976221e-05, 5.976231e-05, 5.976223e-05, 5.976237e-05, 
    5.976229e-05, 5.976225e-05, 5.976206e-05, 5.976202e-05, 5.976199e-05, 
    5.976191e-05, 5.976182e-05, 5.976166e-05, 5.976151e-05, 5.976138e-05, 
    5.976139e-05, 5.976139e-05, 5.976136e-05, 5.976143e-05, 5.976135e-05, 
    5.976134e-05, 5.976137e-05, 5.976116e-05, 5.976122e-05, 5.976116e-05, 
    5.97612e-05, 5.976219e-05, 5.976215e-05, 5.976217e-05, 5.976212e-05, 
    5.976216e-05, 5.9762e-05, 5.976195e-05, 5.976173e-05, 5.976182e-05, 
    5.976168e-05, 5.976181e-05, 5.976178e-05, 5.976167e-05, 5.97618e-05, 
    5.976152e-05, 5.976171e-05, 5.976136e-05, 5.976155e-05, 5.976135e-05, 
    5.976139e-05, 5.976133e-05, 5.976127e-05, 5.976121e-05, 5.976108e-05, 
    5.976111e-05, 5.976101e-05, 5.976207e-05, 5.976201e-05, 5.976201e-05, 
    5.976195e-05, 5.97619e-05, 5.976179e-05, 5.976162e-05, 5.976168e-05, 
    5.976156e-05, 5.976154e-05, 5.976172e-05, 5.976161e-05, 5.976197e-05, 
    5.976191e-05, 5.976194e-05, 5.976207e-05, 5.976167e-05, 5.976187e-05, 
    5.976149e-05, 5.976161e-05, 5.976128e-05, 5.976144e-05, 5.976113e-05, 
    5.976099e-05, 5.976086e-05, 5.976071e-05, 5.976197e-05, 5.976202e-05, 
    5.976194e-05, 5.976183e-05, 5.976173e-05, 5.97616e-05, 5.976158e-05, 
    5.976156e-05, 5.976149e-05, 5.976144e-05, 5.976155e-05, 5.976143e-05, 
    5.976189e-05, 5.976165e-05, 5.976203e-05, 5.976192e-05, 5.976184e-05, 
    5.976187e-05, 5.976169e-05, 5.976165e-05, 5.976147e-05, 5.976156e-05, 
    5.976102e-05, 5.976126e-05, 5.97606e-05, 5.976078e-05, 5.976203e-05, 
    5.976197e-05, 5.976177e-05, 5.976187e-05, 5.976159e-05, 5.976152e-05, 
    5.976146e-05, 5.976139e-05, 5.976139e-05, 5.976134e-05, 5.976141e-05, 
    5.976135e-05, 5.97616e-05, 5.976149e-05, 5.976179e-05, 5.976172e-05, 
    5.976175e-05, 5.976179e-05, 5.976167e-05, 5.976155e-05, 5.976155e-05, 
    5.976151e-05, 5.976139e-05, 5.976159e-05, 5.976099e-05, 5.976136e-05, 
    5.976191e-05, 5.976179e-05, 5.976178e-05, 5.976182e-05, 5.976153e-05, 
    5.976163e-05, 5.976134e-05, 5.976142e-05, 5.97613e-05, 5.976136e-05, 
    5.976137e-05, 5.976145e-05, 5.97615e-05, 5.976163e-05, 5.976173e-05, 
    5.976182e-05, 5.97618e-05, 5.976171e-05, 5.976154e-05, 5.976138e-05, 
    5.976142e-05, 5.97613e-05, 5.976161e-05, 5.976148e-05, 5.976153e-05, 
    5.97614e-05, 5.976168e-05, 5.976145e-05, 5.976174e-05, 5.976172e-05, 
    5.976164e-05, 5.976147e-05, 5.976143e-05, 5.97614e-05, 5.976142e-05, 
    5.976154e-05, 5.976155e-05, 5.976164e-05, 5.976166e-05, 5.976173e-05, 
    5.976178e-05, 5.976173e-05, 5.976168e-05, 5.976154e-05, 5.976141e-05, 
    5.976127e-05, 5.976124e-05, 5.976107e-05, 5.976121e-05, 5.976099e-05, 
    5.976118e-05, 5.976086e-05, 5.976143e-05, 5.976118e-05, 5.976163e-05, 
    5.976158e-05, 5.97615e-05, 5.976129e-05, 5.97614e-05, 5.976127e-05, 
    5.976156e-05, 5.97617e-05, 5.976174e-05, 5.976181e-05, 5.976174e-05, 
    5.976175e-05, 5.976168e-05, 5.97617e-05, 5.976153e-05, 5.976162e-05, 
    5.976137e-05, 5.976127e-05, 5.976102e-05, 5.976086e-05, 5.976069e-05, 
    5.976062e-05, 5.97606e-05, 5.976059e-05 ;

 LITTERC_HR =
  9.681104e-13, 9.707342e-13, 9.702246e-13, 9.723389e-13, 9.711665e-13, 
    9.725504e-13, 9.686429e-13, 9.70838e-13, 9.694371e-13, 9.683471e-13, 
    9.764359e-13, 9.724333e-13, 9.805901e-13, 9.780419e-13, 9.84439e-13, 
    9.801932e-13, 9.852943e-13, 9.843174e-13, 9.872582e-13, 9.864161e-13, 
    9.901719e-13, 9.876468e-13, 9.921177e-13, 9.895696e-13, 9.899681e-13, 
    9.875633e-13, 9.7324e-13, 9.759378e-13, 9.730799e-13, 9.734648e-13, 
    9.732923e-13, 9.711905e-13, 9.701301e-13, 9.679102e-13, 9.683135e-13, 
    9.699442e-13, 9.736379e-13, 9.723851e-13, 9.755428e-13, 9.754715e-13, 
    9.789815e-13, 9.773996e-13, 9.832922e-13, 9.816191e-13, 9.864514e-13, 
    9.85237e-13, 9.863941e-13, 9.860434e-13, 9.863988e-13, 9.846174e-13, 
    9.853807e-13, 9.83813e-13, 9.776958e-13, 9.794949e-13, 9.741246e-13, 
    9.708887e-13, 9.687391e-13, 9.67212e-13, 9.674279e-13, 9.678393e-13, 
    9.699537e-13, 9.719406e-13, 9.734535e-13, 9.744651e-13, 9.754612e-13, 
    9.784723e-13, 9.800662e-13, 9.836301e-13, 9.82988e-13, 9.840761e-13, 
    9.851161e-13, 9.868602e-13, 9.865733e-13, 9.873413e-13, 9.840479e-13, 
    9.862369e-13, 9.82622e-13, 9.836112e-13, 9.757294e-13, 9.727233e-13, 
    9.714423e-13, 9.703225e-13, 9.675938e-13, 9.694783e-13, 9.687355e-13, 
    9.705029e-13, 9.716248e-13, 9.7107e-13, 9.744927e-13, 9.731625e-13, 
    9.801606e-13, 9.771488e-13, 9.849949e-13, 9.831198e-13, 9.854441e-13, 
    9.842585e-13, 9.862894e-13, 9.844618e-13, 9.876273e-13, 9.883157e-13, 
    9.878452e-13, 9.896528e-13, 9.843603e-13, 9.863939e-13, 9.710544e-13, 
    9.711448e-13, 9.715666e-13, 9.697122e-13, 9.695989e-13, 9.67899e-13, 
    9.694118e-13, 9.700555e-13, 9.7169e-13, 9.726558e-13, 9.735737e-13, 
    9.755907e-13, 9.77841e-13, 9.809848e-13, 9.832414e-13, 9.847526e-13, 
    9.838262e-13, 9.846441e-13, 9.837297e-13, 9.833011e-13, 9.880576e-13, 
    9.853878e-13, 9.893929e-13, 9.891715e-13, 9.873595e-13, 9.891965e-13, 
    9.712084e-13, 9.706877e-13, 9.688782e-13, 9.702944e-13, 9.677139e-13, 
    9.691583e-13, 9.699883e-13, 9.731897e-13, 9.738932e-13, 9.745446e-13, 
    9.75831e-13, 9.774806e-13, 9.803716e-13, 9.828846e-13, 9.851767e-13, 
    9.850088e-13, 9.850679e-13, 9.855795e-13, 9.843119e-13, 9.857875e-13, 
    9.860348e-13, 9.853878e-13, 9.891419e-13, 9.8807e-13, 9.891669e-13, 
    9.884691e-13, 9.708571e-13, 9.717332e-13, 9.712597e-13, 9.721498e-13, 
    9.715226e-13, 9.743097e-13, 9.751447e-13, 9.790488e-13, 9.774479e-13, 
    9.799959e-13, 9.777072e-13, 9.781127e-13, 9.800779e-13, 9.77831e-13, 
    9.827456e-13, 9.794138e-13, 9.855993e-13, 9.822751e-13, 9.858074e-13, 
    9.851668e-13, 9.862276e-13, 9.871769e-13, 9.883713e-13, 9.905725e-13, 
    9.900631e-13, 9.919032e-13, 9.73039e-13, 9.741741e-13, 9.740747e-13, 
    9.752625e-13, 9.761404e-13, 9.780428e-13, 9.810904e-13, 9.79945e-13, 
    9.820479e-13, 9.824696e-13, 9.792749e-13, 9.812365e-13, 9.74934e-13, 
    9.759528e-13, 9.753466e-13, 9.731283e-13, 9.802082e-13, 9.765771e-13, 
    9.832786e-13, 9.813147e-13, 9.870416e-13, 9.841947e-13, 9.897825e-13, 
    9.921658e-13, 9.944088e-13, 9.970244e-13, 9.74794e-13, 9.740228e-13, 
    9.754039e-13, 9.773123e-13, 9.79083e-13, 9.814344e-13, 9.816752e-13, 
    9.821152e-13, 9.832554e-13, 9.842133e-13, 9.822539e-13, 9.844534e-13, 
    9.761881e-13, 9.805235e-13, 9.737309e-13, 9.757776e-13, 9.772001e-13, 
    9.765767e-13, 9.798141e-13, 9.805764e-13, 9.836712e-13, 9.820722e-13, 
    9.915773e-13, 9.873767e-13, 9.990156e-13, 9.957689e-13, 9.737533e-13, 
    9.747916e-13, 9.78401e-13, 9.766843e-13, 9.815917e-13, 9.827977e-13, 
    9.837783e-13, 9.850302e-13, 9.851656e-13, 9.859071e-13, 9.846919e-13, 
    9.858593e-13, 9.814395e-13, 9.834157e-13, 9.779893e-13, 9.793108e-13, 
    9.787031e-13, 9.78036e-13, 9.800944e-13, 9.822847e-13, 9.823322e-13, 
    9.830339e-13, 9.850087e-13, 9.816115e-13, 9.921174e-13, 9.856334e-13, 
    9.759232e-13, 9.779198e-13, 9.782058e-13, 9.774325e-13, 9.826768e-13, 
    9.807779e-13, 9.858892e-13, 9.84509e-13, 9.867701e-13, 9.856468e-13, 
    9.854814e-13, 9.840378e-13, 9.831385e-13, 9.808648e-13, 9.790134e-13, 
    9.775448e-13, 9.778864e-13, 9.794995e-13, 9.824187e-13, 9.851775e-13, 
    9.845734e-13, 9.865984e-13, 9.812361e-13, 9.834858e-13, 9.826162e-13, 
    9.848829e-13, 9.799144e-13, 9.841435e-13, 9.788318e-13, 9.792982e-13, 
    9.807402e-13, 9.836377e-13, 9.842794e-13, 9.84963e-13, 9.845413e-13, 
    9.824929e-13, 9.821575e-13, 9.807053e-13, 9.803037e-13, 9.791968e-13, 
    9.782794e-13, 9.791173e-13, 9.799968e-13, 9.824941e-13, 9.847419e-13, 
    9.871904e-13, 9.877895e-13, 9.906442e-13, 9.883195e-13, 9.921533e-13, 
    9.888926e-13, 9.94535e-13, 9.843895e-13, 9.887982e-13, 9.80806e-13, 
    9.816685e-13, 9.83227e-13, 9.867991e-13, 9.848722e-13, 9.87126e-13, 
    9.821445e-13, 9.795547e-13, 9.788852e-13, 9.77634e-13, 9.789138e-13, 
    9.788098e-13, 9.800338e-13, 9.796405e-13, 9.82577e-13, 9.810002e-13, 
    9.85477e-13, 9.871084e-13, 9.917101e-13, 9.94526e-13, 9.9739e-13, 
    9.986528e-13, 9.99037e-13, 9.991976e-13 ;

 LITTERC_LOSS =
  1.792931e-12, 1.79779e-12, 1.796847e-12, 1.800762e-12, 1.798591e-12, 
    1.801154e-12, 1.793917e-12, 1.797983e-12, 1.795388e-12, 1.79337e-12, 
    1.80835e-12, 1.800937e-12, 1.816044e-12, 1.811324e-12, 1.823172e-12, 
    1.815309e-12, 1.824756e-12, 1.822947e-12, 1.828393e-12, 1.826834e-12, 
    1.833789e-12, 1.829113e-12, 1.837393e-12, 1.832674e-12, 1.833412e-12, 
    1.828958e-12, 1.802431e-12, 1.807427e-12, 1.802135e-12, 1.802848e-12, 
    1.802528e-12, 1.798635e-12, 1.796672e-12, 1.79256e-12, 1.793307e-12, 
    1.796327e-12, 1.803168e-12, 1.800848e-12, 1.806696e-12, 1.806564e-12, 
    1.813065e-12, 1.810135e-12, 1.821048e-12, 1.81795e-12, 1.826899e-12, 
    1.82465e-12, 1.826793e-12, 1.826143e-12, 1.826802e-12, 1.823503e-12, 
    1.824916e-12, 1.822013e-12, 1.810683e-12, 1.814015e-12, 1.804069e-12, 
    1.798077e-12, 1.794095e-12, 1.791267e-12, 1.791667e-12, 1.792429e-12, 
    1.796345e-12, 1.800025e-12, 1.802827e-12, 1.8047e-12, 1.806545e-12, 
    1.812122e-12, 1.815073e-12, 1.821674e-12, 1.820485e-12, 1.8225e-12, 
    1.824426e-12, 1.827656e-12, 1.827125e-12, 1.828547e-12, 1.822448e-12, 
    1.826502e-12, 1.819807e-12, 1.821639e-12, 1.807042e-12, 1.801474e-12, 
    1.799102e-12, 1.797028e-12, 1.791974e-12, 1.795464e-12, 1.794089e-12, 
    1.797362e-12, 1.79944e-12, 1.798412e-12, 1.804751e-12, 1.802288e-12, 
    1.815248e-12, 1.80967e-12, 1.824201e-12, 1.820729e-12, 1.825033e-12, 
    1.822838e-12, 1.826599e-12, 1.823214e-12, 1.829077e-12, 1.830352e-12, 
    1.82948e-12, 1.832828e-12, 1.823026e-12, 1.826792e-12, 1.798383e-12, 
    1.798551e-12, 1.799332e-12, 1.795898e-12, 1.795688e-12, 1.79254e-12, 
    1.795341e-12, 1.796534e-12, 1.799561e-12, 1.801349e-12, 1.803049e-12, 
    1.806785e-12, 1.810952e-12, 1.816775e-12, 1.820954e-12, 1.823753e-12, 
    1.822037e-12, 1.823552e-12, 1.821858e-12, 1.821065e-12, 1.829873e-12, 
    1.824929e-12, 1.832347e-12, 1.831937e-12, 1.828581e-12, 1.831983e-12, 
    1.798669e-12, 1.797704e-12, 1.794353e-12, 1.796976e-12, 1.792197e-12, 
    1.794872e-12, 1.796409e-12, 1.802338e-12, 1.803641e-12, 1.804847e-12, 
    1.80723e-12, 1.810285e-12, 1.815639e-12, 1.820293e-12, 1.824538e-12, 
    1.824227e-12, 1.824337e-12, 1.825284e-12, 1.822937e-12, 1.825669e-12, 
    1.826127e-12, 1.824929e-12, 1.831882e-12, 1.829897e-12, 1.831928e-12, 
    1.830636e-12, 1.798018e-12, 1.799641e-12, 1.798764e-12, 1.800412e-12, 
    1.799251e-12, 1.804412e-12, 1.805959e-12, 1.813189e-12, 1.810224e-12, 
    1.814943e-12, 1.810704e-12, 1.811455e-12, 1.815095e-12, 1.810934e-12, 
    1.820036e-12, 1.813865e-12, 1.825321e-12, 1.819164e-12, 1.825706e-12, 
    1.82452e-12, 1.826484e-12, 1.828243e-12, 1.830455e-12, 1.834531e-12, 
    1.833588e-12, 1.836996e-12, 1.802059e-12, 1.804161e-12, 1.803977e-12, 
    1.806177e-12, 1.807803e-12, 1.811326e-12, 1.81697e-12, 1.814849e-12, 
    1.818744e-12, 1.819525e-12, 1.813608e-12, 1.817241e-12, 1.805568e-12, 
    1.807455e-12, 1.806333e-12, 1.802224e-12, 1.815337e-12, 1.808612e-12, 
    1.821023e-12, 1.817386e-12, 1.827992e-12, 1.822719e-12, 1.833068e-12, 
    1.837482e-12, 1.841636e-12, 1.84648e-12, 1.805309e-12, 1.803881e-12, 
    1.806439e-12, 1.809973e-12, 1.813253e-12, 1.817607e-12, 1.818053e-12, 
    1.818868e-12, 1.82098e-12, 1.822754e-12, 1.819125e-12, 1.823198e-12, 
    1.807891e-12, 1.81592e-12, 1.80334e-12, 1.807131e-12, 1.809765e-12, 
    1.808611e-12, 1.814607e-12, 1.816018e-12, 1.82175e-12, 1.818789e-12, 
    1.836392e-12, 1.828613e-12, 1.850168e-12, 1.844155e-12, 1.803382e-12, 
    1.805305e-12, 1.811989e-12, 1.80881e-12, 1.817899e-12, 1.820132e-12, 
    1.821948e-12, 1.824267e-12, 1.824518e-12, 1.825891e-12, 1.82364e-12, 
    1.825802e-12, 1.817617e-12, 1.821277e-12, 1.811227e-12, 1.813675e-12, 
    1.812549e-12, 1.811313e-12, 1.815126e-12, 1.819182e-12, 1.81927e-12, 
    1.82057e-12, 1.824227e-12, 1.817935e-12, 1.837392e-12, 1.825384e-12, 
    1.807401e-12, 1.811098e-12, 1.811628e-12, 1.810196e-12, 1.819908e-12, 
    1.816392e-12, 1.825858e-12, 1.823302e-12, 1.827489e-12, 1.825409e-12, 
    1.825103e-12, 1.822429e-12, 1.820763e-12, 1.816553e-12, 1.813124e-12, 
    1.810404e-12, 1.811036e-12, 1.814024e-12, 1.81943e-12, 1.82454e-12, 
    1.823421e-12, 1.827171e-12, 1.81724e-12, 1.821407e-12, 1.819796e-12, 
    1.823994e-12, 1.814792e-12, 1.822625e-12, 1.812787e-12, 1.813651e-12, 
    1.816322e-12, 1.821688e-12, 1.822876e-12, 1.824142e-12, 1.823362e-12, 
    1.819568e-12, 1.818947e-12, 1.816257e-12, 1.815513e-12, 1.813463e-12, 
    1.811764e-12, 1.813316e-12, 1.814945e-12, 1.81957e-12, 1.823733e-12, 
    1.828268e-12, 1.829377e-12, 1.834664e-12, 1.830359e-12, 1.837459e-12, 
    1.83142e-12, 1.84187e-12, 1.82308e-12, 1.831245e-12, 1.816444e-12, 
    1.818041e-12, 1.820927e-12, 1.827543e-12, 1.823974e-12, 1.828148e-12, 
    1.818922e-12, 1.814126e-12, 1.812886e-12, 1.810569e-12, 1.812939e-12, 
    1.812746e-12, 1.815013e-12, 1.814285e-12, 1.819723e-12, 1.816803e-12, 
    1.825094e-12, 1.828116e-12, 1.836638e-12, 1.841853e-12, 1.847157e-12, 
    1.849496e-12, 1.850208e-12, 1.850505e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.698539e-18, 1.698815e-18, 1.698762e-18, 1.698983e-18, 1.698862e-18, 
    1.699005e-18, 1.698597e-18, 1.698824e-18, 1.69868e-18, 1.698567e-18, 
    1.699405e-18, 1.698993e-18, 1.699856e-18, 1.699588e-18, 1.700267e-18, 
    1.699811e-18, 1.70036e-18, 1.700259e-18, 1.700576e-18, 1.700486e-18, 
    1.700882e-18, 1.700618e-18, 1.701096e-18, 1.700822e-18, 1.700863e-18, 
    1.700609e-18, 1.699081e-18, 1.699352e-18, 1.699063e-18, 1.699102e-18, 
    1.699086e-18, 1.698863e-18, 1.698748e-18, 1.698521e-18, 1.698563e-18, 
    1.698731e-18, 1.69912e-18, 1.698991e-18, 1.699326e-18, 1.699318e-18, 
    1.699689e-18, 1.699521e-18, 1.700149e-18, 1.699972e-18, 1.70049e-18, 
    1.700358e-18, 1.700483e-18, 1.700446e-18, 1.700483e-18, 1.700291e-18, 
    1.700373e-18, 1.700206e-18, 1.699552e-18, 1.699742e-18, 1.699173e-18, 
    1.698825e-18, 1.698606e-18, 1.698447e-18, 1.69847e-18, 1.698511e-18, 
    1.698732e-18, 1.698944e-18, 1.699105e-18, 1.699211e-18, 1.699317e-18, 
    1.699625e-18, 1.6998e-18, 1.700183e-18, 1.700118e-18, 1.700231e-18, 
    1.700346e-18, 1.700532e-18, 1.700502e-18, 1.700583e-18, 1.700231e-18, 
    1.700464e-18, 1.70008e-18, 1.700184e-18, 1.699329e-18, 1.699027e-18, 
    1.698884e-18, 1.698772e-18, 1.698487e-18, 1.698683e-18, 1.698605e-18, 
    1.698793e-18, 1.698911e-18, 1.698853e-18, 1.699214e-18, 1.699073e-18, 
    1.69981e-18, 1.699492e-18, 1.700332e-18, 1.700131e-18, 1.700381e-18, 
    1.700254e-18, 1.70047e-18, 1.700276e-18, 1.700615e-18, 1.700687e-18, 
    1.700637e-18, 1.700834e-18, 1.700265e-18, 1.700481e-18, 1.698851e-18, 
    1.69886e-18, 1.698905e-18, 1.698707e-18, 1.698696e-18, 1.698519e-18, 
    1.698678e-18, 1.698744e-18, 1.698919e-18, 1.699019e-18, 1.699116e-18, 
    1.699329e-18, 1.699565e-18, 1.6999e-18, 1.700144e-18, 1.700307e-18, 
    1.700208e-18, 1.700296e-18, 1.700197e-18, 1.700152e-18, 1.700659e-18, 
    1.700373e-18, 1.700806e-18, 1.700782e-18, 1.700585e-18, 1.700785e-18, 
    1.698867e-18, 1.698813e-18, 1.698621e-18, 1.698772e-18, 1.6985e-18, 
    1.69865e-18, 1.698735e-18, 1.699072e-18, 1.699151e-18, 1.699218e-18, 
    1.699356e-18, 1.69953e-18, 1.699835e-18, 1.700104e-18, 1.700353e-18, 
    1.700335e-18, 1.700341e-18, 1.700395e-18, 1.700259e-18, 1.700417e-18, 
    1.700442e-18, 1.700375e-18, 1.700779e-18, 1.700663e-18, 1.700782e-18, 
    1.700707e-18, 1.698831e-18, 1.698922e-18, 1.698873e-18, 1.698965e-18, 
    1.698899e-18, 1.69919e-18, 1.699277e-18, 1.699691e-18, 1.699526e-18, 
    1.699794e-18, 1.699554e-18, 1.699596e-18, 1.699796e-18, 1.699568e-18, 
    1.700086e-18, 1.699728e-18, 1.700397e-18, 1.700032e-18, 1.70042e-18, 
    1.700352e-18, 1.700466e-18, 1.700566e-18, 1.700696e-18, 1.70093e-18, 
    1.700876e-18, 1.701075e-18, 1.69906e-18, 1.699177e-18, 1.69917e-18, 
    1.699295e-18, 1.699387e-18, 1.69959e-18, 1.699913e-18, 1.699793e-18, 
    1.700018e-18, 1.700062e-18, 1.699722e-18, 1.699928e-18, 1.699259e-18, 
    1.699363e-18, 1.699303e-18, 1.699068e-18, 1.699816e-18, 1.69943e-18, 
    1.700148e-18, 1.699938e-18, 1.700551e-18, 1.700243e-18, 1.700846e-18, 
    1.701097e-18, 1.701348e-18, 1.701625e-18, 1.699245e-18, 1.699165e-18, 
    1.699311e-18, 1.699508e-18, 1.6997e-18, 1.69995e-18, 1.699978e-18, 
    1.700024e-18, 1.700147e-18, 1.700249e-18, 1.700035e-18, 1.700275e-18, 
    1.699381e-18, 1.699851e-18, 1.699132e-18, 1.699344e-18, 1.699498e-18, 
    1.699433e-18, 1.69978e-18, 1.699861e-18, 1.700188e-18, 1.70002e-18, 
    1.701032e-18, 1.700583e-18, 1.701847e-18, 1.70149e-18, 1.699136e-18, 
    1.699246e-18, 1.699625e-18, 1.699445e-18, 1.699969e-18, 1.700096e-18, 
    1.700203e-18, 1.700335e-18, 1.700351e-18, 1.700429e-18, 1.700301e-18, 
    1.700426e-18, 1.699951e-18, 1.700163e-18, 1.699586e-18, 1.699724e-18, 
    1.699661e-18, 1.69959e-18, 1.699809e-18, 1.700038e-18, 1.700048e-18, 
    1.70012e-18, 1.700315e-18, 1.699971e-18, 1.701081e-18, 1.700385e-18, 
    1.699366e-18, 1.699571e-18, 1.699607e-18, 1.699526e-18, 1.700084e-18, 
    1.699881e-18, 1.700428e-18, 1.700281e-18, 1.700524e-18, 1.700403e-18, 
    1.700385e-18, 1.700231e-18, 1.700133e-18, 1.699889e-18, 1.699692e-18, 
    1.699539e-18, 1.699575e-18, 1.699743e-18, 1.700053e-18, 1.70035e-18, 
    1.700284e-18, 1.700505e-18, 1.699931e-18, 1.700169e-18, 1.700075e-18, 
    1.70032e-18, 1.699788e-18, 1.700226e-18, 1.699675e-18, 1.699724e-18, 
    1.699877e-18, 1.700181e-18, 1.700256e-18, 1.700327e-18, 1.700285e-18, 
    1.700062e-18, 1.700028e-18, 1.699874e-18, 1.699829e-18, 1.699714e-18, 
    1.699616e-18, 1.699704e-18, 1.699796e-18, 1.700064e-18, 1.700303e-18, 
    1.700567e-18, 1.700633e-18, 1.700929e-18, 1.700681e-18, 1.701083e-18, 
    1.700731e-18, 1.701347e-18, 1.700259e-18, 1.700731e-18, 1.699885e-18, 
    1.699977e-18, 1.700138e-18, 1.70052e-18, 1.700319e-18, 1.700556e-18, 
    1.700027e-18, 1.699746e-18, 1.69968e-18, 1.699547e-18, 1.699683e-18, 
    1.699673e-18, 1.699803e-18, 1.699761e-18, 1.700073e-18, 1.699906e-18, 
    1.700383e-18, 1.700556e-18, 1.701053e-18, 1.701355e-18, 1.701672e-18, 
    1.70181e-18, 1.701852e-18, 1.70187e-18 ;

 MEG_acetic_acid =
  2.547808e-19, 2.548222e-19, 2.548143e-19, 2.548474e-19, 2.548293e-19, 
    2.548508e-19, 2.547895e-19, 2.548236e-19, 2.54802e-19, 2.54785e-19, 
    2.549108e-19, 2.548489e-19, 2.549783e-19, 2.549382e-19, 2.550401e-19, 
    2.549716e-19, 2.55054e-19, 2.550389e-19, 2.550864e-19, 2.550729e-19, 
    2.551323e-19, 2.550928e-19, 2.551644e-19, 2.551233e-19, 2.551294e-19, 
    2.550913e-19, 2.548621e-19, 2.549028e-19, 2.548595e-19, 2.548653e-19, 
    2.548629e-19, 2.548295e-19, 2.548121e-19, 2.547782e-19, 2.547844e-19, 
    2.548097e-19, 2.54868e-19, 2.548487e-19, 2.548989e-19, 2.548978e-19, 
    2.549533e-19, 2.549282e-19, 2.550224e-19, 2.549957e-19, 2.550734e-19, 
    2.550537e-19, 2.550724e-19, 2.550668e-19, 2.550724e-19, 2.550436e-19, 
    2.550559e-19, 2.550308e-19, 2.549327e-19, 2.549613e-19, 2.548759e-19, 
    2.548237e-19, 2.547909e-19, 2.547671e-19, 2.547705e-19, 2.547767e-19, 
    2.548098e-19, 2.548416e-19, 2.548657e-19, 2.548817e-19, 2.548976e-19, 
    2.549438e-19, 2.549699e-19, 2.550274e-19, 2.550176e-19, 2.550346e-19, 
    2.550518e-19, 2.550798e-19, 2.550753e-19, 2.550875e-19, 2.550347e-19, 
    2.550695e-19, 2.55012e-19, 2.550276e-19, 2.548994e-19, 2.54854e-19, 
    2.548326e-19, 2.548158e-19, 2.54773e-19, 2.548024e-19, 2.547907e-19, 
    2.54819e-19, 2.548366e-19, 2.54828e-19, 2.548822e-19, 2.54861e-19, 
    2.549715e-19, 2.549238e-19, 2.550498e-19, 2.550197e-19, 2.550571e-19, 
    2.550382e-19, 2.550705e-19, 2.550414e-19, 2.550922e-19, 2.55103e-19, 
    2.550956e-19, 2.551251e-19, 2.550397e-19, 2.550721e-19, 2.548276e-19, 
    2.54829e-19, 2.548358e-19, 2.54806e-19, 2.548043e-19, 2.547779e-19, 
    2.548016e-19, 2.548116e-19, 2.548378e-19, 2.548529e-19, 2.548674e-19, 
    2.548994e-19, 2.549347e-19, 2.54985e-19, 2.550216e-19, 2.550461e-19, 
    2.550313e-19, 2.550443e-19, 2.550296e-19, 2.550228e-19, 2.550988e-19, 
    2.550559e-19, 2.551208e-19, 2.551173e-19, 2.550877e-19, 2.551177e-19, 
    2.5483e-19, 2.54822e-19, 2.547932e-19, 2.548157e-19, 2.54775e-19, 
    2.547975e-19, 2.548102e-19, 2.548609e-19, 2.548726e-19, 2.548828e-19, 
    2.549033e-19, 2.549295e-19, 2.549753e-19, 2.550156e-19, 2.550529e-19, 
    2.550502e-19, 2.550512e-19, 2.550592e-19, 2.550389e-19, 2.550626e-19, 
    2.550663e-19, 2.550562e-19, 2.551168e-19, 2.550995e-19, 2.551172e-19, 
    2.55106e-19, 2.548247e-19, 2.548384e-19, 2.548309e-19, 2.548448e-19, 
    2.548348e-19, 2.548785e-19, 2.548916e-19, 2.549537e-19, 2.549288e-19, 
    2.549691e-19, 2.549331e-19, 2.549393e-19, 2.549694e-19, 2.549352e-19, 
    2.550129e-19, 2.549592e-19, 2.550595e-19, 2.550048e-19, 2.550629e-19, 
    2.550528e-19, 2.550699e-19, 2.550849e-19, 2.551043e-19, 2.551395e-19, 
    2.551315e-19, 2.551613e-19, 2.548591e-19, 2.548766e-19, 2.548755e-19, 
    2.548943e-19, 2.549081e-19, 2.549386e-19, 2.54987e-19, 2.549689e-19, 
    2.550026e-19, 2.550093e-19, 2.549583e-19, 2.549891e-19, 2.548888e-19, 
    2.549044e-19, 2.548955e-19, 2.548602e-19, 2.549724e-19, 2.549144e-19, 
    2.550221e-19, 2.549907e-19, 2.550827e-19, 2.550364e-19, 2.551269e-19, 
    2.551645e-19, 2.552022e-19, 2.552438e-19, 2.548868e-19, 2.548747e-19, 
    2.548967e-19, 2.549262e-19, 2.54955e-19, 2.549925e-19, 2.549966e-19, 
    2.550035e-19, 2.550221e-19, 2.550374e-19, 2.550053e-19, 2.550413e-19, 
    2.549071e-19, 2.549777e-19, 2.548698e-19, 2.549015e-19, 2.549247e-19, 
    2.54915e-19, 2.54967e-19, 2.549791e-19, 2.550282e-19, 2.550031e-19, 
    2.551548e-19, 2.550874e-19, 2.552771e-19, 2.552236e-19, 2.548704e-19, 
    2.548869e-19, 2.549438e-19, 2.549168e-19, 2.549953e-19, 2.550145e-19, 
    2.550305e-19, 2.550502e-19, 2.550527e-19, 2.550644e-19, 2.550451e-19, 
    2.550638e-19, 2.549926e-19, 2.550245e-19, 2.549378e-19, 2.549586e-19, 
    2.549492e-19, 2.549386e-19, 2.549714e-19, 2.550057e-19, 2.550072e-19, 
    2.55018e-19, 2.550473e-19, 2.549956e-19, 2.551621e-19, 2.550578e-19, 
    2.549049e-19, 2.549357e-19, 2.54941e-19, 2.549289e-19, 2.550125e-19, 
    2.549821e-19, 2.550642e-19, 2.550422e-19, 2.550785e-19, 2.550604e-19, 
    2.550577e-19, 2.550346e-19, 2.5502e-19, 2.549833e-19, 2.549538e-19, 
    2.549308e-19, 2.549362e-19, 2.549615e-19, 2.550079e-19, 2.550525e-19, 
    2.550427e-19, 2.550758e-19, 2.549896e-19, 2.550253e-19, 2.550112e-19, 
    2.55048e-19, 2.549683e-19, 2.550338e-19, 2.549513e-19, 2.549586e-19, 
    2.549815e-19, 2.550272e-19, 2.550384e-19, 2.550491e-19, 2.550427e-19, 
    2.550093e-19, 2.550041e-19, 2.549811e-19, 2.549744e-19, 2.549571e-19, 
    2.549425e-19, 2.549557e-19, 2.549694e-19, 2.550096e-19, 2.550455e-19, 
    2.55085e-19, 2.55095e-19, 2.551394e-19, 2.551022e-19, 2.551625e-19, 
    2.551096e-19, 2.552021e-19, 2.550388e-19, 2.551096e-19, 2.549828e-19, 
    2.549966e-19, 2.550208e-19, 2.55078e-19, 2.550479e-19, 2.550834e-19, 
    2.55004e-19, 2.54962e-19, 2.549521e-19, 2.54932e-19, 2.549525e-19, 
    2.549509e-19, 2.549705e-19, 2.549642e-19, 2.550109e-19, 2.549859e-19, 
    2.550574e-19, 2.550834e-19, 2.551579e-19, 2.552033e-19, 2.552508e-19, 
    2.552715e-19, 2.552778e-19, 2.552804e-19 ;

 MEG_acetone =
  8.502781e-17, 8.503699e-17, 8.503524e-17, 8.504256e-17, 8.503855e-17, 
    8.504331e-17, 8.502975e-17, 8.503728e-17, 8.503251e-17, 8.502874e-17, 
    8.505659e-17, 8.50429e-17, 8.507154e-17, 8.506266e-17, 8.508522e-17, 
    8.507006e-17, 8.508831e-17, 8.508495e-17, 8.509549e-17, 8.509248e-17, 
    8.510564e-17, 8.509689e-17, 8.511276e-17, 8.510364e-17, 8.5105e-17, 
    8.509657e-17, 8.504581e-17, 8.505483e-17, 8.504524e-17, 8.504653e-17, 
    8.504599e-17, 8.503858e-17, 8.503475e-17, 8.502723e-17, 8.502862e-17, 
    8.503421e-17, 8.504712e-17, 8.504284e-17, 8.505395e-17, 8.505371e-17, 
    8.5066e-17, 8.506045e-17, 8.50813e-17, 8.50754e-17, 8.509261e-17, 
    8.508824e-17, 8.509237e-17, 8.509114e-17, 8.509239e-17, 8.508601e-17, 
    8.508873e-17, 8.508318e-17, 8.506146e-17, 8.506777e-17, 8.504887e-17, 
    8.50373e-17, 8.503004e-17, 8.502478e-17, 8.502552e-17, 8.502691e-17, 
    8.503424e-17, 8.504128e-17, 8.504661e-17, 8.505015e-17, 8.505367e-17, 
    8.50639e-17, 8.506969e-17, 8.508241e-17, 8.508025e-17, 8.508402e-17, 
    8.508782e-17, 8.509402e-17, 8.509302e-17, 8.509572e-17, 8.508402e-17, 
    8.509174e-17, 8.507899e-17, 8.508245e-17, 8.505407e-17, 8.504402e-17, 
    8.503928e-17, 8.503556e-17, 8.502609e-17, 8.503259e-17, 8.503001e-17, 
    8.503627e-17, 8.504017e-17, 8.503826e-17, 8.505025e-17, 8.504556e-17, 
    8.507003e-17, 8.505948e-17, 8.508738e-17, 8.508071e-17, 8.5089e-17, 
    8.508479e-17, 8.509196e-17, 8.508551e-17, 8.509677e-17, 8.509916e-17, 
    8.509752e-17, 8.510404e-17, 8.508514e-17, 8.509232e-17, 8.503818e-17, 
    8.503849e-17, 8.503999e-17, 8.50334e-17, 8.503302e-17, 8.502717e-17, 
    8.503243e-17, 8.503463e-17, 8.504044e-17, 8.504378e-17, 8.504698e-17, 
    8.505407e-17, 8.506189e-17, 8.507302e-17, 8.508113e-17, 8.508655e-17, 
    8.508326e-17, 8.508616e-17, 8.50829e-17, 8.50814e-17, 8.509823e-17, 
    8.508872e-17, 8.51031e-17, 8.510233e-17, 8.509576e-17, 8.510241e-17, 
    8.503871e-17, 8.503693e-17, 8.503055e-17, 8.503554e-17, 8.502653e-17, 
    8.50315e-17, 8.503433e-17, 8.504554e-17, 8.504814e-17, 8.505039e-17, 
    8.505495e-17, 8.506073e-17, 8.507087e-17, 8.507981e-17, 8.508807e-17, 
    8.508747e-17, 8.508768e-17, 8.508946e-17, 8.508496e-17, 8.509021e-17, 
    8.509104e-17, 8.508879e-17, 8.510221e-17, 8.509838e-17, 8.510231e-17, 
    8.509983e-17, 8.503752e-17, 8.504056e-17, 8.503891e-17, 8.504198e-17, 
    8.503977e-17, 8.504944e-17, 8.505234e-17, 8.50661e-17, 8.506058e-17, 
    8.506952e-17, 8.506154e-17, 8.506291e-17, 8.506957e-17, 8.506201e-17, 
    8.507921e-17, 8.506732e-17, 8.508954e-17, 8.507741e-17, 8.509028e-17, 
    8.508803e-17, 8.509182e-17, 8.509515e-17, 8.509945e-17, 8.510724e-17, 
    8.510546e-17, 8.511207e-17, 8.504513e-17, 8.504902e-17, 8.504878e-17, 
    8.505295e-17, 8.505599e-17, 8.506274e-17, 8.507347e-17, 8.506946e-17, 
    8.507694e-17, 8.50784e-17, 8.506711e-17, 8.507394e-17, 8.505172e-17, 
    8.505519e-17, 8.50532e-17, 8.504538e-17, 8.507023e-17, 8.50574e-17, 
    8.508124e-17, 8.507429e-17, 8.509466e-17, 8.508441e-17, 8.510445e-17, 
    8.511278e-17, 8.512113e-17, 8.513033e-17, 8.505127e-17, 8.504861e-17, 
    8.505347e-17, 8.506e-17, 8.506637e-17, 8.507469e-17, 8.507561e-17, 
    8.507713e-17, 8.508123e-17, 8.508462e-17, 8.507752e-17, 8.508549e-17, 
    8.505579e-17, 8.507141e-17, 8.504751e-17, 8.505455e-17, 8.505966e-17, 
    8.505753e-17, 8.506903e-17, 8.507171e-17, 8.508259e-17, 8.507702e-17, 
    8.511062e-17, 8.50957e-17, 8.513772e-17, 8.512585e-17, 8.504765e-17, 
    8.505131e-17, 8.506389e-17, 8.505792e-17, 8.507531e-17, 8.507955e-17, 
    8.50831e-17, 8.508746e-17, 8.508801e-17, 8.509061e-17, 8.508633e-17, 
    8.509048e-17, 8.507471e-17, 8.508177e-17, 8.506258e-17, 8.506717e-17, 
    8.50651e-17, 8.506274e-17, 8.507001e-17, 8.50776e-17, 8.507793e-17, 
    8.508034e-17, 8.508682e-17, 8.507538e-17, 8.511224e-17, 8.508914e-17, 
    8.505529e-17, 8.506211e-17, 8.506328e-17, 8.506061e-17, 8.507912e-17, 
    8.507238e-17, 8.509057e-17, 8.508568e-17, 8.509374e-17, 8.508972e-17, 
    8.508912e-17, 8.5084e-17, 8.508077e-17, 8.507265e-17, 8.506611e-17, 
    8.506101e-17, 8.506221e-17, 8.506781e-17, 8.507811e-17, 8.508798e-17, 
    8.508579e-17, 8.509313e-17, 8.507404e-17, 8.508194e-17, 8.507883e-17, 
    8.508698e-17, 8.506932e-17, 8.508384e-17, 8.506555e-17, 8.506719e-17, 
    8.507225e-17, 8.508236e-17, 8.508486e-17, 8.508722e-17, 8.50858e-17, 
    8.50784e-17, 8.507726e-17, 8.507216e-17, 8.507067e-17, 8.506684e-17, 
    8.50636e-17, 8.506653e-17, 8.506956e-17, 8.507847e-17, 8.508642e-17, 
    8.509517e-17, 8.509738e-17, 8.510721e-17, 8.509897e-17, 8.511234e-17, 
    8.510062e-17, 8.512111e-17, 8.508494e-17, 8.510061e-17, 8.507253e-17, 
    8.507559e-17, 8.508095e-17, 8.509361e-17, 8.508695e-17, 8.509483e-17, 
    8.507723e-17, 8.506792e-17, 8.506573e-17, 8.50613e-17, 8.506583e-17, 
    8.506547e-17, 8.50698e-17, 8.506842e-17, 8.507877e-17, 8.507322e-17, 
    8.508906e-17, 8.509481e-17, 8.511131e-17, 8.512137e-17, 8.51319e-17, 
    8.513647e-17, 8.513788e-17, 8.513845e-17 ;

 MEG_carene_3 =
  3.286486e-17, 3.286848e-17, 3.286779e-17, 3.287068e-17, 3.28691e-17, 
    3.287097e-17, 3.286562e-17, 3.28686e-17, 3.286671e-17, 3.286523e-17, 
    3.287621e-17, 3.287081e-17, 3.288211e-17, 3.287861e-17, 3.288751e-17, 
    3.288153e-17, 3.288873e-17, 3.28874e-17, 3.289156e-17, 3.289037e-17, 
    3.289557e-17, 3.289211e-17, 3.289837e-17, 3.289478e-17, 3.289531e-17, 
    3.289199e-17, 3.287196e-17, 3.287552e-17, 3.287173e-17, 3.287225e-17, 
    3.287203e-17, 3.286911e-17, 3.286759e-17, 3.286463e-17, 3.286518e-17, 
    3.286738e-17, 3.287248e-17, 3.287079e-17, 3.287518e-17, 3.287508e-17, 
    3.287993e-17, 3.287774e-17, 3.288596e-17, 3.288364e-17, 3.289042e-17, 
    3.28887e-17, 3.289033e-17, 3.288985e-17, 3.289034e-17, 3.288782e-17, 
    3.28889e-17, 3.28867e-17, 3.287813e-17, 3.288062e-17, 3.287317e-17, 
    3.28686e-17, 3.286574e-17, 3.286366e-17, 3.286396e-17, 3.28645e-17, 
    3.28674e-17, 3.287017e-17, 3.287228e-17, 3.287368e-17, 3.287506e-17, 
    3.28791e-17, 3.288138e-17, 3.28864e-17, 3.288555e-17, 3.288704e-17, 
    3.288854e-17, 3.289098e-17, 3.289059e-17, 3.289165e-17, 3.288704e-17, 
    3.289008e-17, 3.288505e-17, 3.288642e-17, 3.287522e-17, 3.287125e-17, 
    3.286938e-17, 3.286792e-17, 3.286418e-17, 3.286674e-17, 3.286573e-17, 
    3.28682e-17, 3.286974e-17, 3.286898e-17, 3.287371e-17, 3.287186e-17, 
    3.288151e-17, 3.287736e-17, 3.288836e-17, 3.288573e-17, 3.2889e-17, 
    3.288734e-17, 3.289017e-17, 3.288763e-17, 3.289207e-17, 3.289301e-17, 
    3.289236e-17, 3.289493e-17, 3.288748e-17, 3.289031e-17, 3.286895e-17, 
    3.286907e-17, 3.286966e-17, 3.286706e-17, 3.286692e-17, 3.28646e-17, 
    3.286668e-17, 3.286755e-17, 3.286984e-17, 3.287116e-17, 3.287243e-17, 
    3.287522e-17, 3.287831e-17, 3.28827e-17, 3.28859e-17, 3.288803e-17, 
    3.288674e-17, 3.288788e-17, 3.28866e-17, 3.2886e-17, 3.289264e-17, 
    3.288889e-17, 3.289456e-17, 3.289426e-17, 3.289167e-17, 3.289429e-17, 
    3.286916e-17, 3.286846e-17, 3.286594e-17, 3.286791e-17, 3.286436e-17, 
    3.286632e-17, 3.286743e-17, 3.287185e-17, 3.287288e-17, 3.287377e-17, 
    3.287557e-17, 3.287785e-17, 3.288185e-17, 3.288538e-17, 3.288863e-17, 
    3.28884e-17, 3.288848e-17, 3.288918e-17, 3.288741e-17, 3.288948e-17, 
    3.288981e-17, 3.288892e-17, 3.289421e-17, 3.28927e-17, 3.289425e-17, 
    3.289327e-17, 3.286869e-17, 3.286989e-17, 3.286924e-17, 3.287045e-17, 
    3.286958e-17, 3.287339e-17, 3.287454e-17, 3.287997e-17, 3.287779e-17, 
    3.288131e-17, 3.287817e-17, 3.287871e-17, 3.288134e-17, 3.287835e-17, 
    3.288514e-17, 3.288045e-17, 3.288921e-17, 3.288443e-17, 3.288951e-17, 
    3.288862e-17, 3.289011e-17, 3.289143e-17, 3.289312e-17, 3.28962e-17, 
    3.289549e-17, 3.28981e-17, 3.287169e-17, 3.287323e-17, 3.287314e-17, 
    3.287477e-17, 3.287598e-17, 3.287864e-17, 3.288287e-17, 3.288129e-17, 
    3.288424e-17, 3.288482e-17, 3.288037e-17, 3.288306e-17, 3.287429e-17, 
    3.287566e-17, 3.287488e-17, 3.287179e-17, 3.28816e-17, 3.287653e-17, 
    3.288594e-17, 3.28832e-17, 3.289123e-17, 3.288719e-17, 3.28951e-17, 
    3.289838e-17, 3.290168e-17, 3.290531e-17, 3.287412e-17, 3.287306e-17, 
    3.287498e-17, 3.287756e-17, 3.288007e-17, 3.288336e-17, 3.288371e-17, 
    3.288432e-17, 3.288594e-17, 3.288728e-17, 3.288447e-17, 3.288762e-17, 
    3.28759e-17, 3.288206e-17, 3.287263e-17, 3.287541e-17, 3.287743e-17, 
    3.287658e-17, 3.288112e-17, 3.288218e-17, 3.288647e-17, 3.288428e-17, 
    3.289753e-17, 3.289165e-17, 3.290822e-17, 3.290354e-17, 3.287269e-17, 
    3.287413e-17, 3.28791e-17, 3.287674e-17, 3.28836e-17, 3.288527e-17, 
    3.288667e-17, 3.288839e-17, 3.288861e-17, 3.288964e-17, 3.288795e-17, 
    3.288958e-17, 3.288336e-17, 3.288615e-17, 3.287858e-17, 3.288039e-17, 
    3.287957e-17, 3.287864e-17, 3.288151e-17, 3.28845e-17, 3.288463e-17, 
    3.288558e-17, 3.288814e-17, 3.288363e-17, 3.289817e-17, 3.288906e-17, 
    3.28757e-17, 3.287839e-17, 3.287885e-17, 3.28778e-17, 3.28851e-17, 
    3.288244e-17, 3.288962e-17, 3.288769e-17, 3.289087e-17, 3.288928e-17, 
    3.288905e-17, 3.288703e-17, 3.288575e-17, 3.288255e-17, 3.287997e-17, 
    3.287796e-17, 3.287843e-17, 3.288064e-17, 3.28847e-17, 3.28886e-17, 
    3.288774e-17, 3.289063e-17, 3.28831e-17, 3.288622e-17, 3.288499e-17, 
    3.28882e-17, 3.288124e-17, 3.288696e-17, 3.287975e-17, 3.28804e-17, 
    3.288239e-17, 3.288638e-17, 3.288737e-17, 3.28883e-17, 3.288774e-17, 
    3.288482e-17, 3.288437e-17, 3.288236e-17, 3.288177e-17, 3.288026e-17, 
    3.287898e-17, 3.288013e-17, 3.288133e-17, 3.288485e-17, 3.288798e-17, 
    3.289143e-17, 3.289231e-17, 3.289619e-17, 3.289294e-17, 3.289821e-17, 
    3.289358e-17, 3.290167e-17, 3.28874e-17, 3.289358e-17, 3.288251e-17, 
    3.288371e-17, 3.288582e-17, 3.289082e-17, 3.288819e-17, 3.28913e-17, 
    3.288436e-17, 3.288068e-17, 3.287982e-17, 3.287807e-17, 3.287986e-17, 
    3.287972e-17, 3.288143e-17, 3.288088e-17, 3.288497e-17, 3.288278e-17, 
    3.288903e-17, 3.289129e-17, 3.28978e-17, 3.290177e-17, 3.290593e-17, 
    3.290773e-17, 3.290828e-17, 3.290851e-17 ;

 MEG_ethanol =
  1.698539e-18, 1.698815e-18, 1.698762e-18, 1.698983e-18, 1.698862e-18, 
    1.699005e-18, 1.698597e-18, 1.698824e-18, 1.69868e-18, 1.698567e-18, 
    1.699405e-18, 1.698993e-18, 1.699856e-18, 1.699588e-18, 1.700267e-18, 
    1.699811e-18, 1.70036e-18, 1.700259e-18, 1.700576e-18, 1.700486e-18, 
    1.700882e-18, 1.700618e-18, 1.701096e-18, 1.700822e-18, 1.700863e-18, 
    1.700609e-18, 1.699081e-18, 1.699352e-18, 1.699063e-18, 1.699102e-18, 
    1.699086e-18, 1.698863e-18, 1.698748e-18, 1.698521e-18, 1.698563e-18, 
    1.698731e-18, 1.69912e-18, 1.698991e-18, 1.699326e-18, 1.699318e-18, 
    1.699689e-18, 1.699521e-18, 1.700149e-18, 1.699972e-18, 1.70049e-18, 
    1.700358e-18, 1.700483e-18, 1.700446e-18, 1.700483e-18, 1.700291e-18, 
    1.700373e-18, 1.700206e-18, 1.699552e-18, 1.699742e-18, 1.699173e-18, 
    1.698825e-18, 1.698606e-18, 1.698447e-18, 1.69847e-18, 1.698511e-18, 
    1.698732e-18, 1.698944e-18, 1.699105e-18, 1.699211e-18, 1.699317e-18, 
    1.699625e-18, 1.6998e-18, 1.700183e-18, 1.700118e-18, 1.700231e-18, 
    1.700346e-18, 1.700532e-18, 1.700502e-18, 1.700583e-18, 1.700231e-18, 
    1.700464e-18, 1.70008e-18, 1.700184e-18, 1.699329e-18, 1.699027e-18, 
    1.698884e-18, 1.698772e-18, 1.698487e-18, 1.698683e-18, 1.698605e-18, 
    1.698793e-18, 1.698911e-18, 1.698853e-18, 1.699214e-18, 1.699073e-18, 
    1.69981e-18, 1.699492e-18, 1.700332e-18, 1.700131e-18, 1.700381e-18, 
    1.700254e-18, 1.70047e-18, 1.700276e-18, 1.700615e-18, 1.700687e-18, 
    1.700637e-18, 1.700834e-18, 1.700265e-18, 1.700481e-18, 1.698851e-18, 
    1.69886e-18, 1.698905e-18, 1.698707e-18, 1.698696e-18, 1.698519e-18, 
    1.698678e-18, 1.698744e-18, 1.698919e-18, 1.699019e-18, 1.699116e-18, 
    1.699329e-18, 1.699565e-18, 1.6999e-18, 1.700144e-18, 1.700307e-18, 
    1.700208e-18, 1.700296e-18, 1.700197e-18, 1.700152e-18, 1.700659e-18, 
    1.700373e-18, 1.700806e-18, 1.700782e-18, 1.700585e-18, 1.700785e-18, 
    1.698867e-18, 1.698813e-18, 1.698621e-18, 1.698772e-18, 1.6985e-18, 
    1.69865e-18, 1.698735e-18, 1.699072e-18, 1.699151e-18, 1.699218e-18, 
    1.699356e-18, 1.69953e-18, 1.699835e-18, 1.700104e-18, 1.700353e-18, 
    1.700335e-18, 1.700341e-18, 1.700395e-18, 1.700259e-18, 1.700417e-18, 
    1.700442e-18, 1.700375e-18, 1.700779e-18, 1.700663e-18, 1.700782e-18, 
    1.700707e-18, 1.698831e-18, 1.698922e-18, 1.698873e-18, 1.698965e-18, 
    1.698899e-18, 1.69919e-18, 1.699277e-18, 1.699691e-18, 1.699526e-18, 
    1.699794e-18, 1.699554e-18, 1.699596e-18, 1.699796e-18, 1.699568e-18, 
    1.700086e-18, 1.699728e-18, 1.700397e-18, 1.700032e-18, 1.70042e-18, 
    1.700352e-18, 1.700466e-18, 1.700566e-18, 1.700696e-18, 1.70093e-18, 
    1.700876e-18, 1.701075e-18, 1.69906e-18, 1.699177e-18, 1.69917e-18, 
    1.699295e-18, 1.699387e-18, 1.69959e-18, 1.699913e-18, 1.699793e-18, 
    1.700018e-18, 1.700062e-18, 1.699722e-18, 1.699928e-18, 1.699259e-18, 
    1.699363e-18, 1.699303e-18, 1.699068e-18, 1.699816e-18, 1.69943e-18, 
    1.700148e-18, 1.699938e-18, 1.700551e-18, 1.700243e-18, 1.700846e-18, 
    1.701097e-18, 1.701348e-18, 1.701625e-18, 1.699245e-18, 1.699165e-18, 
    1.699311e-18, 1.699508e-18, 1.6997e-18, 1.69995e-18, 1.699978e-18, 
    1.700024e-18, 1.700147e-18, 1.700249e-18, 1.700035e-18, 1.700275e-18, 
    1.699381e-18, 1.699851e-18, 1.699132e-18, 1.699344e-18, 1.699498e-18, 
    1.699433e-18, 1.69978e-18, 1.699861e-18, 1.700188e-18, 1.70002e-18, 
    1.701032e-18, 1.700583e-18, 1.701847e-18, 1.70149e-18, 1.699136e-18, 
    1.699246e-18, 1.699625e-18, 1.699445e-18, 1.699969e-18, 1.700096e-18, 
    1.700203e-18, 1.700335e-18, 1.700351e-18, 1.700429e-18, 1.700301e-18, 
    1.700426e-18, 1.699951e-18, 1.700163e-18, 1.699586e-18, 1.699724e-18, 
    1.699661e-18, 1.69959e-18, 1.699809e-18, 1.700038e-18, 1.700048e-18, 
    1.70012e-18, 1.700315e-18, 1.699971e-18, 1.701081e-18, 1.700385e-18, 
    1.699366e-18, 1.699571e-18, 1.699607e-18, 1.699526e-18, 1.700084e-18, 
    1.699881e-18, 1.700428e-18, 1.700281e-18, 1.700524e-18, 1.700403e-18, 
    1.700385e-18, 1.700231e-18, 1.700133e-18, 1.699889e-18, 1.699692e-18, 
    1.699539e-18, 1.699575e-18, 1.699743e-18, 1.700053e-18, 1.70035e-18, 
    1.700284e-18, 1.700505e-18, 1.699931e-18, 1.700169e-18, 1.700075e-18, 
    1.70032e-18, 1.699788e-18, 1.700226e-18, 1.699675e-18, 1.699724e-18, 
    1.699877e-18, 1.700181e-18, 1.700256e-18, 1.700327e-18, 1.700285e-18, 
    1.700062e-18, 1.700028e-18, 1.699874e-18, 1.699829e-18, 1.699714e-18, 
    1.699616e-18, 1.699704e-18, 1.699796e-18, 1.700064e-18, 1.700303e-18, 
    1.700567e-18, 1.700633e-18, 1.700929e-18, 1.700681e-18, 1.701083e-18, 
    1.700731e-18, 1.701347e-18, 1.700259e-18, 1.700731e-18, 1.699885e-18, 
    1.699977e-18, 1.700138e-18, 1.70052e-18, 1.700319e-18, 1.700556e-18, 
    1.700027e-18, 1.699746e-18, 1.69968e-18, 1.699547e-18, 1.699683e-18, 
    1.699673e-18, 1.699803e-18, 1.699761e-18, 1.700073e-18, 1.699906e-18, 
    1.700383e-18, 1.700556e-18, 1.701053e-18, 1.701355e-18, 1.701672e-18, 
    1.70181e-18, 1.701852e-18, 1.70187e-18 ;

 MEG_formaldehyde =
  3.397077e-19, 3.39763e-19, 3.397525e-19, 3.397965e-19, 3.397724e-19, 
    3.39801e-19, 3.397194e-19, 3.397648e-19, 3.39736e-19, 3.397133e-19, 
    3.39881e-19, 3.397986e-19, 3.399711e-19, 3.399176e-19, 3.400534e-19, 
    3.399622e-19, 3.40072e-19, 3.400518e-19, 3.401153e-19, 3.400971e-19, 
    3.401764e-19, 3.401237e-19, 3.402192e-19, 3.401643e-19, 3.401725e-19, 
    3.401218e-19, 3.398161e-19, 3.398704e-19, 3.398127e-19, 3.398205e-19, 
    3.398172e-19, 3.397726e-19, 3.397495e-19, 3.397042e-19, 3.397126e-19, 
    3.397462e-19, 3.39824e-19, 3.397982e-19, 3.398652e-19, 3.398637e-19, 
    3.399377e-19, 3.399043e-19, 3.400298e-19, 3.399943e-19, 3.400979e-19, 
    3.400717e-19, 3.400965e-19, 3.400891e-19, 3.400966e-19, 3.400582e-19, 
    3.400746e-19, 3.400411e-19, 3.399104e-19, 3.399484e-19, 3.398346e-19, 
    3.397649e-19, 3.397212e-19, 3.396895e-19, 3.396939e-19, 3.397023e-19, 
    3.397464e-19, 3.397888e-19, 3.398209e-19, 3.398423e-19, 3.398635e-19, 
    3.39925e-19, 3.399599e-19, 3.400365e-19, 3.400235e-19, 3.400462e-19, 
    3.400691e-19, 3.401064e-19, 3.401004e-19, 3.401167e-19, 3.400462e-19, 
    3.400927e-19, 3.400159e-19, 3.400368e-19, 3.398658e-19, 3.398053e-19, 
    3.397768e-19, 3.397544e-19, 3.396973e-19, 3.397365e-19, 3.39721e-19, 
    3.397586e-19, 3.397821e-19, 3.397707e-19, 3.398429e-19, 3.398146e-19, 
    3.39962e-19, 3.398984e-19, 3.400664e-19, 3.400263e-19, 3.400762e-19, 
    3.400509e-19, 3.40094e-19, 3.400552e-19, 3.40123e-19, 3.401374e-19, 
    3.401275e-19, 3.401667e-19, 3.400529e-19, 3.400962e-19, 3.397702e-19, 
    3.39772e-19, 3.397811e-19, 3.397414e-19, 3.397391e-19, 3.397038e-19, 
    3.397355e-19, 3.397488e-19, 3.397838e-19, 3.398039e-19, 3.398232e-19, 
    3.398658e-19, 3.39913e-19, 3.3998e-19, 3.400288e-19, 3.400614e-19, 
    3.400417e-19, 3.400591e-19, 3.400395e-19, 3.400304e-19, 3.401318e-19, 
    3.400745e-19, 3.401611e-19, 3.401564e-19, 3.401169e-19, 3.401569e-19, 
    3.397734e-19, 3.397626e-19, 3.397242e-19, 3.397543e-19, 3.397e-19, 
    3.3973e-19, 3.397469e-19, 3.398145e-19, 3.398301e-19, 3.398437e-19, 
    3.398711e-19, 3.39906e-19, 3.399671e-19, 3.400209e-19, 3.400706e-19, 
    3.40067e-19, 3.400682e-19, 3.40079e-19, 3.400519e-19, 3.400835e-19, 
    3.400885e-19, 3.400749e-19, 3.401558e-19, 3.401327e-19, 3.401563e-19, 
    3.401414e-19, 3.397662e-19, 3.397845e-19, 3.397745e-19, 3.39793e-19, 
    3.397797e-19, 3.39838e-19, 3.398554e-19, 3.399383e-19, 3.399051e-19, 
    3.399589e-19, 3.399108e-19, 3.399191e-19, 3.399592e-19, 3.399136e-19, 
    3.400172e-19, 3.399457e-19, 3.400794e-19, 3.400064e-19, 3.400839e-19, 
    3.400703e-19, 3.400931e-19, 3.401132e-19, 3.401391e-19, 3.40186e-19, 
    3.401753e-19, 3.402151e-19, 3.398121e-19, 3.398355e-19, 3.39834e-19, 
    3.398591e-19, 3.398775e-19, 3.399181e-19, 3.399827e-19, 3.399585e-19, 
    3.400035e-19, 3.400124e-19, 3.399444e-19, 3.399855e-19, 3.398517e-19, 
    3.398726e-19, 3.398606e-19, 3.398135e-19, 3.399632e-19, 3.398859e-19, 
    3.400295e-19, 3.399876e-19, 3.401102e-19, 3.400485e-19, 3.401692e-19, 
    3.402193e-19, 3.402696e-19, 3.40325e-19, 3.39849e-19, 3.39833e-19, 
    3.398623e-19, 3.399016e-19, 3.399399e-19, 3.399901e-19, 3.399955e-19, 
    3.400047e-19, 3.400294e-19, 3.400498e-19, 3.40007e-19, 3.40055e-19, 
    3.398762e-19, 3.399703e-19, 3.398263e-19, 3.398687e-19, 3.398995e-19, 
    3.398867e-19, 3.39956e-19, 3.399721e-19, 3.400376e-19, 3.400041e-19, 
    3.402064e-19, 3.401166e-19, 3.403694e-19, 3.40298e-19, 3.398272e-19, 
    3.398492e-19, 3.39925e-19, 3.398891e-19, 3.399937e-19, 3.400193e-19, 
    3.400406e-19, 3.400669e-19, 3.400702e-19, 3.400859e-19, 3.400602e-19, 
    3.400851e-19, 3.399902e-19, 3.400326e-19, 3.399171e-19, 3.399448e-19, 
    3.399323e-19, 3.399181e-19, 3.399618e-19, 3.400076e-19, 3.400096e-19, 
    3.40024e-19, 3.400631e-19, 3.399942e-19, 3.402161e-19, 3.40077e-19, 
    3.398732e-19, 3.399142e-19, 3.399214e-19, 3.399052e-19, 3.400167e-19, 
    3.399761e-19, 3.400856e-19, 3.400562e-19, 3.401047e-19, 3.400805e-19, 
    3.400769e-19, 3.400461e-19, 3.400267e-19, 3.399778e-19, 3.399384e-19, 
    3.399077e-19, 3.399149e-19, 3.399486e-19, 3.400106e-19, 3.400701e-19, 
    3.400569e-19, 3.40101e-19, 3.399861e-19, 3.400337e-19, 3.400149e-19, 
    3.400641e-19, 3.399577e-19, 3.400451e-19, 3.39935e-19, 3.399449e-19, 
    3.399753e-19, 3.400362e-19, 3.400513e-19, 3.400655e-19, 3.400569e-19, 
    3.400124e-19, 3.400055e-19, 3.399749e-19, 3.399658e-19, 3.399428e-19, 
    3.399233e-19, 3.399409e-19, 3.399591e-19, 3.400128e-19, 3.400607e-19, 
    3.401133e-19, 3.401267e-19, 3.401858e-19, 3.401362e-19, 3.402167e-19, 
    3.401461e-19, 3.402695e-19, 3.400517e-19, 3.401461e-19, 3.399771e-19, 
    3.399955e-19, 3.400277e-19, 3.40104e-19, 3.400638e-19, 3.401113e-19, 
    3.400053e-19, 3.399493e-19, 3.399361e-19, 3.399094e-19, 3.399367e-19, 
    3.399345e-19, 3.399606e-19, 3.399523e-19, 3.400146e-19, 3.399812e-19, 
    3.400765e-19, 3.401112e-19, 3.402105e-19, 3.40271e-19, 3.403344e-19, 
    3.403619e-19, 3.403704e-19, 3.403739e-19 ;

 MEG_isoprene =
  2.334197e-19, 2.334649e-19, 2.334563e-19, 2.334924e-19, 2.334727e-19, 
    2.334961e-19, 2.334293e-19, 2.334664e-19, 2.334429e-19, 2.334243e-19, 
    2.335616e-19, 2.334941e-19, 2.336353e-19, 2.335915e-19, 2.337027e-19, 
    2.33628e-19, 2.337179e-19, 2.337014e-19, 2.337533e-19, 2.337385e-19, 
    2.338033e-19, 2.337602e-19, 2.338384e-19, 2.337935e-19, 2.338002e-19, 
    2.337587e-19, 2.335084e-19, 2.335529e-19, 2.335056e-19, 2.33512e-19, 
    2.335093e-19, 2.334728e-19, 2.334539e-19, 2.334168e-19, 2.334237e-19, 
    2.334513e-19, 2.335149e-19, 2.334938e-19, 2.335486e-19, 2.335474e-19, 
    2.33608e-19, 2.335806e-19, 2.336834e-19, 2.336543e-19, 2.337391e-19, 
    2.337176e-19, 2.33738e-19, 2.337319e-19, 2.337381e-19, 2.337066e-19, 
    2.3372e-19, 2.336926e-19, 2.335856e-19, 2.336167e-19, 2.335235e-19, 
    2.334665e-19, 2.334307e-19, 2.334048e-19, 2.334084e-19, 2.334153e-19, 
    2.334514e-19, 2.334861e-19, 2.335124e-19, 2.335299e-19, 2.335472e-19, 
    2.335976e-19, 2.336262e-19, 2.336889e-19, 2.336782e-19, 2.336968e-19, 
    2.337155e-19, 2.337461e-19, 2.337412e-19, 2.337545e-19, 2.336968e-19, 
    2.337348e-19, 2.33672e-19, 2.336891e-19, 2.335491e-19, 2.334996e-19, 
    2.334762e-19, 2.334579e-19, 2.334112e-19, 2.334433e-19, 2.334305e-19, 
    2.334614e-19, 2.334806e-19, 2.334712e-19, 2.335304e-19, 2.335072e-19, 
    2.336278e-19, 2.335758e-19, 2.337133e-19, 2.336805e-19, 2.337213e-19, 
    2.337006e-19, 2.337359e-19, 2.337042e-19, 2.337597e-19, 2.337715e-19, 
    2.337633e-19, 2.337955e-19, 2.337023e-19, 2.337377e-19, 2.334708e-19, 
    2.334723e-19, 2.334797e-19, 2.334472e-19, 2.334454e-19, 2.334165e-19, 
    2.334425e-19, 2.334533e-19, 2.33482e-19, 2.334984e-19, 2.335143e-19, 
    2.335492e-19, 2.335877e-19, 2.336426e-19, 2.336826e-19, 2.337093e-19, 
    2.336931e-19, 2.337073e-19, 2.336913e-19, 2.336839e-19, 2.337668e-19, 
    2.3372e-19, 2.337908e-19, 2.33787e-19, 2.337547e-19, 2.337874e-19, 
    2.334735e-19, 2.334647e-19, 2.334332e-19, 2.334578e-19, 2.334134e-19, 
    2.334379e-19, 2.334518e-19, 2.335071e-19, 2.335199e-19, 2.33531e-19, 
    2.335535e-19, 2.33582e-19, 2.33632e-19, 2.33676e-19, 2.337168e-19, 
    2.337138e-19, 2.337148e-19, 2.337236e-19, 2.337014e-19, 2.337273e-19, 
    2.337314e-19, 2.337203e-19, 2.337865e-19, 2.337676e-19, 2.337869e-19, 
    2.337747e-19, 2.334676e-19, 2.334826e-19, 2.334744e-19, 2.334896e-19, 
    2.334787e-19, 2.335263e-19, 2.335406e-19, 2.336084e-19, 2.335813e-19, 
    2.336253e-19, 2.33586e-19, 2.335928e-19, 2.336256e-19, 2.335883e-19, 
    2.336731e-19, 2.336145e-19, 2.33724e-19, 2.336642e-19, 2.337277e-19, 
    2.337166e-19, 2.337352e-19, 2.337517e-19, 2.337728e-19, 2.338112e-19, 
    2.338024e-19, 2.33835e-19, 2.335051e-19, 2.335243e-19, 2.335231e-19, 
    2.335436e-19, 2.335587e-19, 2.335919e-19, 2.336448e-19, 2.33625e-19, 
    2.336619e-19, 2.336691e-19, 2.336135e-19, 2.336471e-19, 2.335376e-19, 
    2.335547e-19, 2.335449e-19, 2.335063e-19, 2.336289e-19, 2.335656e-19, 
    2.336831e-19, 2.336488e-19, 2.337492e-19, 2.336987e-19, 2.337975e-19, 
    2.338385e-19, 2.338797e-19, 2.33925e-19, 2.335354e-19, 2.335222e-19, 
    2.335462e-19, 2.335784e-19, 2.336098e-19, 2.336508e-19, 2.336553e-19, 
    2.336629e-19, 2.33683e-19, 2.336998e-19, 2.336647e-19, 2.33704e-19, 
    2.335576e-19, 2.336346e-19, 2.335168e-19, 2.335515e-19, 2.335767e-19, 
    2.335662e-19, 2.336229e-19, 2.336362e-19, 2.336897e-19, 2.336623e-19, 
    2.338279e-19, 2.337544e-19, 2.339614e-19, 2.339029e-19, 2.335175e-19, 
    2.335356e-19, 2.335976e-19, 2.335681e-19, 2.336539e-19, 2.336748e-19, 
    2.336922e-19, 2.337138e-19, 2.337164e-19, 2.337293e-19, 2.337082e-19, 
    2.337286e-19, 2.336509e-19, 2.336857e-19, 2.335911e-19, 2.336138e-19, 
    2.336035e-19, 2.335919e-19, 2.336277e-19, 2.336652e-19, 2.336668e-19, 
    2.336787e-19, 2.337106e-19, 2.336542e-19, 2.338359e-19, 2.33722e-19, 
    2.335552e-19, 2.335888e-19, 2.335946e-19, 2.335814e-19, 2.336726e-19, 
    2.336394e-19, 2.337291e-19, 2.33705e-19, 2.337447e-19, 2.337249e-19, 
    2.337219e-19, 2.336967e-19, 2.336808e-19, 2.336408e-19, 2.336085e-19, 
    2.335834e-19, 2.335893e-19, 2.336169e-19, 2.336676e-19, 2.337163e-19, 
    2.337055e-19, 2.337417e-19, 2.336476e-19, 2.336866e-19, 2.336712e-19, 
    2.337114e-19, 2.336243e-19, 2.336959e-19, 2.336058e-19, 2.336138e-19, 
    2.336388e-19, 2.336886e-19, 2.337009e-19, 2.337126e-19, 2.337056e-19, 
    2.336691e-19, 2.336635e-19, 2.336384e-19, 2.33631e-19, 2.336122e-19, 
    2.335962e-19, 2.336106e-19, 2.336255e-19, 2.336694e-19, 2.337086e-19, 
    2.337518e-19, 2.337626e-19, 2.338111e-19, 2.337705e-19, 2.338363e-19, 
    2.337786e-19, 2.338796e-19, 2.337013e-19, 2.337786e-19, 2.336402e-19, 
    2.336553e-19, 2.336817e-19, 2.337441e-19, 2.337112e-19, 2.337501e-19, 
    2.336633e-19, 2.336174e-19, 2.336067e-19, 2.335848e-19, 2.336072e-19, 
    2.336054e-19, 2.336267e-19, 2.336199e-19, 2.336709e-19, 2.336436e-19, 
    2.337216e-19, 2.3375e-19, 2.338313e-19, 2.338808e-19, 2.339327e-19, 
    2.339552e-19, 2.339621e-19, 2.33965e-19 ;

 MEG_methanol =
  5.843022e-17, 5.843617e-17, 5.843504e-17, 5.843978e-17, 5.843719e-17, 
    5.844026e-17, 5.843147e-17, 5.843636e-17, 5.843326e-17, 5.843082e-17, 
    5.844888e-17, 5.844001e-17, 5.845859e-17, 5.845282e-17, 5.846746e-17, 
    5.845762e-17, 5.846946e-17, 5.846728e-17, 5.847412e-17, 5.847217e-17, 
    5.84807e-17, 5.847502e-17, 5.848532e-17, 5.84794e-17, 5.848029e-17, 
    5.847481e-17, 5.844189e-17, 5.844774e-17, 5.844152e-17, 5.844236e-17, 
    5.8442e-17, 5.843721e-17, 5.843471e-17, 5.842983e-17, 5.843074e-17, 
    5.843437e-17, 5.844274e-17, 5.843997e-17, 5.844718e-17, 5.844701e-17, 
    5.845499e-17, 5.845139e-17, 5.846491e-17, 5.846109e-17, 5.847225e-17, 
    5.846942e-17, 5.847209e-17, 5.84713e-17, 5.847211e-17, 5.846796e-17, 
    5.846973e-17, 5.846613e-17, 5.845204e-17, 5.845614e-17, 5.844388e-17, 
    5.843637e-17, 5.843167e-17, 5.842825e-17, 5.842873e-17, 5.842963e-17, 
    5.843439e-17, 5.843895e-17, 5.844241e-17, 5.844471e-17, 5.844699e-17, 
    5.845362e-17, 5.845738e-17, 5.846564e-17, 5.846423e-17, 5.846667e-17, 
    5.846914e-17, 5.847317e-17, 5.847252e-17, 5.847426e-17, 5.846668e-17, 
    5.847168e-17, 5.846342e-17, 5.846566e-17, 5.844725e-17, 5.844073e-17, 
    5.843766e-17, 5.843524e-17, 5.842909e-17, 5.843332e-17, 5.843164e-17, 
    5.84357e-17, 5.843823e-17, 5.843699e-17, 5.844478e-17, 5.844173e-17, 
    5.84576e-17, 5.845076e-17, 5.846886e-17, 5.846453e-17, 5.84699e-17, 
    5.846718e-17, 5.847182e-17, 5.846765e-17, 5.847495e-17, 5.84765e-17, 
    5.847544e-17, 5.847966e-17, 5.84674e-17, 5.847206e-17, 5.843694e-17, 
    5.843714e-17, 5.843811e-17, 5.843384e-17, 5.84336e-17, 5.84298e-17, 
    5.843321e-17, 5.843464e-17, 5.843841e-17, 5.844057e-17, 5.844265e-17, 
    5.844725e-17, 5.845233e-17, 5.845955e-17, 5.846481e-17, 5.846832e-17, 
    5.846619e-17, 5.846806e-17, 5.846595e-17, 5.846498e-17, 5.847589e-17, 
    5.846973e-17, 5.847906e-17, 5.847855e-17, 5.84743e-17, 5.847861e-17, 
    5.843729e-17, 5.843613e-17, 5.843199e-17, 5.843523e-17, 5.842938e-17, 
    5.843261e-17, 5.843444e-17, 5.844171e-17, 5.844341e-17, 5.844486e-17, 
    5.844781e-17, 5.845157e-17, 5.845815e-17, 5.846395e-17, 5.84693e-17, 
    5.846892e-17, 5.846905e-17, 5.847021e-17, 5.846729e-17, 5.847069e-17, 
    5.847123e-17, 5.846977e-17, 5.847848e-17, 5.847599e-17, 5.847854e-17, 
    5.847692e-17, 5.843652e-17, 5.843848e-17, 5.843742e-17, 5.84394e-17, 
    5.843797e-17, 5.844425e-17, 5.844613e-17, 5.845505e-17, 5.845148e-17, 
    5.845727e-17, 5.84521e-17, 5.845299e-17, 5.84573e-17, 5.84524e-17, 
    5.846356e-17, 5.845585e-17, 5.847025e-17, 5.846239e-17, 5.847074e-17, 
    5.846928e-17, 5.847174e-17, 5.847389e-17, 5.847669e-17, 5.848174e-17, 
    5.848058e-17, 5.848487e-17, 5.844146e-17, 5.844398e-17, 5.844382e-17, 
    5.844652e-17, 5.84485e-17, 5.845288e-17, 5.845983e-17, 5.845724e-17, 
    5.846208e-17, 5.846303e-17, 5.845571e-17, 5.846014e-17, 5.844572e-17, 
    5.844798e-17, 5.844669e-17, 5.844161e-17, 5.845774e-17, 5.844941e-17, 
    5.846488e-17, 5.846037e-17, 5.847358e-17, 5.846693e-17, 5.847993e-17, 
    5.848533e-17, 5.849074e-17, 5.849671e-17, 5.844544e-17, 5.844371e-17, 
    5.844686e-17, 5.84511e-17, 5.845523e-17, 5.846063e-17, 5.846122e-17, 
    5.846221e-17, 5.846487e-17, 5.846707e-17, 5.846246e-17, 5.846763e-17, 
    5.844836e-17, 5.84585e-17, 5.8443e-17, 5.844756e-17, 5.845088e-17, 
    5.84495e-17, 5.845695e-17, 5.84587e-17, 5.846575e-17, 5.846214e-17, 
    5.848393e-17, 5.847426e-17, 5.85015e-17, 5.849381e-17, 5.844309e-17, 
    5.844547e-17, 5.845362e-17, 5.844975e-17, 5.846103e-17, 5.846378e-17, 
    5.846608e-17, 5.846891e-17, 5.846926e-17, 5.847095e-17, 5.846818e-17, 
    5.847087e-17, 5.846064e-17, 5.846522e-17, 5.845277e-17, 5.845576e-17, 
    5.845441e-17, 5.845288e-17, 5.845759e-17, 5.846251e-17, 5.846273e-17, 
    5.846429e-17, 5.846849e-17, 5.846108e-17, 5.848498e-17, 5.847e-17, 
    5.844804e-17, 5.845246e-17, 5.845323e-17, 5.845149e-17, 5.84635e-17, 
    5.845913e-17, 5.847093e-17, 5.846775e-17, 5.847298e-17, 5.847037e-17, 
    5.846998e-17, 5.846667e-17, 5.846457e-17, 5.845931e-17, 5.845506e-17, 
    5.845176e-17, 5.845253e-17, 5.845617e-17, 5.846284e-17, 5.846925e-17, 
    5.846783e-17, 5.847258e-17, 5.84602e-17, 5.846533e-17, 5.846331e-17, 
    5.84686e-17, 5.845715e-17, 5.846656e-17, 5.84547e-17, 5.845576e-17, 
    5.845904e-17, 5.84656e-17, 5.846722e-17, 5.846875e-17, 5.846783e-17, 
    5.846303e-17, 5.846229e-17, 5.845899e-17, 5.845802e-17, 5.845554e-17, 
    5.845343e-17, 5.845533e-17, 5.84573e-17, 5.846308e-17, 5.846824e-17, 
    5.847391e-17, 5.847534e-17, 5.848172e-17, 5.847638e-17, 5.848504e-17, 
    5.847744e-17, 5.849073e-17, 5.846727e-17, 5.847744e-17, 5.845923e-17, 
    5.846121e-17, 5.846468e-17, 5.84729e-17, 5.846857e-17, 5.847369e-17, 
    5.846227e-17, 5.845624e-17, 5.845482e-17, 5.845194e-17, 5.845488e-17, 
    5.845464e-17, 5.845746e-17, 5.845656e-17, 5.846327e-17, 5.845967e-17, 
    5.846994e-17, 5.847368e-17, 5.848438e-17, 5.849089e-17, 5.849772e-17, 
    5.850069e-17, 5.85016e-17, 5.850198e-17 ;

 MEG_pinene_a =
  4.837514e-17, 4.838066e-17, 4.837961e-17, 4.838402e-17, 4.838161e-17, 
    4.838447e-17, 4.83763e-17, 4.838084e-17, 4.837797e-17, 4.837569e-17, 
    4.839247e-17, 4.838423e-17, 4.840148e-17, 4.839613e-17, 4.840972e-17, 
    4.840058e-17, 4.841158e-17, 4.840955e-17, 4.84159e-17, 4.841409e-17, 
    4.842202e-17, 4.841674e-17, 4.842631e-17, 4.842081e-17, 4.842163e-17, 
    4.841655e-17, 4.838598e-17, 4.839141e-17, 4.838563e-17, 4.838641e-17, 
    4.838608e-17, 4.838162e-17, 4.837931e-17, 4.837478e-17, 4.837562e-17, 
    4.837899e-17, 4.838676e-17, 4.838419e-17, 4.839088e-17, 4.839073e-17, 
    4.839814e-17, 4.83948e-17, 4.840735e-17, 4.84038e-17, 4.841417e-17, 
    4.841154e-17, 4.841403e-17, 4.841329e-17, 4.841404e-17, 4.841019e-17, 
    4.841183e-17, 4.840849e-17, 4.83954e-17, 4.839921e-17, 4.838782e-17, 
    4.838085e-17, 4.837648e-17, 4.837331e-17, 4.837376e-17, 4.837459e-17, 
    4.8379e-17, 4.838325e-17, 4.838646e-17, 4.838859e-17, 4.839071e-17, 
    4.839687e-17, 4.840036e-17, 4.840803e-17, 4.840673e-17, 4.840899e-17, 
    4.841128e-17, 4.841502e-17, 4.841442e-17, 4.841604e-17, 4.8409e-17, 
    4.841365e-17, 4.840596e-17, 4.840805e-17, 4.839095e-17, 4.83849e-17, 
    4.838204e-17, 4.83798e-17, 4.837409e-17, 4.837801e-17, 4.837646e-17, 
    4.838023e-17, 4.838258e-17, 4.838143e-17, 4.838865e-17, 4.838583e-17, 
    4.840056e-17, 4.839421e-17, 4.841102e-17, 4.8407e-17, 4.841199e-17, 
    4.840946e-17, 4.841378e-17, 4.840989e-17, 4.841668e-17, 4.841812e-17, 
    4.841712e-17, 4.842106e-17, 4.840967e-17, 4.841399e-17, 4.838138e-17, 
    4.838157e-17, 4.838247e-17, 4.83785e-17, 4.837827e-17, 4.837474e-17, 
    4.837792e-17, 4.837924e-17, 4.838274e-17, 4.838475e-17, 4.838668e-17, 
    4.839095e-17, 4.839566e-17, 4.840237e-17, 4.840725e-17, 4.841052e-17, 
    4.840854e-17, 4.841029e-17, 4.840832e-17, 4.840742e-17, 4.841755e-17, 
    4.841183e-17, 4.842049e-17, 4.842002e-17, 4.841607e-17, 4.842007e-17, 
    4.83817e-17, 4.838063e-17, 4.837678e-17, 4.837979e-17, 4.837436e-17, 
    4.837736e-17, 4.837906e-17, 4.838581e-17, 4.838738e-17, 4.838873e-17, 
    4.839148e-17, 4.839497e-17, 4.840108e-17, 4.840646e-17, 4.841143e-17, 
    4.841107e-17, 4.84112e-17, 4.841227e-17, 4.840956e-17, 4.841272e-17, 
    4.841322e-17, 4.841187e-17, 4.841996e-17, 4.841765e-17, 4.842001e-17, 
    4.841851e-17, 4.838098e-17, 4.838281e-17, 4.838182e-17, 4.838367e-17, 
    4.838234e-17, 4.838816e-17, 4.838991e-17, 4.83982e-17, 4.839488e-17, 
    4.840026e-17, 4.839545e-17, 4.839628e-17, 4.840029e-17, 4.839573e-17, 
    4.84061e-17, 4.839894e-17, 4.841232e-17, 4.840501e-17, 4.841277e-17, 
    4.841141e-17, 4.841369e-17, 4.84157e-17, 4.841829e-17, 4.842298e-17, 
    4.842191e-17, 4.842589e-17, 4.838557e-17, 4.838792e-17, 4.838777e-17, 
    4.839027e-17, 4.839211e-17, 4.839618e-17, 4.840264e-17, 4.840022e-17, 
    4.840473e-17, 4.840561e-17, 4.839881e-17, 4.840292e-17, 4.838954e-17, 
    4.839163e-17, 4.839043e-17, 4.838572e-17, 4.840069e-17, 4.839296e-17, 
    4.840732e-17, 4.840313e-17, 4.84154e-17, 4.840923e-17, 4.84213e-17, 
    4.842632e-17, 4.843135e-17, 4.843689e-17, 4.838927e-17, 4.838766e-17, 
    4.839059e-17, 4.839452e-17, 4.839836e-17, 4.840338e-17, 4.840393e-17, 
    4.840485e-17, 4.840731e-17, 4.840936e-17, 4.840508e-17, 4.840988e-17, 
    4.839198e-17, 4.84014e-17, 4.8387e-17, 4.839124e-17, 4.839432e-17, 
    4.839303e-17, 4.839997e-17, 4.840158e-17, 4.840813e-17, 4.840478e-17, 
    4.842502e-17, 4.841603e-17, 4.844134e-17, 4.843419e-17, 4.838709e-17, 
    4.838929e-17, 4.839687e-17, 4.839327e-17, 4.840374e-17, 4.84063e-17, 
    4.840844e-17, 4.841107e-17, 4.84114e-17, 4.841297e-17, 4.841039e-17, 
    4.841289e-17, 4.840339e-17, 4.840764e-17, 4.839608e-17, 4.839885e-17, 
    4.83976e-17, 4.839618e-17, 4.840055e-17, 4.840513e-17, 4.840533e-17, 
    4.840678e-17, 4.841068e-17, 4.840379e-17, 4.8426e-17, 4.841208e-17, 
    4.839169e-17, 4.839579e-17, 4.83965e-17, 4.839489e-17, 4.840604e-17, 
    4.840198e-17, 4.841294e-17, 4.840999e-17, 4.841485e-17, 4.841243e-17, 
    4.841207e-17, 4.840898e-17, 4.840704e-17, 4.840215e-17, 4.839821e-17, 
    4.839514e-17, 4.839586e-17, 4.839923e-17, 4.840543e-17, 4.841138e-17, 
    4.841006e-17, 4.841448e-17, 4.840298e-17, 4.840774e-17, 4.840587e-17, 
    4.841078e-17, 4.840014e-17, 4.840889e-17, 4.839787e-17, 4.839886e-17, 
    4.84019e-17, 4.8408e-17, 4.84095e-17, 4.841092e-17, 4.841007e-17, 
    4.840561e-17, 4.840493e-17, 4.840185e-17, 4.840095e-17, 4.839865e-17, 
    4.83967e-17, 4.839845e-17, 4.840028e-17, 4.840565e-17, 4.841044e-17, 
    4.841571e-17, 4.841705e-17, 4.842296e-17, 4.8418e-17, 4.842605e-17, 
    4.841899e-17, 4.843134e-17, 4.840955e-17, 4.841899e-17, 4.840208e-17, 
    4.840392e-17, 4.840714e-17, 4.841477e-17, 4.841076e-17, 4.84155e-17, 
    4.840491e-17, 4.83993e-17, 4.839798e-17, 4.839531e-17, 4.839804e-17, 
    4.839782e-17, 4.840043e-17, 4.83996e-17, 4.840583e-17, 4.840249e-17, 
    4.841203e-17, 4.841549e-17, 4.842544e-17, 4.843149e-17, 4.843783e-17, 
    4.844059e-17, 4.844143e-17, 4.844178e-17 ;

 MEG_thujene_a =
  1.220108e-18, 1.220242e-18, 1.220217e-18, 1.220324e-18, 1.220265e-18, 
    1.220335e-18, 1.220136e-18, 1.220247e-18, 1.220177e-18, 1.220121e-18, 
    1.220529e-18, 1.220329e-18, 1.220748e-18, 1.220618e-18, 1.220949e-18, 
    1.220727e-18, 1.220994e-18, 1.220945e-18, 1.221099e-18, 1.221055e-18, 
    1.221248e-18, 1.22112e-18, 1.221352e-18, 1.221219e-18, 1.221238e-18, 
    1.221115e-18, 1.220372e-18, 1.220504e-18, 1.220363e-18, 1.220382e-18, 
    1.220374e-18, 1.220266e-18, 1.220209e-18, 1.220099e-18, 1.22012e-18, 
    1.220202e-18, 1.220391e-18, 1.220328e-18, 1.220491e-18, 1.220487e-18, 
    1.220667e-18, 1.220586e-18, 1.220891e-18, 1.220805e-18, 1.221057e-18, 
    1.220993e-18, 1.221054e-18, 1.221036e-18, 1.221054e-18, 1.22096e-18, 
    1.221e-18, 1.220919e-18, 1.220601e-18, 1.220693e-18, 1.220416e-18, 
    1.220247e-18, 1.220141e-18, 1.220063e-18, 1.220074e-18, 1.220095e-18, 
    1.220202e-18, 1.220305e-18, 1.220383e-18, 1.220435e-18, 1.220487e-18, 
    1.220637e-18, 1.220721e-18, 1.220908e-18, 1.220876e-18, 1.220931e-18, 
    1.220987e-18, 1.221078e-18, 1.221063e-18, 1.221103e-18, 1.220931e-18, 
    1.221044e-18, 1.220858e-18, 1.220908e-18, 1.220492e-18, 1.220345e-18, 
    1.220276e-18, 1.220221e-18, 1.220083e-18, 1.220178e-18, 1.22014e-18, 
    1.220232e-18, 1.220289e-18, 1.220261e-18, 1.220437e-18, 1.220368e-18, 
    1.220726e-18, 1.220572e-18, 1.22098e-18, 1.220883e-18, 1.221004e-18, 
    1.220943e-18, 1.221047e-18, 1.220953e-18, 1.221118e-18, 1.221153e-18, 
    1.221129e-18, 1.221224e-18, 1.220948e-18, 1.221053e-18, 1.22026e-18, 
    1.220264e-18, 1.220286e-18, 1.22019e-18, 1.220184e-18, 1.220098e-18, 
    1.220176e-18, 1.220208e-18, 1.220293e-18, 1.220342e-18, 1.220389e-18, 
    1.220492e-18, 1.220607e-18, 1.22077e-18, 1.220889e-18, 1.220968e-18, 
    1.22092e-18, 1.220963e-18, 1.220915e-18, 1.220893e-18, 1.221139e-18, 
    1.221e-18, 1.221211e-18, 1.221199e-18, 1.221103e-18, 1.221201e-18, 
    1.220268e-18, 1.220241e-18, 1.220148e-18, 1.220221e-18, 1.220089e-18, 
    1.220162e-18, 1.220203e-18, 1.220368e-18, 1.220406e-18, 1.220439e-18, 
    1.220505e-18, 1.22059e-18, 1.220739e-18, 1.22087e-18, 1.22099e-18, 
    1.220982e-18, 1.220985e-18, 1.221011e-18, 1.220945e-18, 1.221022e-18, 
    1.221034e-18, 1.221001e-18, 1.221198e-18, 1.221142e-18, 1.221199e-18, 
    1.221163e-18, 1.22025e-18, 1.220295e-18, 1.22027e-18, 1.220315e-18, 
    1.220283e-18, 1.220425e-18, 1.220467e-18, 1.220669e-18, 1.220588e-18, 
    1.220719e-18, 1.220602e-18, 1.220622e-18, 1.22072e-18, 1.220609e-18, 
    1.220861e-18, 1.220687e-18, 1.221012e-18, 1.220834e-18, 1.221023e-18, 
    1.22099e-18, 1.221045e-18, 1.221094e-18, 1.221157e-18, 1.221271e-18, 
    1.221245e-18, 1.221342e-18, 1.220362e-18, 1.220419e-18, 1.220415e-18, 
    1.220476e-18, 1.220521e-18, 1.22062e-18, 1.220777e-18, 1.220718e-18, 
    1.220827e-18, 1.220849e-18, 1.220684e-18, 1.220784e-18, 1.220458e-18, 
    1.220509e-18, 1.22048e-18, 1.220365e-18, 1.220729e-18, 1.220541e-18, 
    1.220891e-18, 1.220789e-18, 1.221087e-18, 1.220937e-18, 1.22123e-18, 
    1.221352e-18, 1.221475e-18, 1.22161e-18, 1.220452e-18, 1.220413e-18, 
    1.220484e-18, 1.220579e-18, 1.220673e-18, 1.220795e-18, 1.220808e-18, 
    1.22083e-18, 1.22089e-18, 1.22094e-18, 1.220836e-18, 1.220953e-18, 
    1.220518e-18, 1.220747e-18, 1.220396e-18, 1.2205e-18, 1.220574e-18, 
    1.220543e-18, 1.220712e-18, 1.220751e-18, 1.22091e-18, 1.220829e-18, 
    1.221321e-18, 1.221102e-18, 1.221718e-18, 1.221544e-18, 1.220399e-18, 
    1.220452e-18, 1.220636e-18, 1.220549e-18, 1.220804e-18, 1.220866e-18, 
    1.220918e-18, 1.220982e-18, 1.22099e-18, 1.221028e-18, 1.220965e-18, 
    1.221026e-18, 1.220795e-18, 1.220898e-18, 1.220617e-18, 1.220684e-18, 
    1.220654e-18, 1.22062e-18, 1.220726e-18, 1.220837e-18, 1.220842e-18, 
    1.220877e-18, 1.220972e-18, 1.220805e-18, 1.221345e-18, 1.221006e-18, 
    1.22051e-18, 1.22061e-18, 1.220628e-18, 1.220588e-18, 1.220859e-18, 
    1.220761e-18, 1.221027e-18, 1.220956e-18, 1.221074e-18, 1.221015e-18, 
    1.221006e-18, 1.220931e-18, 1.220884e-18, 1.220765e-18, 1.220669e-18, 
    1.220594e-18, 1.220612e-18, 1.220694e-18, 1.220845e-18, 1.220989e-18, 
    1.220957e-18, 1.221065e-18, 1.220785e-18, 1.220901e-18, 1.220855e-18, 
    1.220975e-18, 1.220716e-18, 1.220929e-18, 1.220661e-18, 1.220685e-18, 
    1.220759e-18, 1.220907e-18, 1.220944e-18, 1.220978e-18, 1.220957e-18, 
    1.220849e-18, 1.220832e-18, 1.220758e-18, 1.220736e-18, 1.22068e-18, 
    1.220632e-18, 1.220675e-18, 1.220719e-18, 1.22085e-18, 1.220966e-18, 
    1.221095e-18, 1.221127e-18, 1.221271e-18, 1.22115e-18, 1.221346e-18, 
    1.221174e-18, 1.221474e-18, 1.220945e-18, 1.221174e-18, 1.220763e-18, 
    1.220808e-18, 1.220886e-18, 1.221072e-18, 1.220974e-18, 1.22109e-18, 
    1.220832e-18, 1.220695e-18, 1.220663e-18, 1.220598e-18, 1.220665e-18, 
    1.220659e-18, 1.220723e-18, 1.220703e-18, 1.220854e-18, 1.220773e-18, 
    1.221005e-18, 1.221089e-18, 1.221331e-18, 1.221478e-18, 1.221632e-18, 
    1.221699e-18, 1.22172e-18, 1.221728e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  1.263632e-25, 1.400983e-25, -4.944636e-26, -4.477649e-25, 1.620745e-25, 
    6.86757e-26, 2.307502e-25, -9.065174e-26, 3.076668e-25, 1.593275e-25, 
    2.554734e-25, 1.236162e-25, 2.774496e-25, 2.582204e-25, -7.691661e-26, 
    -1.648207e-26, -3.40631e-25, -3.021727e-25, -3.873304e-25, 1.840507e-25, 
    -3.351369e-25, -2.197612e-26, 6.098396e-25, -1.043869e-25, -5.768744e-26, 
    3.955716e-25, -5.411638e-25, -1.648214e-25, 1.703156e-25, 1.373513e-25, 
    -2.087738e-25, 2.032799e-25, 8.790487e-26, -4.450179e-25, -3.43378e-25, 
    -1.648214e-25, 6.043463e-26, 6.318165e-26, 1.428454e-25, -6.043454e-25, 
    9.339892e-26, 2.032799e-25, 8.790487e-26, -5.219339e-26, -2.28003e-25, 
    2.472331e-26, 2.582204e-25, -3.46125e-25, 5.603931e-25, -2.33497e-25, 
    -4.120529e-26, -3.516191e-25, -5.768744e-26, -1.428452e-25, 
    -2.527262e-25, 5.768753e-25, -8.240992e-27, 2.582204e-25, 2.14268e-25, 
    -3.873304e-25, 1.483394e-25, -1.318571e-25, -2.115208e-25, 2.774496e-25, 
    2.362442e-25, 6.56539e-25, 6.86757e-26, -2.582203e-25, -2.3075e-25, 
    -2.801964e-25, -3.214018e-25, 4.395248e-26, -6.867554e-26, -1.895446e-25, 
    -4.807293e-25, 4.66995e-26, 1.510864e-25, -3.571131e-25, 2.801966e-25, 
    -2.389911e-25, 1.483394e-25, -3.186548e-25, 1.181221e-25, -5.906102e-25, 
    1.510864e-25, 4.148008e-25, 2.774496e-25, 2.747033e-26, -3.488721e-25, 
    2.225091e-25, -3.818364e-25, -1.126279e-25, 5.219355e-26, 1.840507e-25, 
    -2.609673e-25, 2.692085e-25, 7.96638e-26, -9.339876e-26, -4.615001e-25, 
    -2.692083e-25, -2.527262e-25, -6.043446e-26, -4.669934e-26, 1.126281e-25, 
    1.758097e-25, 3.763425e-25, 3.378841e-25, 2.060269e-25, -2.25256e-25, 
    -3.626072e-25, -4.038125e-25, 1.648223e-26, 1.455924e-25, -4.917174e-25, 
    -2.884375e-25, 1.840507e-25, -2.966786e-25, -1.18122e-25, 1.428454e-25, 
    2.719555e-25, -2.170149e-25, -3.37884e-25, -1.016398e-25, -4.395231e-26, 
    3.076668e-25, 1.730626e-25, -6.043446e-26, -3.351369e-25, -2.25256e-25, 
    -4.56006e-25, -2.142679e-25, 2.444853e-25, -1.291101e-25, -4.669934e-26, 
    -5.493967e-27, 5.494132e-27, 7.96638e-26, 1.813037e-25, 8.790487e-26, 
    1.977859e-25, -2.3075e-25, -2.801964e-25, -6.263216e-25, -6.455508e-25, 
    1.813037e-25, -7.142256e-26, 7.96638e-26, 1.04387e-25, -2.911845e-25, 
    -4.422709e-25, -1.950387e-25, -5.933573e-25, -1.20869e-25, 2.609674e-25, 
    3.598603e-25, 3.516192e-25, 1.840507e-25, 1.181221e-25, 4.944653e-26, 
    -4.148007e-25, -9.614578e-26, -1.263631e-25, -4.038125e-25, -2.28003e-25, 
    -2.582203e-25, -3.159078e-25, 1.730626e-25, 6.592867e-26, -4.779822e-25, 
    1.758097e-25, -1.291101e-25, -1.648214e-25, 2.14268e-25, 9.889298e-26, 
    2.307502e-25, -1.400982e-25, 2.280031e-25, -2.005327e-25, -1.483393e-25, 
    -1.126279e-25, -2.472314e-26, 8.257385e-32, -4.065596e-25, 1.0164e-25, 
    -1.648207e-26, -1.043869e-25, -4.340298e-25, -2.747024e-25, 2.747026e-25, 
    2.747033e-26, -1.922916e-25, 2.747033e-26, -7.416958e-26, -1.922916e-25, 
    1.730626e-25, 2.472331e-26, -1.675684e-25, -8.515768e-26, 5.219355e-26, 
    -4.120536e-25, -5.356697e-25, -2.582203e-25, -1.922909e-26, 
    -1.922916e-25, 1.208692e-25, 3.021728e-25, -6.208275e-25, -4.50512e-25, 
    -3.571131e-25, -4.340298e-25, -9.889281e-26, 6.043463e-26, 3.406311e-25, 
    4.395248e-26, -3.186548e-25, -2.884375e-25, 6.318165e-26, -5.768744e-26, 
    -2.582203e-25, -3.049197e-25, -2.801964e-25, -1.538333e-25, 
    -2.801964e-25, 3.131609e-25, 1.181221e-25, -5.494041e-26, -1.922916e-25, 
    3.21402e-25, -1.455922e-25, -6.592851e-26, 2.252561e-25, 2.252561e-25, 
    2.252561e-25, 5.274289e-25, 8.257613e-32, 1.04387e-25, -2.664613e-25, 
    3.57114e-26, 1.373521e-26, 1.318573e-25, -8.790471e-26, 4.999586e-25, 
    1.675686e-25, -2.856905e-25, -1.428452e-25, -1.730625e-25, -1.373512e-25, 
    5.054526e-25, -1.922916e-25, 2.472323e-25, 7.416975e-26, -1.648214e-25, 
    -3.43378e-25, 4.230419e-25, 5.988515e-25, -2.25256e-25, -3.296421e-26, 
    -2.966786e-25, -4.642471e-25, 1.291103e-25, 1.346043e-25, -2.3075e-25, 
    5.494058e-26, -5.60393e-25, 8.257501e-32, 5.136937e-25, -6.620329e-25, 
    -2.554732e-25, -1.895446e-25, -7.416958e-26, -8.240992e-27, 
    -4.120529e-26, 1.648216e-25, -1.730625e-25, -3.268959e-25, 8.241157e-27, 
    -1.098809e-25, -3.763423e-25, -5.219339e-26, -1.483393e-25, 
    -9.339876e-26, 2.966788e-25, -3.571131e-25, -1.648207e-26, -2.142679e-25, 
    -1.648214e-25, 2.801966e-25, 1.758097e-25, 4.230419e-25, -2.115208e-25, 
    4.944653e-26, -3.296429e-25, 2.280031e-25, -1.318571e-25, -9.065174e-26, 
    -1.895446e-25, -3.186548e-25, -1.126279e-25, 4.120545e-26, 4.615002e-25, 
    3.461252e-25, 3.516192e-25, -2.582203e-25, 8.515785e-26, 3.131609e-25, 
    -1.455922e-25, 5.027056e-25, 2.307502e-25, 1.867978e-25, 1.04387e-25, 
    4.66995e-26, 3.021735e-26, -1.538333e-25, -6.043446e-26, 1.04387e-25, 
    2.197628e-26, -3.873304e-25, 3.18655e-25, -2.417381e-25, 2.280031e-25, 
    4.36777e-25, -2.856905e-25, -2.36244e-25, -2.719554e-25, -2.197612e-26, 
    1.977859e-25, 3.021735e-26, -3.296421e-26, 4.66995e-26, -2.197612e-26, 
    4.120538e-25, 1.0164e-25, -4.862233e-25, 7.691677e-26, -5.768744e-26, 
    -1.922916e-25, -9.889281e-26, -2.472314e-26 ;

 M_LITR2C_TO_LEACHING =
  1.291102e-25, -2.746971e-27, -7.142259e-26, 1.181221e-25, 3.571138e-26, 
    -9.889284e-26, -2.197614e-26, -2.197614e-26, 1.593275e-25, -1.483393e-25, 
    1.593275e-25, -1.703155e-25, -2.362441e-25, -1.758095e-25, -2.28003e-25, 
    -2.746971e-27, -3.735953e-25, -4.202947e-25, 1.098815e-26, -4.669937e-26, 
    -1.510863e-25, 1.922918e-25, 4.395245e-26, -3.021722e-26, 6.592865e-26, 
    -1.263631e-25, 1.565805e-25, 1.758096e-25, -1.428452e-25, 4.038127e-25, 
    4.395245e-26, -3.543661e-25, -1.593274e-25, -4.944639e-26, 5.768757e-26, 
    -1.538333e-25, 6.318163e-26, -3.131608e-25, 1.373513e-25, 9.339889e-26, 
    -2.74702e-26, 7.14227e-26, 1.263632e-25, -1.593274e-25, -1.098809e-25, 
    1.153751e-25, 5.494055e-26, -1.20869e-25, -2.74702e-26, 8.24108e-26, 
    -1.291101e-25, -1.263631e-25, -3.241489e-25, -2.225089e-25, 1.483394e-25, 
    3.021733e-26, -1.483393e-25, 3.021733e-26, 1.373518e-26, -1.098805e-26, 
    -2.472317e-26, 2.472323e-25, -1.538333e-25, 2.005329e-25, 5.494103e-27, 
    8.515782e-26, -9.889284e-26, 1.867977e-25, 1.950388e-25, 2.719555e-25, 
    2.060269e-25, -1.675685e-25, -1.648209e-26, -2.472317e-26, -1.236161e-25, 
    5.494055e-26, 2.74703e-26, -1.895447e-25, -1.043869e-25, 4.669947e-26, 
    -5.054525e-25, 1.0164e-25, -8.515771e-26, -3.845834e-25, 4.395245e-26, 
    1.483394e-25, 1.565805e-25, 5.219352e-26, 2.829436e-25, -5.768747e-26, 
    -3.571127e-26, -3.845829e-26, 1.703156e-25, -1.15375e-25, -3.296424e-26, 
    -2.994256e-25, 5.494103e-27, -4.120532e-26, -1.043869e-25, -4.395234e-26, 
    1.648215e-25, -1.016399e-25, -2.362441e-25, -3.845829e-26, -1.263631e-25, 
    1.346043e-25, -2.499792e-25, -1.373512e-25, -3.571127e-26, -2.197614e-26, 
    1.428453e-25, -6.867557e-26, -8.790474e-26, -1.675685e-25, -2.444852e-25, 
    9.889295e-26, 1.538334e-25, 1.64822e-26, -2.197614e-26, 1.565805e-25, 
    -1.346042e-25, -2.142679e-25, 5.494103e-27, 1.09881e-25, 2.774496e-25, 
    1.428453e-25, 4.94465e-26, -9.889284e-26, -3.296429e-25, 7.14227e-26, 
    8.790485e-26, -7.416961e-26, 4.669947e-26, 3.021733e-26, -1.291101e-25, 
    6.592865e-26, -2.472322e-25, -2.389911e-25, 1.922923e-26, -1.922912e-26, 
    -1.977857e-25, -2.197614e-26, -1.620744e-25, -8.790474e-26, 1.126281e-25, 
    1.153751e-25, -9.614581e-26, -2.472317e-26, -2.911846e-25, 3.076668e-25, 
    1.318572e-25, -1.428452e-25, -1.703155e-25, 5.494103e-27, 2.609674e-25, 
    -1.648209e-26, -2.197614e-26, -1.373512e-25, -2.884375e-25, 1.400983e-25, 
    -2.472322e-25, 5.494055e-26, -1.016399e-25, 1.64822e-26, 2.197625e-26, 
    9.065187e-26, -5.494044e-26, -1.922912e-26, -6.043449e-26, 9.065187e-26, 
    -1.730625e-25, -2.472322e-25, 2.197625e-26, -2.417381e-25, 1.126281e-25, 
    6.318163e-26, 4.395245e-26, -2.692084e-25, 3.021733e-26, 8.790485e-26, 
    -2.170149e-25, 9.339889e-26, -3.021722e-26, 9.889295e-26, -1.538333e-25, 
    9.065187e-26, 6.592865e-26, 9.339889e-26, 2.389912e-25, 1.07134e-25, 
    5.351444e-32, -2.060268e-25, -1.648209e-26, -1.593274e-25, -3.241489e-25, 
    -4.065596e-25, -7.691664e-26, 1.703156e-25, 2.19762e-25, 7.966377e-26, 
    -4.395234e-26, 7.691675e-26, -1.373512e-25, -2.74702e-26, 4.395245e-26, 
    3.84584e-26, 2.472323e-25, 1.538334e-25, 3.571138e-26, 1.236162e-25, 
    5.351459e-32, -4.120532e-26, -8.790474e-26, 1.09881e-25, -1.043869e-25, 
    8.790485e-26, -1.15375e-25, -4.395234e-26, -2.417381e-25, -1.730625e-25, 
    4.120543e-26, 6.04346e-26, 6.592865e-26, 1.263632e-25, -2.856905e-25, 
    -3.845829e-26, 7.691675e-26, -1.922917e-25, 9.339889e-26, 1.373513e-25, 
    -6.592854e-26, 2.032799e-25, 3.571138e-26, 1.648215e-25, 2.472328e-26, 
    1.703156e-25, -7.142259e-26, -1.428452e-25, 1.181221e-25, -1.455923e-25, 
    -4.120532e-26, -2.28003e-25, 3.845835e-25, -2.637143e-25, -1.373512e-25, 
    -9.065177e-26, 2.74703e-26, -3.845829e-26, -3.021727e-25, -5.494044e-26, 
    -1.18122e-25, 3.021728e-25, 2.472328e-26, 2.747078e-27, -1.043869e-25, 
    1.318572e-25, 8.241128e-27, -1.236161e-25, -1.730625e-25, -6.318152e-26, 
    -4.47765e-25, -3.296424e-26, -2.197614e-26, -2.197619e-25, -5.768747e-26, 
    9.339889e-26, 1.483394e-25, -2.197619e-25, -1.813036e-25, 1.64822e-26, 
    -2.142679e-25, 6.04346e-26, -7.691664e-26, -2.74702e-26, -5.768747e-26, 
    -2.115208e-25, -2.746971e-27, 8.790485e-26, -1.291101e-25, -1.620744e-25, 
    7.14227e-26, -8.241069e-26, -1.428452e-25, -5.768747e-26, -1.016399e-25, 
    5.494055e-26, 7.14227e-26, 8.790485e-26, -2.74702e-26, -1.346042e-25, 
    -2.444852e-25, 3.159079e-25, 1.098815e-26, -9.065177e-26, -2.362441e-25, 
    2.74703e-26, -2.499792e-25, 1.04387e-25, -2.582203e-25, 9.614592e-26, 
    -8.241021e-27, -1.15375e-25, -1.098805e-26, -4.395239e-25, 1.428453e-25, 
    4.120543e-26, 3.873306e-25, -2.692084e-25, -2.087738e-25, 3.021733e-26, 
    5.219352e-26, -1.675685e-25, -1.428452e-25, 7.691675e-26, -6.318152e-26, 
    2.14268e-25, 4.120543e-26, -1.20869e-25, 9.339889e-26, -2.472317e-26, 
    -2.197619e-25, -3.021722e-26, -3.296424e-26, 3.84584e-26, 1.263632e-25, 
    4.94465e-26, -3.296424e-26, -8.515771e-26, -7.966367e-26, -1.565804e-25, 
    7.691675e-26, 2.939317e-25, 7.14227e-26, -2.829435e-25, 1.126281e-25, 
    -1.236161e-25, 1.373513e-25, -1.15375e-25 ;

 M_LITR3C_TO_LEACHING =
  -9.065179e-26, -8.10372e-26, -4.257886e-26, 8.653131e-26, 5.494076e-27, 
    -3.983183e-26, -7.691667e-26, -1.071339e-25, 1.263632e-25, -1.703155e-25, 
    1.373539e-27, -4.669939e-26, 1.785569e-26, -9.20253e-26, 5.768755e-26, 
    -2.47232e-26, -3.296427e-26, 8.241077e-26, -7.416964e-26, -5.219344e-26, 
    -3.021725e-26, 4.257891e-26, -3.021725e-26, 3.708486e-26, -9.614584e-26, 
    8.653131e-26, -9.889287e-26, -1.263631e-25, -4.257886e-26, -1.09881e-25, 
    -7.691667e-26, 4.669945e-26, 2.675734e-32, 1.140016e-25, 7.279618e-26, 
    -3.433778e-26, -8.790477e-26, 3.845837e-26, 8.378428e-26, -8.653126e-26, 
    -7.00491e-26, -9.889287e-26, 2.747028e-26, 2.747028e-26, -7.279613e-26, 
    -3.57113e-26, -1.071339e-25, 2.472325e-26, 1.648217e-26, -1.579539e-25, 
    9.339887e-26, 2.747028e-26, -1.208691e-25, 1.785569e-26, 1.92292e-26, 
    1.92292e-26, 9.614614e-27, -1.249896e-25, 4.807296e-26, 1.304837e-25, 
    -1.098807e-26, 8.790482e-26, -1.648215e-25, -1.167485e-25, 1.510866e-26, 
    -7.966369e-26, 2.609676e-26, -1.400982e-25, 1.181221e-25, -2.746998e-27, 
    6.867565e-26, -5.631398e-26, 5.21935e-26, -3.708481e-26, 1.291102e-25, 
    -5.906101e-26, -3.296427e-26, 5.768755e-26, -1.785563e-26, -3.296427e-26, 
    -1.043869e-25, -4.257886e-26, -8.241071e-26, 8.653131e-26, 7.966375e-26, 
    -1.373486e-27, 3.571135e-26, 9.477238e-26, 9.889292e-26, -5.219344e-26, 
    -4.669939e-26, 8.515779e-26, 8.790482e-26, -5.494023e-27, -1.510861e-26, 
    -9.614584e-26, 5.21935e-26, -7.142262e-26, -8.241047e-27, -1.648212e-26, 
    -1.318572e-25, -3.845832e-26, -3.159076e-26, -3.021725e-26, 3.845837e-26, 
    -9.065179e-26, 9.75194e-26, 6.867589e-27, -2.746998e-27, -7.829018e-26, 
    1.002664e-25, 9.614614e-27, 6.31816e-26, -4.669939e-26, 4.807296e-26, 
    -6.592857e-26, -5.631398e-26, -8.241071e-26, 1.826772e-25, -1.12628e-25, 
    6.867565e-26, 1.12628e-25, -8.790477e-26, 5.494052e-26, -1.071339e-25, 
    5.081998e-26, 3.02173e-26, 4.944647e-26, 4.120564e-27, -7.142262e-26, 
    -1.455923e-25, 3.845837e-26, -1.37351e-26, -2.334968e-26, 3.02173e-26, 
    6.180808e-26, 3.571135e-26, 1.12628e-25, -6.318154e-26, -6.318154e-26, 
    -3.845832e-26, -1.552069e-25, 7.416969e-26, 3.571135e-26, -7.416964e-26, 
    -8.241047e-27, 5.494076e-27, -1.66195e-25, 4.532594e-26, -1.922915e-26, 
    9.889292e-26, 3.571135e-26, -7.691667e-26, -1.648212e-26, -9.614584e-26, 
    8.653131e-26, 5.494076e-27, 1.030135e-25, -1.428453e-25, -8.241047e-27, 
    6.730214e-26, 1.785569e-26, -1.098807e-26, -3.57113e-26, 1.648217e-26, 
    -1.140015e-25, -8.241047e-27, 2.675725e-32, 4.120564e-27, 1.510866e-26, 
    -1.785563e-26, 3.02173e-26, -4.120511e-27, -1.346042e-25, -5.494047e-26, 
    -9.889287e-26, 1.387248e-25, 3.845837e-26, 4.395242e-26, -8.790477e-26, 
    1.098813e-26, 5.768755e-26, 1.346042e-25, 2.747052e-27, 1.09881e-25, 
    2.060271e-26, 1.455923e-25, -2.609671e-26, -1.442188e-25, 1.07134e-25, 
    8.241101e-27, -1.359777e-25, 5.081998e-26, -1.37351e-26, 2.197622e-26, 
    5.768755e-26, 6.592862e-26, -4.120535e-26, 3.708486e-26, -1.373512e-25, 
    2.197622e-26, -1.346042e-25, -4.532588e-26, 6.043457e-26, 2.032799e-25, 
    5.081998e-26, -1.236158e-26, 1.785569e-26, 9.065185e-26, 6.180808e-26, 
    -1.703155e-25, -8.241047e-27, 2.747028e-26, -2.197617e-26, -3.708481e-26, 
    2.472323e-25, 1.483394e-25, 9.614614e-27, 5.768755e-26, -9.889287e-26, 
    -3.845832e-26, -4.120535e-26, 1.648217e-26, -3.296427e-26, -2.746998e-27, 
    -8.241047e-27, -1.291101e-25, 2.884379e-26, -1.09881e-25, -1.414718e-25, 
    1.249896e-25, -7.142262e-26, 4.120564e-27, -7.691667e-26, -5.631398e-26, 
    3.296432e-26, -1.140015e-25, -1.043869e-25, -3.708481e-26, 4.944647e-26, 
    7.279618e-26, -1.291101e-25, -3.021725e-26, 2.675717e-32, -1.758096e-25, 
    7.966375e-26, 1.964123e-25, -1.236158e-26, -8.241047e-27, 3.02173e-26, 
    -4.120535e-26, 3.571135e-26, 6.592862e-26, -1.140015e-25, 1.359778e-25, 
    1.373515e-26, -8.241071e-26, -7.142262e-26, -8.927828e-26, -1.208691e-25, 
    -1.648212e-26, -7.00491e-26, -2.197617e-26, -1.140015e-25, 7.416969e-26, 
    -9.751935e-26, 5.494076e-27, -1.112545e-25, 4.120564e-27, -2.334968e-26, 
    4.669945e-26, 3.708486e-26, -5.494023e-27, -4.807291e-26, -7.554316e-26, 
    -4.395237e-26, 2.675726e-32, -1.37351e-26, -6.043452e-26, 1.04387e-25, 
    -4.669939e-26, 5.356701e-26, -1.840506e-25, -2.197617e-26, -7.691667e-26, 
    -6.592857e-26, -8.241071e-26, -3.296427e-26, -3.845832e-26, 
    -5.906101e-26, 9.477238e-26, 8.241101e-27, -1.771831e-25, 1.620745e-25, 
    1.236164e-26, 1.620745e-25, -5.768749e-26, -6.592857e-26, -9.889287e-26, 
    2.675724e-32, 8.103726e-26, -8.241047e-27, -1.785563e-26, -1.263631e-25, 
    -9.61456e-27, -1.867977e-25, -4.807291e-26, -1.318572e-25, -3.845832e-26, 
    -4.257886e-26, 6.592862e-26, 1.648217e-26, -8.10372e-26, -4.395237e-26, 
    2.884379e-26, 3.983189e-26, -1.922917e-25, -8.515774e-26, -1.112545e-25, 
    -1.400982e-25, -6.730208e-26, 1.400983e-25, -3.57113e-26, 9.614614e-27, 
    4.532594e-26, -7.416964e-26, -6.043452e-26, -7.279613e-26, 4.12054e-26, 
    9.614614e-27, -5.631398e-26, -8.241047e-27, 5.494076e-27, 6.31816e-26, 
    -1.373486e-27, 9.339887e-26, -3.845832e-26, -4.257886e-26 ;

 M_SOIL1C_TO_LEACHING =
  -2.335273e-20, -8.89189e-21, -8.658897e-21, -2.121358e-20, 5.966474e-21, 
    -4.248867e-21, 1.461406e-20, -1.799809e-20, -1.348343e-20, -1.527764e-20, 
    -4.440565e-21, -1.858273e-20, 2.433378e-20, 6.935087e-21, -2.247284e-20, 
    -3.593788e-21, 1.04848e-20, -3.492013e-21, 4.357335e-20, 4.176895e-20, 
    2.112169e-20, -8.833353e-21, 1.766306e-20, 3.885032e-20, -3.692238e-20, 
    -1.653919e-20, -3.702389e-20, 2.645654e-20, -4.432398e-20, 2.353706e-20, 
    2.491848e-20, 1.985702e-20, -7.205669e-21, 9.802308e-22, 2.272023e-20, 
    4.974563e-23, -1.875691e-20, 1.085942e-21, 2.945799e-20, 3.391129e-20, 
    -2.431372e-20, 7.684063e-21, -1.588721e-20, -3.108793e-20, -8.83901e-21, 
    -3.907879e-20, -2.95762e-20, -9.559437e-21, -1.218174e-20, -1.306076e-20, 
    3.065789e-20, -2.769206e-20, -1.907026e-21, 3.797584e-20, -7.217547e-21, 
    -2.956524e-21, 4.56383e-21, -3.229322e-20, 1.753046e-20, 6.306894e-21, 
    2.29651e-20, 5.437563e-20, -1.128604e-20, -1.221341e-20, -1.00542e-20, 
    2.189748e-21, -8.44065e-21, -2.613393e-20, 3.803301e-21, -6.128754e-21, 
    1.701786e-20, 1.467034e-20, -1.301986e-21, -2.196846e-20, -1.465649e-20, 
    -2.319327e-20, -9.370842e-21, 3.808891e-20, -2.890132e-20, 1.456092e-20, 
    -2.771897e-21, 1.027585e-20, 4.4972e-20, 9.553217e-21, 9.236253e-21, 
    -3.176199e-21, -2.309044e-21, 1.079918e-20, -1.851378e-20, -2.271854e-20, 
    1.340794e-20, 2.153194e-20, 7.932299e-21, -2.667254e-20, 5.667064e-21, 
    9.620767e-21, -1.051701e-20, -4.910074e-20, 7.325822e-21, 3.218211e-20, 
    2.359642e-20, -9.066901e-21, -1.713433e-20, 4.921206e-21, 1.192275e-21, 
    1.347636e-20, 3.00424e-20, 7.953217e-21, 1.749793e-20, -4.53474e-21, 
    3.054621e-20, -3.300315e-21, -3.514904e-21, 1.798053e-20, 2.31743e-20, 
    2.25263e-20, 1.026736e-20, 2.546579e-21, -1.431069e-20, -2.081719e-20, 
    -9.387512e-21, 1.733676e-20, -1.24201e-20, 3.152147e-21, -1.014919e-20, 
    -1.657284e-20, -6.798269e-21, -9.424555e-21, 1.138924e-20, 1.698675e-20, 
    -4.601729e-21, 5.406718e-20, -7.028128e-21, -4.97945e-21, -2.595185e-20, 
    -6.03743e-21, 3.007633e-20, -1.026369e-20, 1.869529e-20, 1.37625e-20, 
    5.721601e-21, 8.414129e-22, 2.691617e-21, -3.376399e-20, 4.693132e-20, 
    -3.383214e-20, 5.218647e-21, 5.563834e-21, -2.333857e-20, 4.870604e-21, 
    -1.171465e-20, -3.348092e-21, -1.952482e-20, 2.839097e-20, -1.580493e-20, 
    2.176859e-20, 5.754136e-21, 1.452499e-20, -4.382892e-21, -1.936649e-20, 
    2.307139e-20, 9.720291e-21, -3.863685e-20, -2.069504e-20, 2.101115e-20, 
    6.116876e-21, 1.266491e-20, 1.11108e-22, 3.812342e-20, -2.19611e-20, 
    -2.935961e-20, -2.860445e-20, -9.453383e-21, -3.659129e-20, 
    -2.680202e-20, 2.205186e-20, -7.625524e-21, 1.519988e-20, 1.842698e-20, 
    -3.221915e-20, -3.845138e-22, 1.930206e-21, 3.910732e-20, 1.676876e-20, 
    1.098323e-20, 3.685933e-20, 3.684577e-20, -2.656734e-20, -2.388e-20, 
    -1.993591e-20, -1.181419e-20, -6.689675e-21, -2.093509e-20, 
    -7.054415e-21, 5.388567e-20, 1.070702e-20, 1.690956e-20, 1.562483e-20, 
    -1.207034e-20, 2.298205e-20, 6.336268e-21, -4.857433e-22, 3.397659e-20, 
    -1.678406e-20, 4.000696e-20, -5.021016e-20, -8.47036e-21, 2.165521e-20, 
    1.707015e-20, -1.328494e-20, -1.916359e-21, 8.753644e-21, 1.268443e-20, 
    -1.266548e-20, 2.010769e-21, -3.949975e-20, -3.132401e-20, -6.281232e-20, 
    3.080906e-21, 1.63865e-20, -2.923728e-21, 1.6274e-20, 2.066111e-20, 
    -3.57287e-21, -1.545265e-20, 1.763335e-20, 1.849597e-20, -3.519093e-20, 
    3.657208e-20, 1.289734e-20, 1.036197e-21, -1.56961e-20, -3.0689e-20, 
    -9.52802e-21, 2.704855e-20, -2.619244e-20, 3.409593e-20, 2.196167e-20, 
    6.008602e-21, 3.07009e-20, -6.308012e-21, -2.785154e-20, -2.406265e-20, 
    4.037412e-21, -1.786406e-20, 1.465933e-20, 4.134673e-21, 1.830965e-20, 
    1.735628e-20, -7.319322e-21, -1.456104e-22, 6.048443e-21, -1.775522e-20, 
    -1.14226e-20, -1.471528e-20, 4.122778e-21, -8.642984e-22, -4.887275e-21, 
    4.686549e-21, 3.818138e-20, -1.489539e-20, 1.190664e-20, -3.661055e-21, 
    1.396423e-21, 1.424539e-20, -2.848741e-20, -2.045255e-21, 1.603566e-20, 
    -4.315689e-20, 1.952933e-20, 2.459729e-20, 1.803145e-20, -3.775277e-20, 
    -9.51842e-21, 3.373262e-21, 2.301316e-20, 8.162598e-22, 4.70693e-20, 
    2.553171e-20, -7.151899e-23, 9.50831e-22, 3.974091e-20, -7.350707e-21, 
    1.217383e-20, -2.092293e-20, 2.969918e-20, 9.214471e-21, 1.818948e-20, 
    -2.062831e-20, -1.793079e-20, 2.632875e-20, 9.434745e-21, 7.367127e-21, 
    -6.063867e-20, -3.945515e-21, -5.838678e-21, -9.122295e-21, 
    -2.184463e-20, 9.128231e-21, -2.720123e-20, 8.90008e-21, -8.958617e-21, 
    -1.634691e-20, -2.201284e-20, -2.171685e-20, 2.339117e-20, -1.177884e-20, 
    -4.017492e-20, 3.450702e-20, 9.081572e-21, -1.088258e-20, 1.790051e-20, 
    -1.196942e-20, 2.709974e-20, -7.672184e-21, 8.852302e-21, -1.007678e-20, 
    -6.100538e-20, 9.474178e-22, -1.409356e-20, 1.584736e-20, -4.150488e-21, 
    1.264287e-20, 7.517948e-22, -2.16914e-20, -1.357447e-20, 8.778837e-22, 
    -3.20845e-21, 6.272676e-21, -1.423805e-20, -3.143656e-20, 2.965959e-20, 
    2.305302e-20, -2.175586e-20, -2.87393e-20, 3.07582e-21, 2.941672e-20, 
    4.804995e-21 ;

 M_SOIL2C_TO_LEACHING =
  3.751187e-20, 1.027219e-20, 1.692002e-20, 1.451001e-20, 4.716233e-21, 
    3.176027e-20, 3.592574e-20, 1.883525e-20, 3.028061e-22, 2.655974e-20, 
    -1.280546e-20, -8.739487e-21, 2.851932e-20, -5.718499e-21, 1.099088e-20, 
    1.967843e-22, 3.599724e-21, -1.750498e-20, -3.350916e-21, -1.718071e-20, 
    1.010989e-20, 1.684822e-20, -5.419367e-21, 1.658102e-20, -1.514051e-20, 
    -7.773414e-21, -1.698393e-20, 1.347298e-20, 1.198609e-20, -2.366511e-22, 
    -2.521278e-20, -3.970685e-21, -1.046556e-20, 2.821364e-21, -2.903729e-20, 
    4.399842e-21, -2.171626e-20, 1.182379e-21, -2.922021e-21, 3.05024e-20, 
    2.291872e-20, -2.295717e-20, 4.897742e-21, -3.719606e-20, -7.345346e-22, 
    -4.75881e-20, 3.212104e-20, 4.666177e-21, -1.930316e-20, -4.329457e-21, 
    1.766586e-20, 2.191898e-20, -1.143701e-20, 2.716759e-20, 4.911769e-20, 
    -3.44123e-20, -6.790905e-21, 5.44342e-21, 2.155058e-20, -2.911026e-20, 
    2.212566e-20, 1.922088e-20, 1.35759e-20, 1.714903e-20, 4.569505e-21, 
    2.310928e-20, 4.527509e-20, -1.724121e-20, -2.331596e-20, 2.274852e-21, 
    7.065312e-22, -2.1608e-20, 7.149677e-21, 2.47169e-20, -2.793721e-20, 
    1.112151e-20, 2.91761e-20, 6.648128e-21, 3.078286e-20, 8.188761e-24, 
    -6.126577e-20, 3.396474e-20, -1.914484e-20, -3.599332e-20, -2.790808e-20, 
    1.021252e-20, -2.982327e-20, -1.169601e-20, 5.68894e-20, -8.615651e-21, 
    -1.378455e-20, 2.126418e-20, -1.395134e-20, -1.0601e-20, 1.057526e-20, 
    -1.106976e-20, -2.519303e-20, -1.666499e-20, -1.166548e-20, 
    -1.991753e-20, -1.902127e-20, 2.757246e-20, 2.869407e-20, 1.534777e-20, 
    2.368664e-20, -3.484459e-20, -5.657447e-22, 1.094752e-21, 1.474752e-20, 
    -1.394115e-20, -3.107155e-20, 1.80713e-20, 2.155262e-21, -2.109001e-20, 
    2.086017e-20, -2.405529e-20, 3.893372e-20, 3.615985e-20, -9.073972e-21, 
    1.764581e-20, -1.516791e-20, -2.227918e-20, 3.531307e-20, -1.052382e-20, 
    -1.434209e-20, -2.318923e-21, -2.805341e-20, 4.033748e-20, -5.614157e-20, 
    1.13234e-21, -1.774816e-20, -3.203273e-22, 1.106976e-20, -4.141836e-20, 
    2.223959e-20, 3.352848e-20, -1.791241e-20, 2.2541e-20, 1.426405e-20, 
    -5.661977e-21, 2.347882e-20, 1.231319e-20, -1.953048e-20, -3.945851e-20, 
    4.804077e-20, -4.297141e-20, 3.530457e-21, 8.874631e-21, -6.79237e-24, 
    2.868388e-20, 4.609639e-21, -3.846581e-20, 3.430174e-20, -3.362206e-20, 
    1.252209e-21, -1.14325e-20, 2.234676e-20, 1.514307e-20, -2.668699e-21, 
    -4.302795e-20, 2.538838e-20, 2.468154e-20, -5.44342e-21, 3.543634e-20, 
    -1.33221e-21, 2.769774e-20, 4.01789e-21, -1.629106e-21, -3.713554e-20, 
    -8.734974e-21, 1.681426e-20, -2.963357e-20, -5.550034e-20, -2.253081e-20, 
    3.59232e-20, -2.660072e-20, -1.783692e-20, 3.122309e-20, -4.31583e-20, 
    -3.04811e-21, -3.727241e-21, -3.31584e-20, 1.346448e-20, -2.046321e-20, 
    2.364477e-20, -6.594693e-21, -1.07859e-20, -1.332906e-20, 2.257521e-20, 
    -3.864165e-20, 1.043929e-20, 2.769264e-20, 3.512705e-20, -1.784595e-21, 
    -2.178163e-21, -3.145943e-21, 5.851962e-20, 1.862462e-20, 3.868321e-21, 
    -1.844026e-20, -1.95839e-20, -1.490982e-20, 2.068289e-20, -2.525944e-20, 
    4.986243e-21, -1.699891e-20, 6.755857e-21, -9.735288e-21, -1.721264e-21, 
    1.826948e-20, -8.032101e-21, -4.528209e-21, 2.356053e-20, -4.250859e-20, 
    -4.118809e-21, -2.623967e-20, 2.652176e-22, 2.472227e-20, -1.541249e-20, 
    -2.660412e-20, 3.763713e-21, -1.758926e-20, -2.895446e-20, -2.597446e-20, 
    1.246901e-20, 2.59264e-21, 3.290158e-21, 1.183877e-20, 1.19813e-20, 
    1.806536e-20, 4.782701e-20, 1.671731e-20, -1.718662e-20, 3.818195e-20, 
    2.071739e-20, 4.058883e-20, -4.395612e-21, 4.093378e-21, 1.866757e-20, 
    -7.919832e-21, -4.122215e-20, -1.357702e-20, 2.521278e-20, 1.164878e-20, 
    -4.112327e-21, 8.596139e-21, 2.365893e-21, -7.498983e-20, 1.213849e-20, 
    1.477098e-20, -3.544625e-20, -1.373367e-20, 7.123111e-21, -2.627757e-20, 
    1.790844e-20, -2.51178e-20, 8.742312e-21, 4.013066e-21, 1.06663e-20, 
    -3.552175e-20, 1.085123e-20, 1.016531e-20, 1.516143e-20, 1.750189e-20, 
    -3.00803e-20, -3.020836e-20, -1.812757e-20, -3.467127e-21, -2.103489e-20, 
    -6.705228e-21, -1.768849e-20, 8.43896e-21, -1.689768e-20, -3.782662e-21, 
    -8.234533e-21, -1.902977e-20, -3.689721e-20, 9.055938e-22, 5.904832e-21, 
    1.475542e-21, 3.534687e-21, 8.960848e-21, -1.261063e-20, 9.946465e-21, 
    3.476203e-20, 1.472829e-20, -9.579782e-21, -1.127809e-21, 4.267848e-20, 
    2.260404e-20, -2.203573e-20, -7.41376e-21, -1.227617e-20, -9.443685e-23, 
    -2.802709e-20, -1.613943e-20, 1.144381e-20, 3.428167e-20, 7.936546e-21, 
    2.707261e-20, 1.566921e-20, 2.355601e-20, 2.526906e-20, -7.315119e-21, 
    3.022026e-20, -1.142374e-20, -4.834647e-22, -1.799581e-20, 1.402911e-20, 
    2.657359e-20, -1.767073e-21, 1.968824e-20, 2.361649e-20, 8.009494e-21, 
    2.758153e-20, -6.715989e-21, -1.029422e-20, 2.894539e-20, -1.638412e-21, 
    2.89785e-20, -8.040856e-22, -1.0558e-20, 2.024268e-20, 9.043983e-21, 
    2.554302e-20, -4.35292e-21, -3.140149e-20, 3.80451e-20, -2.345254e-21, 
    -1.456968e-20, -9.132421e-22, -5.45756e-21, 4.911259e-20, -3.114081e-20, 
    3.357709e-21, 3.771799e-20, 7.591497e-22, -1.954149e-20 ;

 M_SOIL3C_TO_LEACHING =
  -2.598407e-20, -2.739605e-20, -3.173766e-20, -6.308868e-21, -1.320126e-20, 
    7.097107e-21, -3.44123e-20, 2.649753e-20, -3.209584e-21, 4.697572e-20, 
    3.21493e-20, -4.84425e-20, 9.322182e-21, 1.469039e-20, -1.21351e-20, 
    -2.851326e-21, -1.193831e-20, -3.204244e-20, 3.312162e-20, -2.691626e-20, 
    7.158185e-21, 2.376973e-20, 1.827318e-20, 2.261006e-21, 7.982355e-21, 
    -2.918064e-20, -8.895859e-21, -9.997633e-21, -4.800791e-21, 1.40667e-20, 
    1.047094e-20, 8.533943e-21, -1.714677e-20, -1.821975e-20, 6.411494e-21, 
    3.963321e-21, -1.895597e-20, -4.255182e-20, -2.695981e-20, -1.731359e-20, 
    -7.94106e-21, 8.252875e-22, -1.521546e-20, 1.327535e-20, 7.634286e-21, 
    -1.12821e-20, 4.936759e-21, 3.940975e-21, 2.441663e-20, 2.989653e-20, 
    -2.91467e-20, 7.263367e-22, -2.125117e-20, -2.014457e-20, 1.091368e-20, 
    9.769203e-21, -2.304792e-20, -2.588118e-20, 1.059024e-20, -5.505354e-21, 
    -3.710729e-20, 1.928252e-20, -3.050127e-20, 3.113005e-20, 1.369406e-20, 
    1.765287e-20, 4.096826e-20, 1.505769e-20, -3.518872e-21, 9.575252e-21, 
    2.7156e-20, 2.111436e-21, -2.566687e-20, 1.046812e-20, -1.435792e-20, 
    -3.217278e-20, 1.494458e-20, 7.730412e-21, -6.353249e-21, 3.842791e-20, 
    -1.585412e-20, -2.084574e-20, 2.154379e-20, 7.876612e-21, -1.866041e-21, 
    5.881941e-21, 2.318688e-21, -2.993214e-20, -2.413052e-20, 5.811447e-20, 
    3.712453e-20, 1.328297e-20, -2.713593e-20, -3.945254e-20, -1.223674e-21, 
    1.540684e-20, -7.40183e-22, 1.78601e-20, 5.280288e-21, -2.65289e-20, 
    -9.70193e-21, -2.949138e-20, 4.142862e-21, 1.045311e-20, 1.429231e-20, 
    -2.890914e-21, 2.288716e-21, 2.526227e-20, -3.996767e-20, 7.874333e-21, 
    -2.277677e-20, -1.558353e-20, -2.954821e-20, 3.807733e-20, -8.544965e-21, 
    -1.693615e-20, -1.47625e-20, 9.95637e-21, 8.168319e-22, -3.143907e-22, 
    -4.162842e-20, 1.368812e-20, 1.585612e-20, 3.398481e-20, 1.308279e-20, 
    -7.352707e-21, -3.771649e-21, 5.244092e-20, 2.263401e-20, 2.141801e-20, 
    6.124241e-21, -2.37949e-20, -2.294729e-20, 1.526212e-20, -5.631705e-21, 
    -7.736366e-21, 2.001819e-20, 3.999198e-20, -2.48735e-20, -2.229416e-20, 
    -2.258538e-20, 1.058884e-20, 3.226255e-21, 1.183965e-20, -1.473028e-21, 
    5.540818e-20, 1.01701e-20, 2.519697e-20, -2.421731e-20, 3.728343e-20, 
    -1.508822e-20, -3.935872e-21, -4.297805e-21, 2.269028e-20, 3.052136e-20, 
    -3.046992e-21, 2.877295e-20, -1.422589e-20, -2.544067e-20, 4.13406e-20, 
    -1.162596e-21, -1.582926e-20, -2.809325e-20, 1.491402e-20, 2.635531e-20, 
    -1.371075e-20, -2.173077e-21, 5.802485e-21, -1.667687e-20, 1.565423e-20, 
    2.524929e-20, 6.406391e-21, -3.715084e-21, 3.656868e-20, -2.234958e-20, 
    -1.965657e-20, -7.293035e-21, -8.500584e-21, 3.058299e-20, -1.165136e-21, 
    -4.41003e-21, -1.479812e-20, 2.518558e-21, 8.688297e-21, 1.159003e-22, 
    2.65428e-21, -6.002666e-21, -1.989125e-20, 1.368671e-20, -5.422764e-21, 
    3.297202e-21, -3.701003e-20, 2.018897e-20, -2.397244e-20, -8.882273e-21, 
    1.07927e-20, 2.849956e-20, 9.623308e-21, 2.134221e-20, 3.172248e-22, 
    -4.799554e-20, -2.242507e-20, 1.337401e-20, -2.970595e-20, 2.302897e-20, 
    -2.858068e-20, 4.498302e-20, 2.731208e-20, -1.381987e-21, -2.534967e-21, 
    1.496351e-20, -5.646686e-21, -3.633376e-21, 2.684586e-20, 2.484665e-20, 
    1.702125e-20, 1.157275e-20, 4.222555e-20, 2.341774e-20, -3.704284e-20, 
    -2.48236e-22, 1.950644e-20, 2.322858e-20, 1.645602e-22, -1.454734e-20, 
    6.390276e-23, 3.973509e-21, -4.742439e-20, 9.285165e-21, 2.240925e-20, 
    -1.354216e-22, 2.715968e-20, -1.744875e-20, 1.481507e-20, -4.840576e-20, 
    -1.098409e-21, -9.322492e-21, 3.223683e-21, -1.25917e-20, 2.334503e-21, 
    1.72446e-20, 6.464635e-21, 4.076783e-20, -8.969346e-21, -1.565763e-20, 
    -1.281337e-20, -4.908264e-20, 1.148454e-20, 2.125854e-20, 2.793097e-20, 
    -5.559613e-21, 2.65326e-20, -2.172872e-20, -3.771687e-20, 6.789215e-21, 
    4.366767e-21, 2.101532e-21, -1.832632e-20, 1.506163e-20, 2.332812e-20, 
    -5.068658e-20, 4.65587e-20, -2.811675e-20, -1.225326e-20, 1.039657e-20, 
    4.650875e-22, 1.100688e-21, 8.047654e-21, -2.052317e-20, -3.345552e-21, 
    2.768245e-20, 7.278338e-21, -1.242461e-20, 1.117608e-20, -1.604214e-20, 
    -4.877968e-21, -1.205196e-20, -1.727061e-20, 4.657086e-20, -3.512137e-20, 
    1.578317e-20, -4.95174e-21, -6.317629e-21, -6.045929e-21, -2.702822e-20, 
    1.923983e-20, -1.840324e-20, 2.805238e-21, -3.395343e-20, -1.487726e-20, 
    -8.481635e-21, 3.399004e-21, -4.245625e-20, 3.100057e-20, 1.560731e-20, 
    -1.786518e-20, -8.880012e-21, -1.331068e-20, 3.215694e-20, -7.135578e-21, 
    -3.684828e-21, 6.498566e-21, -1.389538e-20, -2.509009e-20, 2.07383e-20, 
    -1.646002e-20, 8.27863e-21, -5.597513e-21, -1.500143e-20, -1.023317e-20, 
    -1.913508e-21, -4.213535e-20, 7.288544e-21, 3.198759e-20, 3.232207e-20, 
    8.844113e-21, 3.937592e-20, -2.396679e-20, 2.858183e-20, 2.790862e-20, 
    -3.823368e-21, -8.32897e-21, 3.233899e-21, 2.590578e-20, -8.385508e-21, 
    -4.490032e-21, -2.586845e-20, -3.708292e-21, 5.490625e-21, 9.305805e-21, 
    -1.521318e-20, -4.629749e-21, -1.474158e-20, -6.217109e-20, 
    -2.092999e-20, -3.862663e-21, -5.991887e-20, 1.653126e-20 ;

 NBP =
  -6.194416e-08, -6.221921e-08, -6.216575e-08, -6.238761e-08, -6.226454e-08, 
    -6.240981e-08, -6.199993e-08, -6.223013e-08, -6.208317e-08, 
    -6.196893e-08, -6.281821e-08, -6.239751e-08, -6.325536e-08, 
    -6.298698e-08, -6.366125e-08, -6.321359e-08, -6.375153e-08, 
    -6.364835e-08, -6.395895e-08, -6.386996e-08, -6.426725e-08, 
    -6.400002e-08, -6.447324e-08, -6.420344e-08, -6.424563e-08, -6.39912e-08, 
    -6.248218e-08, -6.276583e-08, -6.246538e-08, -6.250582e-08, 
    -6.248767e-08, -6.226708e-08, -6.215591e-08, -6.192315e-08, -6.19654e-08, 
    -6.213637e-08, -6.2524e-08, -6.239242e-08, -6.272409e-08, -6.27166e-08, 
    -6.308589e-08, -6.291938e-08, -6.354018e-08, -6.336372e-08, 
    -6.387368e-08, -6.374542e-08, -6.386765e-08, -6.383059e-08, 
    -6.386814e-08, -6.368003e-08, -6.376062e-08, -6.359511e-08, 
    -6.295056e-08, -6.313996e-08, -6.25751e-08, -6.223551e-08, -6.201002e-08, 
    -6.185e-08, -6.187263e-08, -6.191575e-08, -6.213737e-08, -6.234576e-08, 
    -6.250459e-08, -6.261083e-08, -6.271553e-08, -6.303241e-08, 
    -6.320018e-08, -6.357585e-08, -6.350807e-08, -6.362291e-08, 
    -6.373266e-08, -6.39169e-08, -6.388658e-08, -6.396775e-08, -6.361989e-08, 
    -6.385107e-08, -6.346945e-08, -6.357381e-08, -6.274394e-08, 
    -6.242792e-08, -6.229357e-08, -6.217602e-08, -6.189002e-08, 
    -6.208752e-08, -6.200966e-08, -6.219491e-08, -6.231262e-08, -6.22544e-08, 
    -6.261374e-08, -6.247403e-08, -6.321012e-08, -6.289304e-08, 
    -6.371985e-08, -6.352198e-08, -6.376729e-08, -6.364211e-08, -6.38566e-08, 
    -6.366356e-08, -6.399797e-08, -6.407078e-08, -6.402102e-08, 
    -6.421219e-08, -6.365286e-08, -6.386765e-08, -6.225277e-08, 
    -6.226226e-08, -6.23065e-08, -6.211204e-08, -6.210015e-08, -6.192198e-08, 
    -6.208052e-08, -6.214803e-08, -6.231944e-08, -6.242083e-08, 
    -6.251722e-08, -6.272915e-08, -6.296587e-08, -6.329692e-08, 
    -6.353481e-08, -6.369427e-08, -6.359649e-08, -6.368282e-08, 
    -6.358631e-08, -6.354109e-08, -6.40435e-08, -6.376137e-08, -6.41847e-08, 
    -6.416128e-08, -6.396969e-08, -6.416391e-08, -6.226892e-08, 
    -6.221429e-08, -6.202459e-08, -6.217304e-08, -6.190258e-08, 
    -6.205396e-08, -6.214101e-08, -6.247694e-08, -6.255076e-08, -6.26192e-08, 
    -6.27544e-08, -6.29279e-08, -6.32323e-08, -6.349719e-08, -6.373904e-08, 
    -6.372132e-08, -6.372756e-08, -6.378159e-08, -6.364776e-08, 
    -6.380356e-08, -6.38297e-08, -6.376134e-08, -6.415814e-08, -6.404477e-08, 
    -6.416078e-08, -6.408697e-08, -6.223205e-08, -6.232399e-08, 
    -6.227431e-08, -6.236773e-08, -6.230191e-08, -6.259458e-08, 
    -6.268234e-08, -6.309303e-08, -6.292449e-08, -6.319274e-08, 
    -6.295173e-08, -6.299444e-08, -6.320148e-08, -6.296477e-08, 
    -6.348257e-08, -6.313149e-08, -6.378369e-08, -6.343302e-08, 
    -6.380566e-08, -6.3738e-08, -6.385004e-08, -6.395038e-08, -6.407663e-08, 
    -6.430958e-08, -6.425564e-08, -6.445048e-08, -6.246106e-08, 
    -6.258032e-08, -6.256982e-08, -6.269464e-08, -6.278695e-08, 
    -6.298706e-08, -6.330801e-08, -6.318732e-08, -6.340892e-08, 
    -6.345341e-08, -6.311675e-08, -6.332343e-08, -6.266014e-08, 
    -6.276728e-08, -6.27035e-08, -6.247047e-08, -6.321512e-08, -6.283292e-08, 
    -6.353874e-08, -6.333165e-08, -6.393607e-08, -6.363545e-08, 
    -6.422594e-08, -6.447839e-08, -6.471606e-08, -6.499378e-08, 
    -6.264541e-08, -6.256438e-08, -6.270949e-08, -6.291025e-08, 
    -6.309657e-08, -6.334428e-08, -6.336963e-08, -6.341604e-08, 
    -6.353626e-08, -6.363734e-08, -6.34307e-08, -6.366268e-08, -6.279212e-08, 
    -6.32483e-08, -6.253374e-08, -6.274887e-08, -6.289842e-08, -6.283283e-08, 
    -6.317353e-08, -6.325383e-08, -6.358018e-08, -6.341148e-08, 
    -6.441608e-08, -6.397156e-08, -6.52053e-08, -6.486045e-08, -6.253607e-08, 
    -6.264514e-08, -6.302479e-08, -6.284415e-08, -6.336082e-08, 
    -6.348802e-08, -6.359143e-08, -6.372361e-08, -6.373789e-08, 
    -6.381621e-08, -6.368786e-08, -6.381114e-08, -6.334481e-08, 
    -6.355319e-08, -6.298141e-08, -6.312055e-08, -6.305654e-08, 
    -6.298632e-08, -6.320305e-08, -6.343395e-08, -6.34389e-08, -6.351294e-08, 
    -6.372157e-08, -6.336292e-08, -6.447343e-08, -6.378752e-08, 
    -6.276409e-08, -6.297419e-08, -6.300422e-08, -6.292283e-08, 
    -6.347526e-08, -6.327508e-08, -6.38143e-08, -6.366856e-08, -6.390736e-08, 
    -6.37887e-08, -6.377123e-08, -6.361883e-08, -6.352395e-08, -6.328425e-08, 
    -6.308925e-08, -6.293464e-08, -6.297059e-08, -6.314043e-08, 
    -6.344808e-08, -6.373917e-08, -6.367541e-08, -6.388921e-08, 
    -6.332336e-08, -6.356061e-08, -6.34689e-08, -6.370803e-08, -6.318411e-08, 
    -6.36302e-08, -6.307009e-08, -6.31192e-08, -6.327111e-08, -6.357669e-08, 
    -6.364433e-08, -6.371651e-08, -6.367197e-08, -6.34559e-08, -6.34205e-08, 
    -6.326741e-08, -6.322514e-08, -6.310851e-08, -6.301195e-08, 
    -6.310017e-08, -6.319282e-08, -6.345599e-08, -6.369318e-08, -6.39518e-08, 
    -6.401511e-08, -6.431729e-08, -6.407128e-08, -6.447725e-08, 
    -6.413207e-08, -6.472964e-08, -6.365608e-08, -6.412193e-08, 
    -6.327802e-08, -6.336893e-08, -6.353335e-08, -6.391052e-08, 
    -6.370691e-08, -6.394504e-08, -6.341912e-08, -6.314629e-08, 
    -6.307572e-08, -6.294403e-08, -6.307872e-08, -6.306777e-08, 
    -6.319667e-08, -6.315525e-08, -6.346473e-08, -6.329849e-08, 
    -6.377079e-08, -6.394317e-08, -6.443005e-08, -6.472857e-08, 
    -6.503251e-08, -6.51667e-08, -6.520754e-08, -6.522462e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.194416e-08, 6.221921e-08, 6.216575e-08, 6.238761e-08, 6.226454e-08, 
    6.240981e-08, 6.199993e-08, 6.223013e-08, 6.208317e-08, 6.196893e-08, 
    6.281821e-08, 6.239751e-08, 6.325536e-08, 6.298698e-08, 6.366125e-08, 
    6.321359e-08, 6.375153e-08, 6.364835e-08, 6.395895e-08, 6.386996e-08, 
    6.426725e-08, 6.400002e-08, 6.447324e-08, 6.420344e-08, 6.424563e-08, 
    6.39912e-08, 6.248218e-08, 6.276583e-08, 6.246538e-08, 6.250582e-08, 
    6.248767e-08, 6.226708e-08, 6.215591e-08, 6.192315e-08, 6.19654e-08, 
    6.213637e-08, 6.2524e-08, 6.239242e-08, 6.272409e-08, 6.27166e-08, 
    6.308589e-08, 6.291938e-08, 6.354018e-08, 6.336372e-08, 6.387368e-08, 
    6.374542e-08, 6.386765e-08, 6.383059e-08, 6.386814e-08, 6.368003e-08, 
    6.376062e-08, 6.359511e-08, 6.295056e-08, 6.313996e-08, 6.25751e-08, 
    6.223551e-08, 6.201002e-08, 6.185e-08, 6.187263e-08, 6.191575e-08, 
    6.213737e-08, 6.234576e-08, 6.250459e-08, 6.261083e-08, 6.271553e-08, 
    6.303241e-08, 6.320018e-08, 6.357585e-08, 6.350807e-08, 6.362291e-08, 
    6.373266e-08, 6.39169e-08, 6.388658e-08, 6.396775e-08, 6.361989e-08, 
    6.385107e-08, 6.346945e-08, 6.357381e-08, 6.274394e-08, 6.242792e-08, 
    6.229357e-08, 6.217602e-08, 6.189002e-08, 6.208752e-08, 6.200966e-08, 
    6.219491e-08, 6.231262e-08, 6.22544e-08, 6.261374e-08, 6.247403e-08, 
    6.321012e-08, 6.289304e-08, 6.371985e-08, 6.352198e-08, 6.376729e-08, 
    6.364211e-08, 6.38566e-08, 6.366356e-08, 6.399797e-08, 6.407078e-08, 
    6.402102e-08, 6.421219e-08, 6.365286e-08, 6.386765e-08, 6.225277e-08, 
    6.226226e-08, 6.23065e-08, 6.211204e-08, 6.210015e-08, 6.192198e-08, 
    6.208052e-08, 6.214803e-08, 6.231944e-08, 6.242083e-08, 6.251722e-08, 
    6.272915e-08, 6.296587e-08, 6.329692e-08, 6.353481e-08, 6.369427e-08, 
    6.359649e-08, 6.368282e-08, 6.358631e-08, 6.354109e-08, 6.40435e-08, 
    6.376137e-08, 6.41847e-08, 6.416128e-08, 6.396969e-08, 6.416391e-08, 
    6.226892e-08, 6.221429e-08, 6.202459e-08, 6.217304e-08, 6.190258e-08, 
    6.205396e-08, 6.214101e-08, 6.247694e-08, 6.255076e-08, 6.26192e-08, 
    6.27544e-08, 6.29279e-08, 6.32323e-08, 6.349719e-08, 6.373904e-08, 
    6.372132e-08, 6.372756e-08, 6.378159e-08, 6.364776e-08, 6.380356e-08, 
    6.38297e-08, 6.376134e-08, 6.415814e-08, 6.404477e-08, 6.416078e-08, 
    6.408697e-08, 6.223205e-08, 6.232399e-08, 6.227431e-08, 6.236773e-08, 
    6.230191e-08, 6.259458e-08, 6.268234e-08, 6.309303e-08, 6.292449e-08, 
    6.319274e-08, 6.295173e-08, 6.299444e-08, 6.320148e-08, 6.296477e-08, 
    6.348257e-08, 6.313149e-08, 6.378369e-08, 6.343302e-08, 6.380566e-08, 
    6.3738e-08, 6.385004e-08, 6.395038e-08, 6.407663e-08, 6.430958e-08, 
    6.425564e-08, 6.445048e-08, 6.246106e-08, 6.258032e-08, 6.256982e-08, 
    6.269464e-08, 6.278695e-08, 6.298706e-08, 6.330801e-08, 6.318732e-08, 
    6.340892e-08, 6.345341e-08, 6.311675e-08, 6.332343e-08, 6.266014e-08, 
    6.276728e-08, 6.27035e-08, 6.247047e-08, 6.321512e-08, 6.283292e-08, 
    6.353874e-08, 6.333165e-08, 6.393607e-08, 6.363545e-08, 6.422594e-08, 
    6.447839e-08, 6.471606e-08, 6.499378e-08, 6.264541e-08, 6.256438e-08, 
    6.270949e-08, 6.291025e-08, 6.309657e-08, 6.334428e-08, 6.336963e-08, 
    6.341604e-08, 6.353626e-08, 6.363734e-08, 6.34307e-08, 6.366268e-08, 
    6.279212e-08, 6.32483e-08, 6.253374e-08, 6.274887e-08, 6.289842e-08, 
    6.283283e-08, 6.317353e-08, 6.325383e-08, 6.358018e-08, 6.341148e-08, 
    6.441608e-08, 6.397156e-08, 6.52053e-08, 6.486045e-08, 6.253607e-08, 
    6.264514e-08, 6.302479e-08, 6.284415e-08, 6.336082e-08, 6.348802e-08, 
    6.359143e-08, 6.372361e-08, 6.373789e-08, 6.381621e-08, 6.368786e-08, 
    6.381114e-08, 6.334481e-08, 6.355319e-08, 6.298141e-08, 6.312055e-08, 
    6.305654e-08, 6.298632e-08, 6.320305e-08, 6.343395e-08, 6.34389e-08, 
    6.351294e-08, 6.372157e-08, 6.336292e-08, 6.447343e-08, 6.378752e-08, 
    6.276409e-08, 6.297419e-08, 6.300422e-08, 6.292283e-08, 6.347526e-08, 
    6.327508e-08, 6.38143e-08, 6.366856e-08, 6.390736e-08, 6.37887e-08, 
    6.377123e-08, 6.361883e-08, 6.352395e-08, 6.328425e-08, 6.308925e-08, 
    6.293464e-08, 6.297059e-08, 6.314043e-08, 6.344808e-08, 6.373917e-08, 
    6.367541e-08, 6.388921e-08, 6.332336e-08, 6.356061e-08, 6.34689e-08, 
    6.370803e-08, 6.318411e-08, 6.36302e-08, 6.307009e-08, 6.31192e-08, 
    6.327111e-08, 6.357669e-08, 6.364433e-08, 6.371651e-08, 6.367197e-08, 
    6.34559e-08, 6.34205e-08, 6.326741e-08, 6.322514e-08, 6.310851e-08, 
    6.301195e-08, 6.310017e-08, 6.319282e-08, 6.345599e-08, 6.369318e-08, 
    6.39518e-08, 6.401511e-08, 6.431729e-08, 6.407128e-08, 6.447725e-08, 
    6.413207e-08, 6.472964e-08, 6.365608e-08, 6.412193e-08, 6.327802e-08, 
    6.336893e-08, 6.353335e-08, 6.391052e-08, 6.370691e-08, 6.394504e-08, 
    6.341912e-08, 6.314629e-08, 6.307572e-08, 6.294403e-08, 6.307872e-08, 
    6.306777e-08, 6.319667e-08, 6.315525e-08, 6.346473e-08, 6.329849e-08, 
    6.377079e-08, 6.394317e-08, 6.443005e-08, 6.472857e-08, 6.503251e-08, 
    6.51667e-08, 6.520754e-08, 6.522462e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.194416e-08, -6.221921e-08, -6.216575e-08, -6.238761e-08, -6.226454e-08, 
    -6.240981e-08, -6.199993e-08, -6.223013e-08, -6.208317e-08, 
    -6.196893e-08, -6.281821e-08, -6.239751e-08, -6.325536e-08, 
    -6.298698e-08, -6.366125e-08, -6.321359e-08, -6.375153e-08, 
    -6.364835e-08, -6.395895e-08, -6.386996e-08, -6.426725e-08, 
    -6.400002e-08, -6.447324e-08, -6.420344e-08, -6.424563e-08, -6.39912e-08, 
    -6.248218e-08, -6.276583e-08, -6.246538e-08, -6.250582e-08, 
    -6.248767e-08, -6.226708e-08, -6.215591e-08, -6.192315e-08, -6.19654e-08, 
    -6.213637e-08, -6.2524e-08, -6.239242e-08, -6.272409e-08, -6.27166e-08, 
    -6.308589e-08, -6.291938e-08, -6.354018e-08, -6.336372e-08, 
    -6.387368e-08, -6.374542e-08, -6.386765e-08, -6.383059e-08, 
    -6.386814e-08, -6.368003e-08, -6.376062e-08, -6.359511e-08, 
    -6.295056e-08, -6.313996e-08, -6.25751e-08, -6.223551e-08, -6.201002e-08, 
    -6.185e-08, -6.187263e-08, -6.191575e-08, -6.213737e-08, -6.234576e-08, 
    -6.250459e-08, -6.261083e-08, -6.271553e-08, -6.303241e-08, 
    -6.320018e-08, -6.357585e-08, -6.350807e-08, -6.362291e-08, 
    -6.373266e-08, -6.39169e-08, -6.388658e-08, -6.396775e-08, -6.361989e-08, 
    -6.385107e-08, -6.346945e-08, -6.357381e-08, -6.274394e-08, 
    -6.242792e-08, -6.229357e-08, -6.217602e-08, -6.189002e-08, 
    -6.208752e-08, -6.200966e-08, -6.219491e-08, -6.231262e-08, -6.22544e-08, 
    -6.261374e-08, -6.247403e-08, -6.321012e-08, -6.289304e-08, 
    -6.371985e-08, -6.352198e-08, -6.376729e-08, -6.364211e-08, -6.38566e-08, 
    -6.366356e-08, -6.399797e-08, -6.407078e-08, -6.402102e-08, 
    -6.421219e-08, -6.365286e-08, -6.386765e-08, -6.225277e-08, 
    -6.226226e-08, -6.23065e-08, -6.211204e-08, -6.210015e-08, -6.192198e-08, 
    -6.208052e-08, -6.214803e-08, -6.231944e-08, -6.242083e-08, 
    -6.251722e-08, -6.272915e-08, -6.296587e-08, -6.329692e-08, 
    -6.353481e-08, -6.369427e-08, -6.359649e-08, -6.368282e-08, 
    -6.358631e-08, -6.354109e-08, -6.40435e-08, -6.376137e-08, -6.41847e-08, 
    -6.416128e-08, -6.396969e-08, -6.416391e-08, -6.226892e-08, 
    -6.221429e-08, -6.202459e-08, -6.217304e-08, -6.190258e-08, 
    -6.205396e-08, -6.214101e-08, -6.247694e-08, -6.255076e-08, -6.26192e-08, 
    -6.27544e-08, -6.29279e-08, -6.32323e-08, -6.349719e-08, -6.373904e-08, 
    -6.372132e-08, -6.372756e-08, -6.378159e-08, -6.364776e-08, 
    -6.380356e-08, -6.38297e-08, -6.376134e-08, -6.415814e-08, -6.404477e-08, 
    -6.416078e-08, -6.408697e-08, -6.223205e-08, -6.232399e-08, 
    -6.227431e-08, -6.236773e-08, -6.230191e-08, -6.259458e-08, 
    -6.268234e-08, -6.309303e-08, -6.292449e-08, -6.319274e-08, 
    -6.295173e-08, -6.299444e-08, -6.320148e-08, -6.296477e-08, 
    -6.348257e-08, -6.313149e-08, -6.378369e-08, -6.343302e-08, 
    -6.380566e-08, -6.3738e-08, -6.385004e-08, -6.395038e-08, -6.407663e-08, 
    -6.430958e-08, -6.425564e-08, -6.445048e-08, -6.246106e-08, 
    -6.258032e-08, -6.256982e-08, -6.269464e-08, -6.278695e-08, 
    -6.298706e-08, -6.330801e-08, -6.318732e-08, -6.340892e-08, 
    -6.345341e-08, -6.311675e-08, -6.332343e-08, -6.266014e-08, 
    -6.276728e-08, -6.27035e-08, -6.247047e-08, -6.321512e-08, -6.283292e-08, 
    -6.353874e-08, -6.333165e-08, -6.393607e-08, -6.363545e-08, 
    -6.422594e-08, -6.447839e-08, -6.471606e-08, -6.499378e-08, 
    -6.264541e-08, -6.256438e-08, -6.270949e-08, -6.291025e-08, 
    -6.309657e-08, -6.334428e-08, -6.336963e-08, -6.341604e-08, 
    -6.353626e-08, -6.363734e-08, -6.34307e-08, -6.366268e-08, -6.279212e-08, 
    -6.32483e-08, -6.253374e-08, -6.274887e-08, -6.289842e-08, -6.283283e-08, 
    -6.317353e-08, -6.325383e-08, -6.358018e-08, -6.341148e-08, 
    -6.441608e-08, -6.397156e-08, -6.52053e-08, -6.486045e-08, -6.253607e-08, 
    -6.264514e-08, -6.302479e-08, -6.284415e-08, -6.336082e-08, 
    -6.348802e-08, -6.359143e-08, -6.372361e-08, -6.373789e-08, 
    -6.381621e-08, -6.368786e-08, -6.381114e-08, -6.334481e-08, 
    -6.355319e-08, -6.298141e-08, -6.312055e-08, -6.305654e-08, 
    -6.298632e-08, -6.320305e-08, -6.343395e-08, -6.34389e-08, -6.351294e-08, 
    -6.372157e-08, -6.336292e-08, -6.447343e-08, -6.378752e-08, 
    -6.276409e-08, -6.297419e-08, -6.300422e-08, -6.292283e-08, 
    -6.347526e-08, -6.327508e-08, -6.38143e-08, -6.366856e-08, -6.390736e-08, 
    -6.37887e-08, -6.377123e-08, -6.361883e-08, -6.352395e-08, -6.328425e-08, 
    -6.308925e-08, -6.293464e-08, -6.297059e-08, -6.314043e-08, 
    -6.344808e-08, -6.373917e-08, -6.367541e-08, -6.388921e-08, 
    -6.332336e-08, -6.356061e-08, -6.34689e-08, -6.370803e-08, -6.318411e-08, 
    -6.36302e-08, -6.307009e-08, -6.31192e-08, -6.327111e-08, -6.357669e-08, 
    -6.364433e-08, -6.371651e-08, -6.367197e-08, -6.34559e-08, -6.34205e-08, 
    -6.326741e-08, -6.322514e-08, -6.310851e-08, -6.301195e-08, 
    -6.310017e-08, -6.319282e-08, -6.345599e-08, -6.369318e-08, -6.39518e-08, 
    -6.401511e-08, -6.431729e-08, -6.407128e-08, -6.447725e-08, 
    -6.413207e-08, -6.472964e-08, -6.365608e-08, -6.412193e-08, 
    -6.327802e-08, -6.336893e-08, -6.353335e-08, -6.391052e-08, 
    -6.370691e-08, -6.394504e-08, -6.341912e-08, -6.314629e-08, 
    -6.307572e-08, -6.294403e-08, -6.307872e-08, -6.306777e-08, 
    -6.319667e-08, -6.315525e-08, -6.346473e-08, -6.329849e-08, 
    -6.377079e-08, -6.394317e-08, -6.443005e-08, -6.472857e-08, 
    -6.503251e-08, -6.51667e-08, -6.520754e-08, -6.522462e-08 ;

 NET_NMIN =
  8.726471e-09, 8.765218e-09, 8.757686e-09, 8.788938e-09, 8.771602e-09, 
    8.792067e-09, 8.734327e-09, 8.766755e-09, 8.746054e-09, 8.729961e-09, 
    8.849597e-09, 8.790334e-09, 8.911176e-09, 8.87337e-09, 8.968351e-09, 
    8.905293e-09, 8.981069e-09, 8.966535e-09, 9.010287e-09, 8.997753e-09, 
    9.053716e-09, 9.016073e-09, 9.082733e-09, 9.044728e-09, 9.050671e-09, 
    9.014831e-09, 8.802261e-09, 8.842217e-09, 8.799893e-09, 8.805591e-09, 
    8.803035e-09, 8.77196e-09, 8.7563e-09, 8.723512e-09, 8.729464e-09, 
    8.753547e-09, 8.808152e-09, 8.789617e-09, 8.836338e-09, 8.835283e-09, 
    8.887303e-09, 8.863848e-09, 8.951297e-09, 8.926441e-09, 8.998275e-09, 
    8.980209e-09, 8.997427e-09, 8.992206e-09, 8.997494e-09, 8.970997e-09, 
    8.982349e-09, 8.959035e-09, 8.86824e-09, 8.89492e-09, 8.815351e-09, 
    8.767515e-09, 8.735749e-09, 8.713209e-09, 8.716395e-09, 8.722469e-09, 
    8.753688e-09, 8.783045e-09, 8.805418e-09, 8.820384e-09, 8.835132e-09, 
    8.879769e-09, 8.903403e-09, 8.956322e-09, 8.946773e-09, 8.962951e-09, 
    8.978411e-09, 9.004364e-09, 9.000093e-09, 9.011528e-09, 8.962527e-09, 
    8.995091e-09, 8.941334e-09, 8.956036e-09, 8.839134e-09, 8.794618e-09, 
    8.775692e-09, 8.759133e-09, 8.718845e-09, 8.746666e-09, 8.735698e-09, 
    8.761793e-09, 8.778375e-09, 8.770175e-09, 8.820793e-09, 8.801113e-09, 
    8.904803e-09, 8.860137e-09, 8.976607e-09, 8.948733e-09, 8.983289e-09, 
    8.965657e-09, 8.99587e-09, 8.968678e-09, 9.015784e-09, 9.026041e-09, 
    9.019032e-09, 9.045961e-09, 8.96717e-09, 8.997426e-09, 8.769945e-09, 
    8.771281e-09, 8.777513e-09, 8.750122e-09, 8.748446e-09, 8.723347e-09, 
    8.745681e-09, 8.75519e-09, 8.779336e-09, 8.793618e-09, 8.807197e-09, 
    8.837051e-09, 8.870396e-09, 8.917031e-09, 8.95054e-09, 8.973003e-09, 
    8.95923e-09, 8.97139e-09, 8.957795e-09, 8.951424e-09, 9.022197e-09, 
    8.982456e-09, 9.042088e-09, 9.038788e-09, 9.011799e-09, 9.03916e-09, 
    8.772221e-09, 8.764524e-09, 8.737802e-09, 8.758715e-09, 8.720614e-09, 
    8.74194e-09, 8.754202e-09, 8.801522e-09, 8.811922e-09, 8.821563e-09, 
    8.840607e-09, 8.865048e-09, 8.907928e-09, 8.945242e-09, 8.979311e-09, 
    8.976814e-09, 8.977693e-09, 8.985303e-09, 8.966452e-09, 8.988398e-09, 
    8.992082e-09, 8.982451e-09, 9.038346e-09, 9.022377e-09, 9.038718e-09, 
    9.02832e-09, 8.767026e-09, 8.779977e-09, 8.772979e-09, 8.786139e-09, 
    8.776867e-09, 8.818095e-09, 8.830457e-09, 8.888309e-09, 8.864567e-09, 
    8.902355e-09, 8.868406e-09, 8.87442e-09, 8.903585e-09, 8.870241e-09, 
    8.943183e-09, 8.893727e-09, 8.985599e-09, 8.936202e-09, 8.988695e-09, 
    8.979163e-09, 8.994945e-09, 9.00908e-09, 9.026865e-09, 9.059679e-09, 
    9.052081e-09, 9.079526e-09, 8.799286e-09, 8.816085e-09, 8.814608e-09, 
    8.832189e-09, 8.845193e-09, 8.87338e-09, 8.918594e-09, 8.901591e-09, 
    8.932806e-09, 8.939073e-09, 8.89165e-09, 8.920765e-09, 8.82733e-09, 
    8.842423e-09, 8.833437e-09, 8.800611e-09, 8.905507e-09, 8.85167e-09, 
    8.951093e-09, 8.921923e-09, 9.007064e-09, 8.964719e-09, 9.047898e-09, 
    9.083459e-09, 9.116938e-09, 9.156059e-09, 8.825255e-09, 8.81384e-09, 
    8.834281e-09, 8.862561e-09, 8.888808e-09, 8.923702e-09, 8.927273e-09, 
    8.93381e-09, 8.950745e-09, 8.964984e-09, 8.935876e-09, 8.968553e-09, 
    8.845921e-09, 8.910181e-09, 8.809524e-09, 8.839828e-09, 8.860895e-09, 
    8.851655e-09, 8.899648e-09, 8.910961e-09, 8.956932e-09, 8.933168e-09, 
    9.074681e-09, 9.012064e-09, 9.185854e-09, 9.137278e-09, 8.809852e-09, 
    8.825217e-09, 8.878697e-09, 8.853251e-09, 8.926031e-09, 8.943949e-09, 
    8.958516e-09, 8.977136e-09, 8.979147e-09, 8.99018e-09, 8.972101e-09, 
    8.989466e-09, 8.923776e-09, 8.95313e-09, 8.872585e-09, 8.892187e-09, 
    8.883169e-09, 8.873278e-09, 8.903807e-09, 8.936333e-09, 8.937031e-09, 
    8.947461e-09, 8.976849e-09, 8.926327e-09, 9.082759e-09, 8.986139e-09, 
    8.841972e-09, 8.871569e-09, 8.875799e-09, 8.864333e-09, 8.942153e-09, 
    8.913954e-09, 8.989912e-09, 8.969382e-09, 9.003021e-09, 8.986304e-09, 
    8.983845e-09, 8.962377e-09, 8.94901e-09, 8.915246e-09, 8.887777e-09, 
    8.865997e-09, 8.871061e-09, 8.894986e-09, 8.938324e-09, 8.979328e-09, 
    8.970345e-09, 9.000464e-09, 8.920755e-09, 8.954175e-09, 8.941257e-09, 
    8.974942e-09, 8.901139e-09, 8.963978e-09, 8.885078e-09, 8.891996e-09, 
    8.913394e-09, 8.95644e-09, 8.965968e-09, 8.976137e-09, 8.969862e-09, 
    8.939425e-09, 8.934439e-09, 8.912874e-09, 8.906919e-09, 8.890489e-09, 
    8.876887e-09, 8.889314e-09, 8.902366e-09, 8.939438e-09, 8.97285e-09, 
    9.00928e-09, 9.018199e-09, 9.060765e-09, 9.026111e-09, 9.083297e-09, 
    9.034674e-09, 9.118851e-09, 8.967624e-09, 9.033246e-09, 8.914369e-09, 
    8.927174e-09, 8.950335e-09, 9.003466e-09, 8.974784e-09, 9.008328e-09, 
    8.934244e-09, 8.895811e-09, 8.88587e-09, 8.86732e-09, 8.886294e-09, 
    8.884751e-09, 8.902908e-09, 8.897073e-09, 8.94067e-09, 8.917251e-09, 
    8.983783e-09, 9.008065e-09, 9.07665e-09, 9.1187e-09, 9.161514e-09, 
    9.180416e-09, 9.18617e-09, 9.188575e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.059954e-14, 5.073669e-14, 5.071005e-14, 5.082057e-14, 5.075929e-14, 
    5.083163e-14, 5.062738e-14, 5.074212e-14, 5.066889e-14, 5.061192e-14, 
    5.103474e-14, 5.082551e-14, 5.125189e-14, 5.111869e-14, 5.145308e-14, 
    5.123114e-14, 5.149779e-14, 5.144673e-14, 5.160045e-14, 5.155644e-14, 
    5.175276e-14, 5.162077e-14, 5.185447e-14, 5.172128e-14, 5.174211e-14, 
    5.16164e-14, 5.086768e-14, 5.10087e-14, 5.085931e-14, 5.087943e-14, 
    5.087041e-14, 5.076055e-14, 5.070512e-14, 5.058908e-14, 5.061016e-14, 
    5.06954e-14, 5.088848e-14, 5.0823e-14, 5.098805e-14, 5.098433e-14, 
    5.116781e-14, 5.108512e-14, 5.139314e-14, 5.130568e-14, 5.155828e-14, 
    5.149479e-14, 5.155529e-14, 5.153695e-14, 5.155552e-14, 5.146241e-14, 
    5.150231e-14, 5.142036e-14, 5.11006e-14, 5.119464e-14, 5.091392e-14, 
    5.074477e-14, 5.06324e-14, 5.055258e-14, 5.056387e-14, 5.058537e-14, 
    5.06959e-14, 5.079976e-14, 5.087884e-14, 5.093172e-14, 5.098379e-14, 
    5.114119e-14, 5.122451e-14, 5.14108e-14, 5.137723e-14, 5.143411e-14, 
    5.148848e-14, 5.157965e-14, 5.156465e-14, 5.160479e-14, 5.143264e-14, 
    5.154707e-14, 5.13581e-14, 5.140981e-14, 5.099781e-14, 5.084067e-14, 
    5.077371e-14, 5.071517e-14, 5.057254e-14, 5.067105e-14, 5.063222e-14, 
    5.07246e-14, 5.078325e-14, 5.075425e-14, 5.093316e-14, 5.086363e-14, 
    5.122944e-14, 5.1072e-14, 5.148214e-14, 5.138413e-14, 5.150562e-14, 
    5.144365e-14, 5.154981e-14, 5.145427e-14, 5.161974e-14, 5.165573e-14, 
    5.163114e-14, 5.172563e-14, 5.144897e-14, 5.155527e-14, 5.075343e-14, 
    5.075816e-14, 5.07802e-14, 5.068327e-14, 5.067735e-14, 5.058849e-14, 
    5.066757e-14, 5.070122e-14, 5.078666e-14, 5.083714e-14, 5.088512e-14, 
    5.099056e-14, 5.110819e-14, 5.127253e-14, 5.139048e-14, 5.146948e-14, 
    5.142105e-14, 5.14638e-14, 5.141601e-14, 5.13936e-14, 5.164224e-14, 
    5.150268e-14, 5.171204e-14, 5.170047e-14, 5.160574e-14, 5.170177e-14, 
    5.076148e-14, 5.073426e-14, 5.063968e-14, 5.071371e-14, 5.057882e-14, 
    5.065432e-14, 5.069771e-14, 5.086505e-14, 5.090182e-14, 5.093587e-14, 
    5.100312e-14, 5.108935e-14, 5.124047e-14, 5.137183e-14, 5.149164e-14, 
    5.148287e-14, 5.148596e-14, 5.15127e-14, 5.144644e-14, 5.152357e-14, 
    5.15365e-14, 5.150268e-14, 5.169892e-14, 5.164289e-14, 5.170022e-14, 
    5.166375e-14, 5.074312e-14, 5.078892e-14, 5.076417e-14, 5.081069e-14, 
    5.077791e-14, 5.09236e-14, 5.096725e-14, 5.117132e-14, 5.108764e-14, 
    5.122083e-14, 5.110119e-14, 5.112239e-14, 5.122512e-14, 5.110767e-14, 
    5.136457e-14, 5.11904e-14, 5.151374e-14, 5.133997e-14, 5.152461e-14, 
    5.149113e-14, 5.154658e-14, 5.159621e-14, 5.165864e-14, 5.17737e-14, 
    5.174707e-14, 5.184326e-14, 5.085717e-14, 5.091651e-14, 5.091131e-14, 
    5.09734e-14, 5.101929e-14, 5.111874e-14, 5.127804e-14, 5.121817e-14, 
    5.132809e-14, 5.135014e-14, 5.118314e-14, 5.128568e-14, 5.095623e-14, 
    5.100949e-14, 5.09778e-14, 5.086184e-14, 5.123193e-14, 5.104212e-14, 
    5.139242e-14, 5.128977e-14, 5.158913e-14, 5.144032e-14, 5.173241e-14, 
    5.185698e-14, 5.197423e-14, 5.211096e-14, 5.094891e-14, 5.09086e-14, 
    5.098079e-14, 5.108055e-14, 5.117311e-14, 5.129603e-14, 5.130861e-14, 
    5.133162e-14, 5.139121e-14, 5.144128e-14, 5.133886e-14, 5.145384e-14, 
    5.102179e-14, 5.124841e-14, 5.089334e-14, 5.100033e-14, 5.107468e-14, 
    5.10421e-14, 5.121133e-14, 5.125118e-14, 5.141295e-14, 5.132936e-14, 
    5.182623e-14, 5.160665e-14, 5.221505e-14, 5.204533e-14, 5.089451e-14, 
    5.094879e-14, 5.113746e-14, 5.104773e-14, 5.130424e-14, 5.136729e-14, 
    5.141855e-14, 5.148399e-14, 5.149107e-14, 5.152983e-14, 5.14663e-14, 
    5.152733e-14, 5.129629e-14, 5.13996e-14, 5.111594e-14, 5.118502e-14, 
    5.115325e-14, 5.111838e-14, 5.122598e-14, 5.134047e-14, 5.134296e-14, 
    5.137964e-14, 5.148286e-14, 5.130528e-14, 5.185446e-14, 5.151552e-14, 
    5.100794e-14, 5.111231e-14, 5.112726e-14, 5.108684e-14, 5.136097e-14, 
    5.126171e-14, 5.152889e-14, 5.145675e-14, 5.157494e-14, 5.151622e-14, 
    5.150757e-14, 5.143211e-14, 5.13851e-14, 5.126625e-14, 5.116947e-14, 
    5.109271e-14, 5.111056e-14, 5.119488e-14, 5.134748e-14, 5.149169e-14, 
    5.146011e-14, 5.156596e-14, 5.128566e-14, 5.140325e-14, 5.13578e-14, 
    5.147628e-14, 5.121657e-14, 5.143764e-14, 5.115998e-14, 5.118436e-14, 
    5.125974e-14, 5.14112e-14, 5.144474e-14, 5.148047e-14, 5.145843e-14, 
    5.135136e-14, 5.133383e-14, 5.125791e-14, 5.123692e-14, 5.117906e-14, 
    5.113111e-14, 5.11749e-14, 5.122088e-14, 5.135142e-14, 5.146892e-14, 
    5.15969e-14, 5.162822e-14, 5.177745e-14, 5.165593e-14, 5.185633e-14, 
    5.168589e-14, 5.198083e-14, 5.14505e-14, 5.168095e-14, 5.126318e-14, 
    5.130827e-14, 5.138973e-14, 5.157645e-14, 5.147573e-14, 5.159354e-14, 
    5.133314e-14, 5.119777e-14, 5.116277e-14, 5.109737e-14, 5.116427e-14, 
    5.115883e-14, 5.122281e-14, 5.120226e-14, 5.135575e-14, 5.127333e-14, 
    5.150735e-14, 5.159262e-14, 5.183317e-14, 5.198036e-14, 5.213007e-14, 
    5.219608e-14, 5.221617e-14, 5.222456e-14 ;

 POT_F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POT_F_NIT =
  3.836991e-11, 3.870249e-11, 3.863771e-11, 3.890682e-11, 3.875741e-11, 
    3.893379e-11, 3.84372e-11, 3.871568e-11, 3.853778e-11, 3.839976e-11, 
    3.943183e-11, 3.891881e-11, 3.996859e-11, 3.96386e-11, 4.047033e-11, 
    3.991713e-11, 4.058237e-11, 4.045433e-11, 4.084039e-11, 4.072958e-11, 
    4.122547e-11, 4.089157e-11, 4.148381e-11, 4.11456e-11, 4.11984e-11, 
    4.088055e-11, 3.902182e-11, 3.93678e-11, 3.900135e-11, 3.905058e-11, 
    3.902848e-11, 3.876047e-11, 3.862577e-11, 3.834453e-11, 3.83955e-11, 
    3.860211e-11, 3.907269e-11, 3.891261e-11, 3.931673e-11, 3.930758e-11, 
    3.976003e-11, 3.955569e-11, 4.032031e-11, 4.010219e-11, 4.07342e-11, 
    4.057475e-11, 4.072669e-11, 4.068058e-11, 4.072728e-11, 4.049358e-11, 
    4.05936e-11, 4.038829e-11, 3.959397e-11, 3.982656e-11, 3.913497e-11, 
    3.872221e-11, 3.844937e-11, 3.825638e-11, 3.828362e-11, 3.83356e-11, 
    3.860331e-11, 3.885593e-11, 3.904903e-11, 3.917848e-11, 3.930626e-11, 
    3.969433e-11, 3.99006e-11, 4.036447e-11, 4.028056e-11, 4.042277e-11, 
    4.05589e-11, 4.078798e-11, 4.075023e-11, 4.085132e-11, 4.0419e-11, 
    4.070604e-11, 4.023275e-11, 4.03619e-11, 3.934102e-11, 3.895579e-11, 
    3.87926e-11, 3.865011e-11, 3.830458e-11, 3.854301e-11, 3.844892e-11, 
    3.867296e-11, 3.881568e-11, 3.874506e-11, 3.918202e-11, 3.901182e-11, 
    3.991283e-11, 3.952339e-11, 4.054301e-11, 4.029776e-11, 4.06019e-11, 
    4.044656e-11, 4.071292e-11, 4.047315e-11, 4.088897e-11, 4.097982e-11, 
    4.091772e-11, 4.115652e-11, 4.045985e-11, 4.072663e-11, 3.874311e-11, 
    3.875462e-11, 3.880827e-11, 3.857267e-11, 3.855828e-11, 3.83431e-11, 
    3.853453e-11, 3.86162e-11, 3.882396e-11, 3.894711e-11, 3.906438e-11, 
    3.932289e-11, 3.961266e-11, 4.001976e-11, 4.031363e-11, 4.051124e-11, 
    4.039e-11, 4.049702e-11, 4.037739e-11, 4.032137e-11, 4.094575e-11, 
    4.059452e-11, 4.112212e-11, 4.109283e-11, 4.085369e-11, 4.109611e-11, 
    3.876269e-11, 3.869646e-11, 3.846694e-11, 3.864649e-11, 3.831969e-11, 
    3.850242e-11, 3.86077e-11, 3.901535e-11, 3.910524e-11, 3.918867e-11, 
    3.935373e-11, 3.95661e-11, 3.994012e-11, 4.026708e-11, 4.056681e-11, 
    4.05448e-11, 4.055255e-11, 4.061964e-11, 4.045353e-11, 4.064693e-11, 
    4.067944e-11, 4.059447e-11, 4.108889e-11, 4.094731e-11, 4.109219e-11, 
    4.099997e-11, 3.871797e-11, 3.882948e-11, 3.87692e-11, 3.888259e-11, 
    3.880267e-11, 3.915865e-11, 3.926571e-11, 3.976877e-11, 3.956191e-11, 
    3.989141e-11, 3.959531e-11, 3.964768e-11, 3.990215e-11, 3.961127e-11, 
    4.024899e-11, 3.981602e-11, 4.062224e-11, 4.018771e-11, 4.064955e-11, 
    4.056547e-11, 4.070471e-11, 4.082962e-11, 4.098706e-11, 4.127841e-11, 
    4.121084e-11, 4.145513e-11, 3.899605e-11, 3.914126e-11, 3.912847e-11, 
    3.928073e-11, 3.939353e-11, 3.963864e-11, 4.003344e-11, 3.988473e-11, 
    4.015796e-11, 4.021293e-11, 3.97979e-11, 4.005244e-11, 3.923857e-11, 
    3.936944e-11, 3.929149e-11, 3.900742e-11, 3.991892e-11, 3.944972e-11, 
    4.031843e-11, 4.006253e-11, 4.081178e-11, 4.043823e-11, 4.117367e-11, 
    4.149019e-11, 4.178932e-11, 4.214028e-11, 3.922064e-11, 3.912182e-11, 
    3.929885e-11, 3.954447e-11, 3.977312e-11, 4.007817e-11, 4.010945e-11, 
    4.016675e-11, 4.03154e-11, 4.044062e-11, 4.018486e-11, 4.047202e-11, 
    3.939981e-11, 3.995978e-11, 3.908443e-11, 3.934691e-11, 3.952991e-11, 
    3.944959e-11, 3.98677e-11, 3.996657e-11, 4.036973e-11, 4.016106e-11, 
    4.141193e-11, 4.085599e-11, 4.240858e-11, 4.197158e-11, 3.908732e-11, 
    3.922029e-11, 3.968494e-11, 3.94635e-11, 4.009857e-11, 4.025572e-11, 
    4.038371e-11, 4.054763e-11, 4.056535e-11, 4.066266e-11, 4.050325e-11, 
    4.065635e-11, 4.007877e-11, 4.033633e-11, 3.963165e-11, 3.980254e-11, 
    3.972387e-11, 3.963766e-11, 3.990402e-11, 4.018882e-11, 4.019493e-11, 
    4.028648e-11, 4.054504e-11, 4.010107e-11, 4.148392e-11, 4.062693e-11, 
    3.936556e-11, 3.962284e-11, 3.965968e-11, 3.955986e-11, 4.023993e-11, 
    3.99928e-11, 4.066029e-11, 4.047931e-11, 4.077605e-11, 4.062845e-11, 
    4.060674e-11, 4.041764e-11, 4.030012e-11, 4.000407e-11, 3.976404e-11, 
    3.957427e-11, 3.961835e-11, 3.982696e-11, 4.020627e-11, 4.056688e-11, 
    4.048774e-11, 4.07534e-11, 4.005225e-11, 4.034545e-11, 4.023198e-11, 
    4.05282e-11, 3.988077e-11, 4.043177e-11, 3.974055e-11, 3.98009e-11, 
    3.998789e-11, 4.036544e-11, 4.044924e-11, 4.05388e-11, 4.048352e-11, 
    4.021596e-11, 4.017222e-11, 3.998331e-11, 3.993122e-11, 3.978771e-11, 
    3.966909e-11, 3.977745e-11, 3.989141e-11, 4.021604e-11, 4.050979e-11, 
    4.083134e-11, 4.091025e-11, 4.128801e-11, 4.098033e-11, 4.148869e-11, 
    4.105623e-11, 4.180639e-11, 4.046384e-11, 4.104367e-11, 3.999642e-11, 
    4.010854e-11, 4.031177e-11, 4.077998e-11, 4.052686e-11, 4.082297e-11, 
    4.01705e-11, 3.983417e-11, 3.974741e-11, 3.958579e-11, 3.97511e-11, 
    3.973764e-11, 3.989614e-11, 3.984516e-11, 4.022683e-11, 4.002158e-11, 
    4.060613e-11, 4.082057e-11, 4.142944e-11, 4.180505e-11, 4.218928e-11, 
    4.23595e-11, 4.241138e-11, 4.243308e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005835613, 0.0005835643, 0.0005835638, 0.0005835661, 0.0005835648, 
    0.0005835664, 0.000583562, 0.0005835644, 0.0005835628, 0.0005835616, 
    0.0005835679, 0.0005835663, 0.00058357, 0.00058357, 0.0005835745, 
    0.0005835724, 0.0005835755, 0.0005835744, 0.0005835778, 0.0005835769, 
    0.0005835812, 0.0005835783, 0.0005835835, 0.0005835805, 0.000583581, 
    0.0005835782, 0.0005835672, 0.0005835674, 0.000583567, 0.0005835674, 
    0.0005835672, 0.0005835649, 0.0005835636, 0.0005835611, 0.0005835615, 
    0.0005835634, 0.0005835677, 0.0005835663, 0.0005835671, 0.000583567, 
    0.000583571, 0.0005835692, 0.0005835732, 0.0005835712, 0.0005835769, 
    0.0005835755, 0.0005835768, 0.0005835764, 0.0005835768, 0.0005835747, 
    0.0005835756, 0.0005835738, 0.0005835696, 0.0005835716, 0.0005835682, 
    0.0005835644, 0.000583562, 0.0005835603, 0.0005835606, 0.000583561, 
    0.0005835634, 0.0005835657, 0.0005835675, 0.0005835659, 0.000583567, 
    0.0005835704, 0.0005835723, 0.0005835735, 0.0005835728, 0.0005835741, 
    0.0005835753, 0.0005835774, 0.000583577, 0.0005835779, 0.0005835741, 
    0.0005835766, 0.0005835724, 0.0005835735, 0.0005835671, 0.0005835666, 
    0.000583565, 0.0005835638, 0.0005835607, 0.0005835629, 0.000583562, 
    0.000583564, 0.0005835654, 0.0005835647, 0.0005835659, 0.0005835671, 
    0.0005835724, 0.0005835689, 0.0005835752, 0.000583573, 0.0005835757, 
    0.0005835743, 0.0005835767, 0.0005835746, 0.0005835783, 0.0005835791, 
    0.0005835785, 0.0005835806, 0.0005835744, 0.0005835768, 0.0005835647, 
    0.0005835648, 0.0005835653, 0.0005835631, 0.000583563, 0.0005835611, 
    0.0005835628, 0.0005835635, 0.0005835654, 0.0005835666, 0.0005835676, 
    0.0005835671, 0.0005835697, 0.0005835705, 0.0005835731, 0.0005835749, 
    0.0005835738, 0.0005835748, 0.0005835737, 0.0005835732, 0.0005835787, 
    0.0005835756, 0.0005835803, 0.0005835801, 0.000583578, 0.0005835801, 
    0.0005835649, 0.0005835643, 0.0005835622, 0.0005835638, 0.0005835608, 
    0.0005835625, 0.0005835634, 0.0005835671, 0.000583568, 0.0005835659, 
    0.0005835674, 0.0005835693, 0.0005835698, 0.0005835727, 0.0005835754, 
    0.0005835752, 0.0005835753, 0.0005835759, 0.0005835744, 0.0005835761, 
    0.0005835764, 0.0005835756, 0.0005835801, 0.0005835788, 0.0005835801, 
    0.0005835792, 0.0005835645, 0.0005835655, 0.0005835649, 0.000583566, 
    0.0005835652, 0.0005835656, 0.0005835666, 0.0005835711, 0.0005835693, 
    0.0005835722, 0.0005835696, 0.00058357, 0.0005835723, 0.0005835698, 
    0.0005835725, 0.0005835715, 0.0005835759, 0.0005835719, 0.0005835761, 
    0.0005835754, 0.0005835766, 0.0005835777, 0.0005835791, 0.0005835817, 
    0.0005835811, 0.0005835833, 0.000583567, 0.0005835683, 0.0005835682, 
    0.0005835668, 0.0005835678, 0.00058357, 0.0005835706, 0.0005835722, 
    0.0005835717, 0.0005835722, 0.0005835714, 0.0005835707, 0.0005835664, 
    0.0005835675, 0.0005835668, 0.0005835671, 0.0005835724, 0.0005835682, 
    0.0005835731, 0.0005835709, 0.0005835776, 0.0005835742, 0.0005835808, 
    0.0005835835, 0.0005835863, 0.0005835893, 0.0005835662, 0.0005835681, 
    0.000583567, 0.0005835691, 0.0005835712, 0.000583571, 0.0005835713, 
    0.0005835718, 0.0005835731, 0.0005835742, 0.0005835719, 0.0005835745, 
    0.0005835677, 0.0005835699, 0.0005835678, 0.0005835673, 0.000583569, 
    0.0005835683, 0.0005835721, 0.00058357, 0.0005835736, 0.0005835718, 
    0.0005835828, 0.0005835779, 0.0005835918, 0.0005835879, 0.0005835678, 
    0.0005835662, 0.0005835704, 0.0005835684, 0.0005835712, 0.0005835726, 
    0.0005835738, 0.0005835752, 0.0005835754, 0.0005835762, 0.0005835748, 
    0.0005835762, 0.000583571, 0.0005835733, 0.0005835699, 0.0005835714, 
    0.0005835707, 0.00058357, 0.0005835724, 0.000583572, 0.0005835721, 
    0.0005835728, 0.000583575, 0.0005835712, 0.0005835834, 0.0005835757, 
    0.0005835675, 0.0005835698, 0.0005835702, 0.0005835693, 0.0005835724, 
    0.0005835702, 0.0005835762, 0.0005835746, 0.0005835773, 0.0005835759, 
    0.0005835757, 0.0005835741, 0.000583573, 0.0005835703, 0.0005835711, 
    0.0005835694, 0.0005835698, 0.0005835717, 0.0005835721, 0.0005835753, 
    0.0005835746, 0.0005835771, 0.0005835708, 0.0005835734, 0.0005835724, 
    0.000583575, 0.0005835721, 0.000583574, 0.0005835709, 0.0005835714, 
    0.0005835702, 0.0005835735, 0.0005835744, 0.0005835751, 0.0005835746, 
    0.0005835722, 0.0005835718, 0.0005835702, 0.0005835726, 0.0005835713, 
    0.0005835703, 0.0005835712, 0.0005835723, 0.0005835723, 0.0005835749, 
    0.0005835777, 0.0005835785, 0.0005835817, 0.000583579, 0.0005835834, 
    0.0005835795, 0.0005835863, 0.0005835744, 0.0005835795, 0.0005835703, 
    0.0005835713, 0.0005835731, 0.0005835772, 0.000583575, 0.0005835776, 
    0.0005835718, 0.0005835717, 0.000583571, 0.0005835695, 0.000583571, 
    0.0005835709, 0.0005835723, 0.0005835718, 0.0005835723, 0.0005835705, 
    0.0005835757, 0.0005835776, 0.000583583, 0.0005835863, 0.0005835898, 
    0.0005835913, 0.0005835918, 0.000583592 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_NODYNLNDUSE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_R =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.24139, 81.24034, 81.24054, 81.23971, 81.24017, 81.23962, 81.24117, 
    81.24031, 81.24085, 81.24128, 81.2377, 81.23967, 81.2356, 81.23701, 
    81.23404, 81.23617, 81.23369, 81.23407, 81.23287, 81.23322, 81.23172, 
    81.23272, 81.23091, 81.23195, 81.2318, 81.23275, 81.23934, 81.2379, 
    81.2394, 81.23926, 81.23932, 81.24016, 81.2406, 81.24146, 81.24129, 
    81.24066, 81.23919, 81.23968, 81.238, 81.23803, 81.23663, 81.23726, 
    81.23449, 81.23516, 81.2332, 81.2337, 81.23323, 81.23337, 81.23323, 
    81.23396, 81.23364, 81.23428, 81.23714, 81.23643, 81.23899, 81.2403, 
    81.24113, 81.24173, 81.24165, 81.24149, 81.24065, 81.23985, 81.23925, 
    81.23843, 81.23803, 81.23687, 81.23621, 81.23436, 81.2346, 81.23418, 
    81.23375, 81.23304, 81.23315, 81.23285, 81.23418, 81.2333, 81.23475, 
    81.23436, 81.23798, 81.23954, 81.24008, 81.24051, 81.24158, 81.24084, 
    81.24113, 81.24043, 81.23998, 81.2402, 81.23842, 81.23936, 81.23617, 
    81.23737, 81.2338, 81.23456, 81.23361, 81.23409, 81.23328, 81.23401, 
    81.23273, 81.23246, 81.23264, 81.2319, 81.23405, 81.23324, 81.2402, 
    81.24017, 81.24, 81.24075, 81.24079, 81.24146, 81.24086, 81.24061, 
    81.23995, 81.23957, 81.2392, 81.23798, 81.2371, 81.23543, 81.2345, 
    81.23389, 81.23426, 81.23393, 81.23431, 81.23447, 81.23257, 81.23364, 
    81.23201, 81.2321, 81.23284, 81.23209, 81.24014, 81.24035, 81.24107, 
    81.24051, 81.24153, 81.24097, 81.24065, 81.23937, 81.23907, 81.2384, 
    81.23788, 81.23723, 81.23567, 81.23466, 81.23372, 81.23379, 81.23376, 
    81.23356, 81.23407, 81.23347, 81.23338, 81.23363, 81.23211, 81.23254, 
    81.2321, 81.23238, 81.24028, 81.23994, 81.24013, 81.23978, 81.24003, 
    81.23851, 81.23818, 81.23662, 81.23724, 81.23623, 81.23714, 81.23698, 
    81.23622, 81.23708, 81.23473, 81.23648, 81.23355, 81.23493, 81.23347, 
    81.23373, 81.23329, 81.23291, 81.23242, 81.23154, 81.23174, 81.231, 
    81.23942, 81.23898, 81.239, 81.23811, 81.23776, 81.237, 81.23537, 
    81.23624, 81.23499, 81.23482, 81.2365, 81.23532, 81.23825, 81.23785, 
    81.23808, 81.23939, 81.23615, 81.2376, 81.2345, 81.23528, 81.23297, 
    81.23413, 81.23186, 81.23091, 81.22997, 81.22892, 81.2383, 81.23902, 
    81.23805, 81.23731, 81.23659, 81.23524, 81.23514, 81.23496, 81.2345, 
    81.23411, 81.23492, 81.23401, 81.23779, 81.23561, 81.23914, 81.23793, 
    81.23735, 81.23759, 81.23628, 81.23558, 81.23434, 81.23497, 81.23116, 
    81.23285, 81.22808, 81.22942, 81.23913, 81.2383, 81.23687, 81.23755, 
    81.23517, 81.23469, 81.23428, 81.23379, 81.23373, 81.23343, 81.23392, 
    81.23344, 81.23524, 81.23444, 81.23701, 81.2365, 81.23673, 81.237, 
    81.23618, 81.23491, 81.23487, 81.2346, 81.23386, 81.23516, 81.23097, 
    81.2336, 81.23785, 81.23707, 81.23694, 81.23724, 81.23473, 81.2355, 
    81.23344, 81.23399, 81.23307, 81.23353, 81.2336, 81.23418, 81.23455, 
    81.23547, 81.23662, 81.2372, 81.23706, 81.23642, 81.23485, 81.23373, 
    81.23398, 81.23315, 81.23531, 81.23441, 81.23477, 81.23384, 81.23625, 
    81.2342, 81.23668, 81.2365, 81.23552, 81.23437, 81.23409, 81.23382, 
    81.23398, 81.23482, 81.23495, 81.23553, 81.2361, 81.23653, 81.2369, 
    81.23657, 81.23622, 81.23481, 81.2339, 81.23291, 81.23266, 81.23154, 
    81.23248, 81.23096, 81.23229, 81.22997, 81.23408, 81.23229, 81.23548, 
    81.23514, 81.23453, 81.23309, 81.23385, 81.23295, 81.23495, 81.23641, 
    81.23666, 81.23716, 81.23665, 81.23669, 81.2362, 81.23635, 81.23477, 
    81.2354, 81.2336, 81.23296, 81.23108, 81.22993, 81.22874, 81.22822, 
    81.22806, 81.228 ;

 RH2M_R =
  81.24139, 81.24034, 81.24054, 81.23971, 81.24017, 81.23962, 81.24117, 
    81.24031, 81.24085, 81.24128, 81.2377, 81.23967, 81.2356, 81.23701, 
    81.23404, 81.23617, 81.23369, 81.23407, 81.23287, 81.23322, 81.23172, 
    81.23272, 81.23091, 81.23195, 81.2318, 81.23275, 81.23934, 81.2379, 
    81.2394, 81.23926, 81.23932, 81.24016, 81.2406, 81.24146, 81.24129, 
    81.24066, 81.23919, 81.23968, 81.238, 81.23803, 81.23663, 81.23726, 
    81.23449, 81.23516, 81.2332, 81.2337, 81.23323, 81.23337, 81.23323, 
    81.23396, 81.23364, 81.23428, 81.23714, 81.23643, 81.23899, 81.2403, 
    81.24113, 81.24173, 81.24165, 81.24149, 81.24065, 81.23985, 81.23925, 
    81.23843, 81.23803, 81.23687, 81.23621, 81.23436, 81.2346, 81.23418, 
    81.23375, 81.23304, 81.23315, 81.23285, 81.23418, 81.2333, 81.23475, 
    81.23436, 81.23798, 81.23954, 81.24008, 81.24051, 81.24158, 81.24084, 
    81.24113, 81.24043, 81.23998, 81.2402, 81.23842, 81.23936, 81.23617, 
    81.23737, 81.2338, 81.23456, 81.23361, 81.23409, 81.23328, 81.23401, 
    81.23273, 81.23246, 81.23264, 81.2319, 81.23405, 81.23324, 81.2402, 
    81.24017, 81.24, 81.24075, 81.24079, 81.24146, 81.24086, 81.24061, 
    81.23995, 81.23957, 81.2392, 81.23798, 81.2371, 81.23543, 81.2345, 
    81.23389, 81.23426, 81.23393, 81.23431, 81.23447, 81.23257, 81.23364, 
    81.23201, 81.2321, 81.23284, 81.23209, 81.24014, 81.24035, 81.24107, 
    81.24051, 81.24153, 81.24097, 81.24065, 81.23937, 81.23907, 81.2384, 
    81.23788, 81.23723, 81.23567, 81.23466, 81.23372, 81.23379, 81.23376, 
    81.23356, 81.23407, 81.23347, 81.23338, 81.23363, 81.23211, 81.23254, 
    81.2321, 81.23238, 81.24028, 81.23994, 81.24013, 81.23978, 81.24003, 
    81.23851, 81.23818, 81.23662, 81.23724, 81.23623, 81.23714, 81.23698, 
    81.23622, 81.23708, 81.23473, 81.23648, 81.23355, 81.23493, 81.23347, 
    81.23373, 81.23329, 81.23291, 81.23242, 81.23154, 81.23174, 81.231, 
    81.23942, 81.23898, 81.239, 81.23811, 81.23776, 81.237, 81.23537, 
    81.23624, 81.23499, 81.23482, 81.2365, 81.23532, 81.23825, 81.23785, 
    81.23808, 81.23939, 81.23615, 81.2376, 81.2345, 81.23528, 81.23297, 
    81.23413, 81.23186, 81.23091, 81.22997, 81.22892, 81.2383, 81.23902, 
    81.23805, 81.23731, 81.23659, 81.23524, 81.23514, 81.23496, 81.2345, 
    81.23411, 81.23492, 81.23401, 81.23779, 81.23561, 81.23914, 81.23793, 
    81.23735, 81.23759, 81.23628, 81.23558, 81.23434, 81.23497, 81.23116, 
    81.23285, 81.22808, 81.22942, 81.23913, 81.2383, 81.23687, 81.23755, 
    81.23517, 81.23469, 81.23428, 81.23379, 81.23373, 81.23343, 81.23392, 
    81.23344, 81.23524, 81.23444, 81.23701, 81.2365, 81.23673, 81.237, 
    81.23618, 81.23491, 81.23487, 81.2346, 81.23386, 81.23516, 81.23097, 
    81.2336, 81.23785, 81.23707, 81.23694, 81.23724, 81.23473, 81.2355, 
    81.23344, 81.23399, 81.23307, 81.23353, 81.2336, 81.23418, 81.23455, 
    81.23547, 81.23662, 81.2372, 81.23706, 81.23642, 81.23485, 81.23373, 
    81.23398, 81.23315, 81.23531, 81.23441, 81.23477, 81.23384, 81.23625, 
    81.2342, 81.23668, 81.2365, 81.23552, 81.23437, 81.23409, 81.23382, 
    81.23398, 81.23482, 81.23495, 81.23553, 81.2361, 81.23653, 81.2369, 
    81.23657, 81.23622, 81.23481, 81.2339, 81.23291, 81.23266, 81.23154, 
    81.23248, 81.23096, 81.23229, 81.22997, 81.23408, 81.23229, 81.23548, 
    81.23514, 81.23453, 81.23309, 81.23385, 81.23295, 81.23495, 81.23641, 
    81.23666, 81.23716, 81.23665, 81.23669, 81.2362, 81.23635, 81.23477, 
    81.2354, 81.2336, 81.23296, 81.23108, 81.22993, 81.22874, 81.22822, 
    81.22806, 81.228 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RSCANOPY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004370575, 0.0004389129, 0.0004385521, 0.0004400488, 0.0004392185, 
    0.0004401984, 0.0004374334, 0.0004389862, 0.0004379949, 0.0004372241, 
    0.0004429528, 0.0004401151, 0.0004459011, 0.0004440909, 0.0004486382, 
    0.0004456192, 0.0004492469, 0.000448551, 0.0004506455, 0.0004500453, 
    0.0004527242, 0.0004509223, 0.000454113, 0.0004522938, 0.0004525783, 
    0.0004508625, 0.0004406866, 0.0004425999, 0.0004405731, 0.000440846, 
    0.0004407235, 0.0004392354, 0.0004384855, 0.0004369152, 0.0004372002, 
    0.0004383535, 0.0004409683, 0.0004400806, 0.0004423177, 0.0004422672, 
    0.0004447578, 0.0004436348, 0.0004478215, 0.0004466314, 0.0004500703, 
    0.0004492053, 0.0004500296, 0.0004497796, 0.0004500327, 0.0004487642, 
    0.0004493076, 0.0004481915, 0.0004438457, 0.000445123, 0.0004413132, 
    0.0004390225, 0.0004375012, 0.0004364218, 0.0004365743, 0.0004368652, 
    0.0004383601, 0.0004397658, 0.0004408371, 0.0004415537, 0.0004422597, 
    0.0004443971, 0.0004455285, 0.0004480619, 0.0004476047, 0.0004483792, 
    0.0004491192, 0.0004503616, 0.0004501571, 0.0004507044, 0.0004483585, 
    0.0004499175, 0.0004473439, 0.0004480477, 0.000442452, 0.0004403203, 
    0.0004394141, 0.000438621, 0.0004366916, 0.0004380239, 0.0004374986, 
    0.0004387482, 0.0004395422, 0.0004391494, 0.0004415732, 0.0004406307, 
    0.0004455954, 0.0004434569, 0.000449033, 0.0004476985, 0.0004493527, 
    0.0004485086, 0.0004499548, 0.0004486531, 0.000450908, 0.000451399, 
    0.0004510634, 0.0004523525, 0.0004485806, 0.000450029, 0.0004391387, 
    0.0004392027, 0.0004395011, 0.0004381893, 0.000438109, 0.0004369071, 
    0.0004379764, 0.0004384319, 0.0004395881, 0.0004402719, 0.000440922, 
    0.0004423515, 0.000443948, 0.0004461807, 0.0004477849, 0.0004488602, 
    0.0004482008, 0.0004487828, 0.0004481321, 0.000447827, 0.0004512149, 
    0.0004493124, 0.0004521669, 0.0004520089, 0.000450717, 0.0004520266, 
    0.0004392476, 0.000438879, 0.0004375993, 0.0004386006, 0.0004367761, 
    0.0004377973, 0.0004383844, 0.0004406503, 0.0004411482, 0.0004416099, 
    0.0004425216, 0.0004436918, 0.0004457448, 0.0004475311, 0.0004491621, 
    0.0004490425, 0.0004490845, 0.0004494488, 0.0004485463, 0.0004495968, 
    0.0004497731, 0.0004493121, 0.0004519876, 0.0004512232, 0.0004520054, 
    0.0004515076, 0.0004389987, 0.0004396188, 0.0004392836, 0.0004399138, 
    0.0004394697, 0.0004414438, 0.0004420357, 0.0004448056, 0.0004436687, 
    0.000445478, 0.0004438524, 0.0004441405, 0.0004455368, 0.0004439402, 
    0.0004474324, 0.0004450645, 0.0004494629, 0.000447098, 0.000449611, 
    0.0004491546, 0.00044991, 0.0004505867, 0.0004514379, 0.0004530087, 
    0.0004526448, 0.0004539585, 0.0004405433, 0.0004413477, 0.0004412768, 
    0.0004421186, 0.0004427412, 0.0004440908, 0.0004462555, 0.0004454414, 
    0.0004469358, 0.0004472358, 0.0004449652, 0.0004463592, 0.0004418855, 
    0.0004426081, 0.0004421778, 0.0004406059, 0.0004456284, 0.0004430506, 
    0.0004478107, 0.0004464141, 0.00045049, 0.0004484629, 0.0004524445, 
    0.0004541468, 0.0004557491, 0.0004576214, 0.0004417867, 0.00044124, 
    0.0004422187, 0.0004435728, 0.0004448293, 0.0004464999, 0.0004466708, 
    0.0004469837, 0.0004477944, 0.0004484761, 0.0004470825, 0.0004486468, 
    0.0004427755, 0.0004458522, 0.0004410326, 0.0004424837, 0.0004434923, 
    0.0004430499, 0.0004453476, 0.0004458891, 0.00044809, 0.0004469523, 
    0.0004537264, 0.0004507291, 0.0004590472, 0.0004567224, 0.000441049, 
    0.0004417846, 0.0004443452, 0.0004431268, 0.0004466113, 0.0004474691, 
    0.0004481664, 0.0004490578, 0.0004491539, 0.0004496821, 0.0004488165, 
    0.0004496479, 0.0004465029, 0.0004479082, 0.000444052, 0.0004449903, 
    0.0004445586, 0.0004440849, 0.0004455466, 0.0004471038, 0.0004471371, 
    0.0004476364, 0.0004490433, 0.0004466245, 0.0004541129, 0.0004494878, 
    0.0004425868, 0.0004440038, 0.0004442063, 0.0004436573, 0.000447383, 
    0.0004460329, 0.0004496693, 0.0004486864, 0.0004502966, 0.0004494964, 
    0.0004493786, 0.0004483509, 0.0004477109, 0.0004460944, 0.0004447791, 
    0.0004437363, 0.0004439787, 0.0004451242, 0.0004471989, 0.0004491619, 
    0.0004487319, 0.0004501736, 0.0004463576, 0.0004479576, 0.000447339, 
    0.0004489516, 0.0004454195, 0.000448428, 0.0004446504, 0.0004449816, 
    0.000446006, 0.0004480669, 0.0004485228, 0.0004490097, 0.0004487092, 
    0.000447252, 0.0004470133, 0.0004459808, 0.0004456956, 0.000444909, 
    0.0004442576, 0.0004448526, 0.0004454774, 0.0004472522, 0.0004488517, 
    0.0004505956, 0.0004510224, 0.00045306, 0.0004514011, 0.0004541384, 
    0.0004518109, 0.00045584, 0.0004486023, 0.0004517437, 0.0004460526, 
    0.0004466656, 0.0004477745, 0.0004503179, 0.0004489447, 0.0004505506, 
    0.0004470039, 0.0004451638, 0.0004446878, 0.0004437996, 0.000444708, 
    0.0004446341, 0.0004455033, 0.0004452239, 0.000447311, 0.0004461899, 
    0.0004493749, 0.0004505373, 0.0004538202, 0.0004558328, 0.0004578819, 
    0.0004587864, 0.0004590617, 0.0004591768 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.512568e-14, 3.522086e-14, 3.520237e-14, 3.527907e-14, 3.523654e-14, 
    3.528675e-14, 3.5145e-14, 3.522463e-14, 3.517381e-14, 3.513427e-14, 
    3.54277e-14, 3.52825e-14, 3.557839e-14, 3.548595e-14, 3.571801e-14, 
    3.5564e-14, 3.574904e-14, 3.57136e-14, 3.582028e-14, 3.578974e-14, 
    3.592598e-14, 3.583438e-14, 3.599656e-14, 3.590413e-14, 3.591858e-14, 
    3.583135e-14, 3.531176e-14, 3.540963e-14, 3.530596e-14, 3.531992e-14, 
    3.531366e-14, 3.523741e-14, 3.519895e-14, 3.511842e-14, 3.513305e-14, 
    3.51922e-14, 3.53262e-14, 3.528075e-14, 3.53953e-14, 3.539271e-14, 
    3.552004e-14, 3.546265e-14, 3.567641e-14, 3.561572e-14, 3.579101e-14, 
    3.574696e-14, 3.578894e-14, 3.577622e-14, 3.57891e-14, 3.572449e-14, 
    3.575218e-14, 3.56953e-14, 3.54734e-14, 3.553866e-14, 3.534385e-14, 
    3.522647e-14, 3.514849e-14, 3.509309e-14, 3.510092e-14, 3.511585e-14, 
    3.519255e-14, 3.526463e-14, 3.531951e-14, 3.53562e-14, 3.539234e-14, 
    3.550157e-14, 3.555939e-14, 3.568867e-14, 3.566538e-14, 3.570485e-14, 
    3.574258e-14, 3.580584e-14, 3.579544e-14, 3.58233e-14, 3.570382e-14, 
    3.578324e-14, 3.56521e-14, 3.568798e-14, 3.540207e-14, 3.529302e-14, 
    3.524655e-14, 3.520592e-14, 3.510694e-14, 3.51753e-14, 3.514836e-14, 
    3.521247e-14, 3.525317e-14, 3.523305e-14, 3.535721e-14, 3.530895e-14, 
    3.556281e-14, 3.545356e-14, 3.573818e-14, 3.567016e-14, 3.575447e-14, 
    3.571146e-14, 3.578514e-14, 3.571884e-14, 3.583367e-14, 3.585864e-14, 
    3.584158e-14, 3.590715e-14, 3.571516e-14, 3.578893e-14, 3.523248e-14, 
    3.523576e-14, 3.525105e-14, 3.518379e-14, 3.517968e-14, 3.511802e-14, 
    3.517289e-14, 3.519625e-14, 3.525553e-14, 3.529057e-14, 3.532387e-14, 
    3.539704e-14, 3.547867e-14, 3.559271e-14, 3.567457e-14, 3.572939e-14, 
    3.569578e-14, 3.572545e-14, 3.569228e-14, 3.567674e-14, 3.584928e-14, 
    3.575243e-14, 3.589772e-14, 3.588969e-14, 3.582395e-14, 3.58906e-14, 
    3.523806e-14, 3.521918e-14, 3.515353e-14, 3.520491e-14, 3.51113e-14, 
    3.51637e-14, 3.519381e-14, 3.530994e-14, 3.533546e-14, 3.535909e-14, 
    3.540575e-14, 3.546559e-14, 3.557047e-14, 3.566163e-14, 3.574477e-14, 
    3.573869e-14, 3.574083e-14, 3.575938e-14, 3.57134e-14, 3.576693e-14, 
    3.57759e-14, 3.575243e-14, 3.588861e-14, 3.584973e-14, 3.588952e-14, 
    3.586421e-14, 3.522532e-14, 3.52571e-14, 3.523993e-14, 3.527221e-14, 
    3.524946e-14, 3.535057e-14, 3.538086e-14, 3.552248e-14, 3.546441e-14, 
    3.555684e-14, 3.547381e-14, 3.548852e-14, 3.555981e-14, 3.547831e-14, 
    3.565658e-14, 3.553572e-14, 3.57601e-14, 3.563952e-14, 3.576765e-14, 
    3.574441e-14, 3.57829e-14, 3.581734e-14, 3.586066e-14, 3.594051e-14, 
    3.592203e-14, 3.598878e-14, 3.530447e-14, 3.534565e-14, 3.534204e-14, 
    3.538513e-14, 3.541698e-14, 3.548599e-14, 3.559654e-14, 3.555499e-14, 
    3.563127e-14, 3.564658e-14, 3.553068e-14, 3.560184e-14, 3.537321e-14, 
    3.541017e-14, 3.538818e-14, 3.530771e-14, 3.556454e-14, 3.543282e-14, 
    3.567592e-14, 3.560468e-14, 3.581242e-14, 3.570915e-14, 3.591185e-14, 
    3.59983e-14, 3.607967e-14, 3.617456e-14, 3.536814e-14, 3.534016e-14, 
    3.539026e-14, 3.545949e-14, 3.552372e-14, 3.560902e-14, 3.561776e-14, 
    3.563372e-14, 3.567508e-14, 3.570982e-14, 3.563875e-14, 3.571854e-14, 
    3.541871e-14, 3.557598e-14, 3.532957e-14, 3.540382e-14, 3.545542e-14, 
    3.54328e-14, 3.555024e-14, 3.55779e-14, 3.569016e-14, 3.563216e-14, 
    3.597696e-14, 3.582458e-14, 3.624679e-14, 3.612901e-14, 3.533038e-14, 
    3.536805e-14, 3.549898e-14, 3.543671e-14, 3.561472e-14, 3.565848e-14, 
    3.569404e-14, 3.573946e-14, 3.574437e-14, 3.577127e-14, 3.572719e-14, 
    3.576954e-14, 3.56092e-14, 3.568089e-14, 3.548405e-14, 3.553199e-14, 
    3.550994e-14, 3.548574e-14, 3.556041e-14, 3.563986e-14, 3.564159e-14, 
    3.566704e-14, 3.573868e-14, 3.561545e-14, 3.599655e-14, 3.576134e-14, 
    3.54091e-14, 3.548153e-14, 3.54919e-14, 3.546385e-14, 3.565409e-14, 
    3.558521e-14, 3.577062e-14, 3.572056e-14, 3.580258e-14, 3.576183e-14, 
    3.575583e-14, 3.570346e-14, 3.567084e-14, 3.558836e-14, 3.55212e-14, 
    3.546792e-14, 3.548032e-14, 3.553883e-14, 3.564473e-14, 3.57448e-14, 
    3.572289e-14, 3.579635e-14, 3.560183e-14, 3.568343e-14, 3.565189e-14, 
    3.573411e-14, 3.555388e-14, 3.570729e-14, 3.551461e-14, 3.553153e-14, 
    3.558384e-14, 3.568894e-14, 3.571222e-14, 3.573702e-14, 3.572173e-14, 
    3.564742e-14, 3.563525e-14, 3.558257e-14, 3.5568e-14, 3.552785e-14, 
    3.549457e-14, 3.552497e-14, 3.555687e-14, 3.564746e-14, 3.5729e-14, 
    3.581782e-14, 3.583956e-14, 3.594311e-14, 3.585878e-14, 3.599785e-14, 
    3.587957e-14, 3.608425e-14, 3.571622e-14, 3.587615e-14, 3.558623e-14, 
    3.561752e-14, 3.567405e-14, 3.580363e-14, 3.573373e-14, 3.581548e-14, 
    3.563478e-14, 3.554083e-14, 3.551655e-14, 3.547116e-14, 3.551758e-14, 
    3.551381e-14, 3.555821e-14, 3.554395e-14, 3.565047e-14, 3.559327e-14, 
    3.575567e-14, 3.581485e-14, 3.598178e-14, 3.608393e-14, 3.618782e-14, 
    3.623363e-14, 3.624757e-14, 3.625339e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.167967e-14, 1.171135e-14, 1.17052e-14, 1.173073e-14, 1.171657e-14, 
    1.173328e-14, 1.16861e-14, 1.171261e-14, 1.169569e-14, 1.168253e-14, 
    1.17802e-14, 1.173187e-14, 1.183036e-14, 1.179959e-14, 1.187683e-14, 
    1.182557e-14, 1.188716e-14, 1.187536e-14, 1.191087e-14, 1.190071e-14, 
    1.194606e-14, 1.191557e-14, 1.196955e-14, 1.193878e-14, 1.19436e-14, 
    1.191456e-14, 1.174161e-14, 1.177418e-14, 1.173968e-14, 1.174432e-14, 
    1.174224e-14, 1.171686e-14, 1.170406e-14, 1.167726e-14, 1.168213e-14, 
    1.170181e-14, 1.174641e-14, 1.173129e-14, 1.176941e-14, 1.176855e-14, 
    1.181094e-14, 1.179183e-14, 1.186299e-14, 1.184278e-14, 1.190113e-14, 
    1.188647e-14, 1.190044e-14, 1.189621e-14, 1.19005e-14, 1.187899e-14, 
    1.18882e-14, 1.186927e-14, 1.179541e-14, 1.181714e-14, 1.175229e-14, 
    1.171322e-14, 1.168726e-14, 1.166882e-14, 1.167143e-14, 1.16764e-14, 
    1.170193e-14, 1.172592e-14, 1.174419e-14, 1.17564e-14, 1.176843e-14, 
    1.180479e-14, 1.182403e-14, 1.186707e-14, 1.185931e-14, 1.187245e-14, 
    1.188501e-14, 1.190607e-14, 1.190261e-14, 1.191188e-14, 1.187211e-14, 
    1.189854e-14, 1.185489e-14, 1.186684e-14, 1.177167e-14, 1.173537e-14, 
    1.17199e-14, 1.170638e-14, 1.167344e-14, 1.169619e-14, 1.168722e-14, 
    1.170856e-14, 1.172211e-14, 1.171541e-14, 1.175674e-14, 1.174067e-14, 
    1.182517e-14, 1.178881e-14, 1.188354e-14, 1.18609e-14, 1.188897e-14, 
    1.187465e-14, 1.189918e-14, 1.187711e-14, 1.191533e-14, 1.192364e-14, 
    1.191796e-14, 1.193979e-14, 1.187588e-14, 1.190044e-14, 1.171522e-14, 
    1.171631e-14, 1.17214e-14, 1.169901e-14, 1.169764e-14, 1.167712e-14, 
    1.169539e-14, 1.170316e-14, 1.172289e-14, 1.173455e-14, 1.174564e-14, 
    1.176999e-14, 1.179716e-14, 1.183513e-14, 1.186237e-14, 1.188062e-14, 
    1.186943e-14, 1.187931e-14, 1.186827e-14, 1.186309e-14, 1.192053e-14, 
    1.188829e-14, 1.193665e-14, 1.193398e-14, 1.19121e-14, 1.193428e-14, 
    1.171708e-14, 1.171079e-14, 1.168894e-14, 1.170604e-14, 1.167488e-14, 
    1.169233e-14, 1.170235e-14, 1.1741e-14, 1.17495e-14, 1.175736e-14, 
    1.177289e-14, 1.179281e-14, 1.182772e-14, 1.185806e-14, 1.188574e-14, 
    1.188371e-14, 1.188443e-14, 1.18906e-14, 1.18753e-14, 1.189312e-14, 
    1.18961e-14, 1.188829e-14, 1.193362e-14, 1.192068e-14, 1.193392e-14, 
    1.19255e-14, 1.171284e-14, 1.172342e-14, 1.17177e-14, 1.172845e-14, 
    1.172087e-14, 1.175453e-14, 1.176461e-14, 1.181175e-14, 1.179242e-14, 
    1.182318e-14, 1.179555e-14, 1.180045e-14, 1.182417e-14, 1.179704e-14, 
    1.185639e-14, 1.181616e-14, 1.189084e-14, 1.185071e-14, 1.189336e-14, 
    1.188562e-14, 1.189843e-14, 1.190989e-14, 1.192431e-14, 1.195089e-14, 
    1.194474e-14, 1.196696e-14, 1.173918e-14, 1.175289e-14, 1.175169e-14, 
    1.176603e-14, 1.177663e-14, 1.17996e-14, 1.18364e-14, 1.182257e-14, 
    1.184796e-14, 1.185305e-14, 1.181448e-14, 1.183816e-14, 1.176206e-14, 
    1.177437e-14, 1.176705e-14, 1.174026e-14, 1.182575e-14, 1.17819e-14, 
    1.186282e-14, 1.183911e-14, 1.190826e-14, 1.187388e-14, 1.194136e-14, 
    1.197013e-14, 1.199722e-14, 1.20288e-14, 1.176037e-14, 1.175106e-14, 
    1.176774e-14, 1.179078e-14, 1.181216e-14, 1.184055e-14, 1.184346e-14, 
    1.184877e-14, 1.186254e-14, 1.187411e-14, 1.185045e-14, 1.187701e-14, 
    1.177721e-14, 1.182955e-14, 1.174754e-14, 1.177225e-14, 1.178943e-14, 
    1.17819e-14, 1.182099e-14, 1.183019e-14, 1.186756e-14, 1.184825e-14, 
    1.196303e-14, 1.191231e-14, 1.205285e-14, 1.201364e-14, 1.174781e-14, 
    1.176034e-14, 1.180393e-14, 1.17832e-14, 1.184245e-14, 1.185702e-14, 
    1.186886e-14, 1.188397e-14, 1.188561e-14, 1.189456e-14, 1.187989e-14, 
    1.189398e-14, 1.184062e-14, 1.186448e-14, 1.179895e-14, 1.181491e-14, 
    1.180757e-14, 1.179952e-14, 1.182437e-14, 1.185082e-14, 1.185139e-14, 
    1.185987e-14, 1.188371e-14, 1.184269e-14, 1.196955e-14, 1.189126e-14, 
    1.177401e-14, 1.179812e-14, 1.180157e-14, 1.179223e-14, 1.185556e-14, 
    1.183263e-14, 1.189434e-14, 1.187768e-14, 1.190498e-14, 1.189142e-14, 
    1.188942e-14, 1.187199e-14, 1.186113e-14, 1.183368e-14, 1.181132e-14, 
    1.179359e-14, 1.179771e-14, 1.181719e-14, 1.185244e-14, 1.188575e-14, 
    1.187846e-14, 1.190291e-14, 1.183816e-14, 1.186532e-14, 1.185482e-14, 
    1.188219e-14, 1.18222e-14, 1.187326e-14, 1.180913e-14, 1.181476e-14, 
    1.183217e-14, 1.186716e-14, 1.187491e-14, 1.188316e-14, 1.187807e-14, 
    1.185334e-14, 1.184929e-14, 1.183175e-14, 1.18269e-14, 1.181353e-14, 
    1.180246e-14, 1.181258e-14, 1.18232e-14, 1.185335e-14, 1.188049e-14, 
    1.191006e-14, 1.191729e-14, 1.195176e-14, 1.192369e-14, 1.196998e-14, 
    1.193061e-14, 1.199874e-14, 1.187624e-14, 1.192947e-14, 1.183297e-14, 
    1.184338e-14, 1.18622e-14, 1.190533e-14, 1.188206e-14, 1.190928e-14, 
    1.184913e-14, 1.181786e-14, 1.180977e-14, 1.179466e-14, 1.181012e-14, 
    1.180886e-14, 1.182364e-14, 1.181889e-14, 1.185435e-14, 1.183531e-14, 
    1.188937e-14, 1.190907e-14, 1.196463e-14, 1.199863e-14, 1.203322e-14, 
    1.204846e-14, 1.20531e-14, 1.205504e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.150457e-11, -8.186674e-11, -8.179634e-11, -8.208847e-11, -8.192642e-11, 
    -8.211771e-11, -8.157801e-11, -8.188111e-11, -8.168762e-11, 
    -8.153719e-11, -8.265545e-11, -8.210151e-11, -8.323106e-11, 
    -8.287768e-11, -8.37655e-11, -8.317606e-11, -8.388438e-11, -8.374853e-11, 
    -8.415749e-11, -8.404033e-11, -8.456345e-11, -8.421158e-11, 
    -8.483469e-11, -8.447942e-11, -8.453498e-11, -8.419997e-11, -8.2213e-11, 
    -8.258648e-11, -8.219087e-11, -8.224412e-11, -8.222022e-11, 
    -8.192977e-11, -8.178339e-11, -8.147691e-11, -8.153255e-11, 
    -8.175766e-11, -8.226807e-11, -8.209481e-11, -8.253152e-11, 
    -8.252166e-11, -8.300792e-11, -8.278867e-11, -8.360609e-11, 
    -8.337375e-11, -8.404522e-11, -8.387634e-11, -8.403728e-11, 
    -8.398848e-11, -8.403792e-11, -8.379024e-11, -8.389635e-11, 
    -8.367842e-11, -8.282972e-11, -8.307911e-11, -8.233535e-11, 
    -8.188821e-11, -8.15913e-11, -8.13806e-11, -8.141039e-11, -8.146717e-11, 
    -8.175897e-11, -8.203337e-11, -8.22425e-11, -8.238239e-11, -8.252025e-11, 
    -8.293749e-11, -8.31584e-11, -8.365306e-11, -8.35638e-11, -8.371503e-11, 
    -8.385953e-11, -8.410213e-11, -8.406221e-11, -8.416909e-11, 
    -8.371105e-11, -8.401545e-11, -8.351296e-11, -8.365039e-11, 
    -8.255766e-11, -8.214156e-11, -8.196466e-11, -8.180987e-11, 
    -8.143329e-11, -8.169334e-11, -8.159082e-11, -8.183473e-11, 
    -8.198973e-11, -8.191307e-11, -8.238622e-11, -8.220227e-11, 
    -8.317149e-11, -8.275398e-11, -8.384268e-11, -8.358213e-11, 
    -8.390513e-11, -8.374031e-11, -8.402273e-11, -8.376855e-11, 
    -8.420888e-11, -8.430476e-11, -8.423923e-11, -8.449096e-11, 
    -8.375446e-11, -8.403727e-11, -8.191093e-11, -8.192343e-11, 
    -8.198167e-11, -8.172563e-11, -8.170997e-11, -8.147538e-11, 
    -8.168412e-11, -8.177302e-11, -8.199872e-11, -8.213222e-11, 
    -8.225913e-11, -8.253819e-11, -8.284988e-11, -8.328579e-11, 
    -8.359901e-11, -8.380899e-11, -8.368024e-11, -8.37939e-11, -8.366684e-11, 
    -8.360728e-11, -8.426882e-11, -8.389734e-11, -8.445476e-11, 
    -8.442391e-11, -8.417163e-11, -8.442738e-11, -8.19322e-11, -8.186026e-11, 
    -8.161048e-11, -8.180596e-11, -8.144983e-11, -8.164916e-11, 
    -8.176378e-11, -8.220609e-11, -8.23033e-11, -8.239342e-11, -8.257143e-11, 
    -8.279989e-11, -8.32007e-11, -8.354949e-11, -8.386794e-11, -8.38446e-11, 
    -8.385282e-11, -8.392396e-11, -8.374774e-11, -8.395289e-11, 
    -8.398732e-11, -8.38973e-11, -8.441978e-11, -8.42705e-11, -8.442325e-11, 
    -8.432606e-11, -8.188365e-11, -8.200471e-11, -8.193929e-11, -8.20623e-11, 
    -8.197563e-11, -8.2361e-11, -8.247655e-11, -8.301731e-11, -8.279539e-11, 
    -8.314861e-11, -8.283127e-11, -8.28875e-11, -8.31601e-11, -8.284842e-11, 
    -8.353024e-11, -8.306795e-11, -8.392672e-11, -8.346499e-11, 
    -8.395566e-11, -8.386657e-11, -8.401409e-11, -8.414621e-11, 
    -8.431245e-11, -8.461919e-11, -8.454817e-11, -8.480471e-11, 
    -8.218519e-11, -8.234222e-11, -8.23284e-11, -8.249275e-11, -8.26143e-11, 
    -8.287777e-11, -8.330039e-11, -8.314147e-11, -8.343325e-11, 
    -8.349183e-11, -8.304855e-11, -8.33207e-11, -8.244733e-11, -8.25884e-11, 
    -8.250441e-11, -8.219758e-11, -8.317807e-11, -8.267483e-11, 
    -8.360419e-11, -8.333152e-11, -8.412737e-11, -8.373154e-11, 
    -8.450906e-11, -8.484147e-11, -8.515442e-11, -8.55201e-11, -8.242793e-11, 
    -8.232123e-11, -8.25123e-11, -8.277665e-11, -8.302198e-11, -8.334814e-11, 
    -8.338152e-11, -8.344263e-11, -8.360093e-11, -8.373403e-11, 
    -8.346194e-11, -8.376739e-11, -8.26211e-11, -8.322176e-11, -8.228088e-11, 
    -8.256415e-11, -8.276107e-11, -8.26747e-11, -8.312331e-11, -8.322905e-11, 
    -8.365876e-11, -8.343663e-11, -8.475941e-11, -8.417411e-11, 
    -8.579862e-11, -8.534454e-11, -8.228395e-11, -8.242757e-11, 
    -8.292746e-11, -8.268961e-11, -8.336992e-11, -8.35374e-11, -8.367357e-11, 
    -8.384762e-11, -8.386642e-11, -8.396955e-11, -8.380055e-11, 
    -8.396287e-11, -8.334884e-11, -8.362323e-11, -8.287034e-11, 
    -8.305356e-11, -8.296927e-11, -8.287682e-11, -8.316219e-11, 
    -8.346621e-11, -8.347274e-11, -8.357023e-11, -8.384494e-11, 
    -8.337269e-11, -8.483492e-11, -8.393177e-11, -8.25842e-11, -8.286084e-11, 
    -8.290038e-11, -8.279321e-11, -8.352061e-11, -8.325703e-11, 
    -8.396703e-11, -8.377513e-11, -8.408957e-11, -8.393332e-11, 
    -8.391032e-11, -8.370966e-11, -8.358472e-11, -8.326911e-11, 
    -8.301233e-11, -8.280875e-11, -8.285609e-11, -8.307973e-11, 
    -8.348482e-11, -8.386811e-11, -8.378415e-11, -8.406567e-11, 
    -8.332059e-11, -8.363299e-11, -8.351224e-11, -8.38271e-11, -8.313725e-11, 
    -8.372462e-11, -8.298712e-11, -8.305177e-11, -8.325179e-11, 
    -8.365416e-11, -8.374322e-11, -8.383828e-11, -8.377962e-11, 
    -8.349511e-11, -8.344851e-11, -8.324694e-11, -8.319127e-11, 
    -8.303769e-11, -8.291055e-11, -8.302671e-11, -8.314871e-11, 
    -8.349524e-11, -8.380755e-11, -8.414808e-11, -8.423144e-11, 
    -8.462934e-11, -8.430541e-11, -8.483995e-11, -8.438545e-11, -8.51723e-11, 
    -8.375871e-11, -8.437211e-11, -8.32609e-11, -8.33806e-11, -8.359709e-11, 
    -8.409373e-11, -8.382563e-11, -8.413919e-11, -8.344668e-11, 
    -8.308744e-11, -8.299451e-11, -8.282113e-11, -8.299848e-11, 
    -8.298406e-11, -8.315378e-11, -8.309924e-11, -8.350674e-11, 
    -8.328784e-11, -8.390975e-11, -8.413672e-11, -8.477782e-11, 
    -8.517089e-11, -8.557109e-11, -8.574778e-11, -8.580157e-11, -8.582406e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -1.964416e-12, -1.973143e-12, -1.971446e-12, -1.978486e-12, -1.974581e-12, 
    -1.97919e-12, -1.966185e-12, -1.973489e-12, -1.968826e-12, -1.965201e-12, 
    -1.992148e-12, -1.9788e-12, -2.006018e-12, -1.997503e-12, -2.018896e-12, 
    -2.004693e-12, -2.021761e-12, -2.018487e-12, -2.028342e-12, 
    -2.025519e-12, -2.038124e-12, -2.029645e-12, -2.04466e-12, -2.036099e-12, 
    -2.037438e-12, -2.029365e-12, -1.981486e-12, -1.990486e-12, 
    -1.980953e-12, -1.982236e-12, -1.98166e-12, -1.974661e-12, -1.971134e-12, 
    -1.963749e-12, -1.96509e-12, -1.970514e-12, -1.982813e-12, -1.978638e-12, 
    -1.989162e-12, -1.988924e-12, -2.000641e-12, -1.995358e-12, 
    -2.015055e-12, -2.009456e-12, -2.025636e-12, -2.021567e-12, 
    -2.025445e-12, -2.024269e-12, -2.025461e-12, -2.019492e-12, 
    -2.022049e-12, -2.016798e-12, -1.996347e-12, -2.002357e-12, 
    -1.984435e-12, -1.97366e-12, -1.966505e-12, -1.961428e-12, -1.962146e-12, 
    -1.963514e-12, -1.970546e-12, -1.977158e-12, -1.982197e-12, 
    -1.985568e-12, -1.98889e-12, -1.998944e-12, -2.004267e-12, -2.016187e-12, 
    -2.014036e-12, -2.01768e-12, -2.021162e-12, -2.027008e-12, -2.026046e-12, 
    -2.028621e-12, -2.017584e-12, -2.024919e-12, -2.012811e-12, 
    -2.016122e-12, -1.989791e-12, -1.979765e-12, -1.975502e-12, 
    -1.971772e-12, -1.962698e-12, -1.968964e-12, -1.966494e-12, 
    -1.972371e-12, -1.976106e-12, -1.974259e-12, -1.98566e-12, -1.981228e-12, 
    -2.004583e-12, -1.994522e-12, -2.020756e-12, -2.014478e-12, 
    -2.022261e-12, -2.018289e-12, -2.025095e-12, -2.01897e-12, -2.02958e-12, 
    -2.03189e-12, -2.030312e-12, -2.036377e-12, -2.01863e-12, -2.025445e-12, 
    -1.974207e-12, -1.974508e-12, -1.975912e-12, -1.969743e-12, 
    -1.969365e-12, -1.963712e-12, -1.968742e-12, -1.970884e-12, 
    -1.976323e-12, -1.97954e-12, -1.982598e-12, -1.989322e-12, -1.996833e-12, 
    -2.007337e-12, -2.014885e-12, -2.019944e-12, -2.016842e-12, 
    -2.019581e-12, -2.016519e-12, -2.015084e-12, -2.031025e-12, 
    -2.022073e-12, -2.035505e-12, -2.034762e-12, -2.028683e-12, 
    -2.034845e-12, -1.97472e-12, -1.972987e-12, -1.966968e-12, -1.971678e-12, 
    -1.963097e-12, -1.9679e-12, -1.970661e-12, -1.98132e-12, -1.983662e-12, 
    -1.985834e-12, -1.990123e-12, -1.995628e-12, -2.005287e-12, 
    -2.013691e-12, -2.021365e-12, -2.020803e-12, -2.021001e-12, 
    -2.022715e-12, -2.018469e-12, -2.023412e-12, -2.024241e-12, 
    -2.022072e-12, -2.034662e-12, -2.031065e-12, -2.034746e-12, 
    -2.032404e-12, -1.97355e-12, -1.976467e-12, -1.974891e-12, -1.977855e-12, 
    -1.975767e-12, -1.985053e-12, -1.987837e-12, -2.000868e-12, -1.99552e-12, 
    -2.004031e-12, -1.996385e-12, -1.997739e-12, -2.004308e-12, 
    -1.996798e-12, -2.013227e-12, -2.002088e-12, -2.022781e-12, 
    -2.011655e-12, -2.023479e-12, -2.021332e-12, -2.024886e-12, -2.02807e-12, 
    -2.032076e-12, -2.039467e-12, -2.037756e-12, -2.043938e-12, 
    -1.980816e-12, -1.9846e-12, -1.984267e-12, -1.988227e-12, -1.991156e-12, 
    -1.997505e-12, -2.007689e-12, -2.003859e-12, -2.01089e-12, -2.012302e-12, 
    -2.00162e-12, -2.008178e-12, -1.987133e-12, -1.990532e-12, -1.988508e-12, 
    -1.981115e-12, -2.004741e-12, -1.992615e-12, -2.015009e-12, 
    -2.008439e-12, -2.027616e-12, -2.018078e-12, -2.036813e-12, 
    -2.044823e-12, -2.052364e-12, -2.061176e-12, -1.986665e-12, 
    -1.984094e-12, -1.988698e-12, -1.995068e-12, -2.00098e-12, -2.008839e-12, 
    -2.009644e-12, -2.011116e-12, -2.014931e-12, -2.018138e-12, 
    -2.011582e-12, -2.018942e-12, -1.99132e-12, -2.005794e-12, -1.983122e-12, 
    -1.989948e-12, -1.994693e-12, -1.992612e-12, -2.003422e-12, -2.00597e-12, 
    -2.016324e-12, -2.010972e-12, -2.042846e-12, -2.028742e-12, 
    -2.067887e-12, -2.056946e-12, -1.983196e-12, -1.986657e-12, 
    -1.998703e-12, -1.992971e-12, -2.009364e-12, -2.0134e-12, -2.016681e-12, 
    -2.020875e-12, -2.021328e-12, -2.023813e-12, -2.019741e-12, 
    -2.023652e-12, -2.008856e-12, -2.015468e-12, -1.997326e-12, 
    -2.001741e-12, -1.99971e-12, -1.997482e-12, -2.004358e-12, -2.011685e-12, 
    -2.011842e-12, -2.014191e-12, -2.02081e-12, -2.009431e-12, -2.044666e-12, 
    -2.022903e-12, -1.990431e-12, -1.997097e-12, -1.99805e-12, -1.995467e-12, 
    -2.012995e-12, -2.006644e-12, -2.023752e-12, -2.019128e-12, 
    -2.026705e-12, -2.02294e-12, -2.022386e-12, -2.017551e-12, -2.01454e-12, 
    -2.006935e-12, -2.000748e-12, -1.995842e-12, -1.996983e-12, 
    -2.002372e-12, -2.012133e-12, -2.021369e-12, -2.019346e-12, 
    -2.026129e-12, -2.008176e-12, -2.015703e-12, -2.012794e-12, 
    -2.020381e-12, -2.003758e-12, -2.017911e-12, -2.00014e-12, -2.001698e-12, 
    -2.006518e-12, -2.016213e-12, -2.018359e-12, -2.02065e-12, -2.019237e-12, 
    -2.012381e-12, -2.011258e-12, -2.006401e-12, -2.005059e-12, 
    -2.001359e-12, -1.998295e-12, -2.001094e-12, -2.004034e-12, 
    -2.012384e-12, -2.01991e-12, -2.028115e-12, -2.030124e-12, -2.039712e-12, 
    -2.031906e-12, -2.044787e-12, -2.033835e-12, -2.052795e-12, 
    -2.018733e-12, -2.033513e-12, -2.006737e-12, -2.009621e-12, 
    -2.014838e-12, -2.026805e-12, -2.020345e-12, -2.027901e-12, 
    -2.011214e-12, -2.002557e-12, -2.000318e-12, -1.99614e-12, -2.000414e-12, 
    -2.000066e-12, -2.004156e-12, -2.002842e-12, -2.012661e-12, 
    -2.007386e-12, -2.022372e-12, -2.027841e-12, -2.04329e-12, -2.052761e-12, 
    -2.062405e-12, -2.066662e-12, -2.067958e-12, -2.0685e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.794188e-15, 3.80448e-15, 3.802481e-15, 3.810774e-15, 3.806176e-15, 
    3.811604e-15, 3.796277e-15, 3.804887e-15, 3.799392e-15, 3.795117e-15, 
    3.826844e-15, 3.811144e-15, 3.843139e-15, 3.833144e-15, 3.858236e-15, 
    3.841582e-15, 3.861591e-15, 3.85776e-15, 3.869295e-15, 3.865992e-15, 
    3.880725e-15, 3.870819e-15, 3.888357e-15, 3.878362e-15, 3.879925e-15, 
    3.870492e-15, 3.814309e-15, 3.82489e-15, 3.813681e-15, 3.815191e-15, 
    3.814514e-15, 3.80627e-15, 3.80211e-15, 3.793403e-15, 3.794985e-15, 
    3.801381e-15, 3.815869e-15, 3.810956e-15, 3.823341e-15, 3.823062e-15, 
    3.83683e-15, 3.830625e-15, 3.853739e-15, 3.847176e-15, 3.86613e-15, 
    3.861367e-15, 3.865906e-15, 3.86453e-15, 3.865924e-15, 3.858937e-15, 
    3.861931e-15, 3.855781e-15, 3.831786e-15, 3.838844e-15, 3.817779e-15, 
    3.805086e-15, 3.796654e-15, 3.790664e-15, 3.791511e-15, 3.793125e-15, 
    3.801418e-15, 3.809212e-15, 3.815147e-15, 3.819114e-15, 3.823022e-15, 
    3.834832e-15, 3.841084e-15, 3.855063e-15, 3.852545e-15, 3.856813e-15, 
    3.860893e-15, 3.867734e-15, 3.866609e-15, 3.869621e-15, 3.856702e-15, 
    3.865289e-15, 3.851109e-15, 3.85499e-15, 3.824073e-15, 3.812282e-15, 
    3.807257e-15, 3.802865e-15, 3.792162e-15, 3.799553e-15, 3.79664e-15, 
    3.803572e-15, 3.807973e-15, 3.805797e-15, 3.819222e-15, 3.814005e-15, 
    3.841455e-15, 3.829641e-15, 3.860417e-15, 3.853062e-15, 3.862179e-15, 
    3.857529e-15, 3.865495e-15, 3.858326e-15, 3.870743e-15, 3.873443e-15, 
    3.871597e-15, 3.878688e-15, 3.857928e-15, 3.865905e-15, 3.805736e-15, 
    3.80609e-15, 3.807745e-15, 3.800471e-15, 3.800027e-15, 3.793359e-15, 
    3.799293e-15, 3.801818e-15, 3.808229e-15, 3.812017e-15, 3.815617e-15, 
    3.823529e-15, 3.832356e-15, 3.844688e-15, 3.853539e-15, 3.859467e-15, 
    3.855833e-15, 3.859041e-15, 3.855454e-15, 3.853773e-15, 3.87243e-15, 
    3.861958e-15, 3.877669e-15, 3.8768e-15, 3.869692e-15, 3.876898e-15, 
    3.80634e-15, 3.804297e-15, 3.7972e-15, 3.802755e-15, 3.792633e-15, 
    3.798299e-15, 3.801554e-15, 3.814111e-15, 3.816871e-15, 3.819426e-15, 
    3.824471e-15, 3.830942e-15, 3.842282e-15, 3.852139e-15, 3.86113e-15, 
    3.860472e-15, 3.860704e-15, 3.86271e-15, 3.857738e-15, 3.863526e-15, 
    3.864496e-15, 3.861958e-15, 3.876684e-15, 3.87248e-15, 3.876782e-15, 
    3.874045e-15, 3.804962e-15, 3.808398e-15, 3.806541e-15, 3.810033e-15, 
    3.807572e-15, 3.818505e-15, 3.82178e-15, 3.837094e-15, 3.830815e-15, 
    3.840809e-15, 3.831831e-15, 3.833422e-15, 3.84113e-15, 3.832317e-15, 
    3.851594e-15, 3.838525e-15, 3.862788e-15, 3.849749e-15, 3.863604e-15, 
    3.861091e-15, 3.865253e-15, 3.868976e-15, 3.873661e-15, 3.882296e-15, 
    3.880297e-15, 3.887515e-15, 3.81352e-15, 3.817973e-15, 3.817583e-15, 
    3.822242e-15, 3.825686e-15, 3.833148e-15, 3.845102e-15, 3.840609e-15, 
    3.848858e-15, 3.850512e-15, 3.83798e-15, 3.845675e-15, 3.820953e-15, 
    3.82495e-15, 3.822572e-15, 3.81387e-15, 3.841641e-15, 3.827398e-15, 
    3.853685e-15, 3.845982e-15, 3.868445e-15, 3.857279e-15, 3.879197e-15, 
    3.888545e-15, 3.897344e-15, 3.907604e-15, 3.820404e-15, 3.817379e-15, 
    3.822796e-15, 3.830282e-15, 3.837228e-15, 3.846451e-15, 3.847396e-15, 
    3.849122e-15, 3.853594e-15, 3.857351e-15, 3.849666e-15, 3.858293e-15, 
    3.825872e-15, 3.842878e-15, 3.816234e-15, 3.824262e-15, 3.829842e-15, 
    3.827397e-15, 3.840095e-15, 3.843086e-15, 3.855225e-15, 3.848953e-15, 
    3.886237e-15, 3.86976e-15, 3.915415e-15, 3.902679e-15, 3.816322e-15, 
    3.820395e-15, 3.834552e-15, 3.827819e-15, 3.847068e-15, 3.851799e-15, 
    3.855645e-15, 3.860556e-15, 3.861087e-15, 3.863995e-15, 3.859229e-15, 
    3.863808e-15, 3.846471e-15, 3.854223e-15, 3.832938e-15, 3.838121e-15, 
    3.835737e-15, 3.833121e-15, 3.841195e-15, 3.849786e-15, 3.849973e-15, 
    3.852725e-15, 3.860471e-15, 3.847146e-15, 3.888356e-15, 3.862922e-15, 
    3.824834e-15, 3.832665e-15, 3.833787e-15, 3.830754e-15, 3.851325e-15, 
    3.843876e-15, 3.863925e-15, 3.858512e-15, 3.86738e-15, 3.862974e-15, 
    3.862325e-15, 3.856663e-15, 3.853136e-15, 3.844217e-15, 3.836955e-15, 
    3.831194e-15, 3.832534e-15, 3.838861e-15, 3.850312e-15, 3.861134e-15, 
    3.858764e-15, 3.866707e-15, 3.845674e-15, 3.854498e-15, 3.851087e-15, 
    3.859977e-15, 3.840488e-15, 3.857078e-15, 3.836243e-15, 3.838072e-15, 
    3.843728e-15, 3.855093e-15, 3.857611e-15, 3.860292e-15, 3.858638e-15, 
    3.850603e-15, 3.849287e-15, 3.843592e-15, 3.842016e-15, 3.837674e-15, 
    3.834076e-15, 3.837362e-15, 3.840812e-15, 3.850608e-15, 3.859425e-15, 
    3.869029e-15, 3.871379e-15, 3.882577e-15, 3.873458e-15, 3.888497e-15, 
    3.875706e-15, 3.897839e-15, 3.858043e-15, 3.875336e-15, 3.843986e-15, 
    3.84737e-15, 3.853482e-15, 3.867494e-15, 3.859936e-15, 3.868776e-15, 
    3.849236e-15, 3.839078e-15, 3.836452e-15, 3.831544e-15, 3.836564e-15, 
    3.836156e-15, 3.840957e-15, 3.839415e-15, 3.850933e-15, 3.844748e-15, 
    3.862308e-15, 3.868707e-15, 3.886758e-15, 3.897803e-15, 3.909038e-15, 
    3.913991e-15, 3.915499e-15, 3.916129e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.533392e-09, -8.571281e-09, -8.563916e-09, -8.594476e-09, -8.577524e-09, 
    -8.597535e-09, -8.541075e-09, -8.572784e-09, -8.552541e-09, 
    -8.536804e-09, -8.653791e-09, -8.595841e-09, -8.714007e-09, 
    -8.677039e-09, -8.769917e-09, -8.708254e-09, -8.782353e-09, 
    -8.768141e-09, -8.810924e-09, -8.798667e-09, -8.853391e-09, 
    -8.816582e-09, -8.881766e-09, -8.844601e-09, -8.850414e-09, 
    -8.815367e-09, -8.607504e-09, -8.646575e-09, -8.605189e-09, -8.61076e-09, 
    -8.60826e-09, -8.577874e-09, -8.56256e-09, -8.530498e-09, -8.536318e-09, 
    -8.559868e-09, -8.613265e-09, -8.59514e-09, -8.640827e-09, -8.639795e-09, 
    -8.690663e-09, -8.667727e-09, -8.75324e-09, -8.728934e-09, -8.799178e-09, 
    -8.781512e-09, -8.798349e-09, -8.793243e-09, -8.798414e-09, 
    -8.772505e-09, -8.783605e-09, -8.760806e-09, -8.672022e-09, 
    -8.698112e-09, -8.620304e-09, -8.573527e-09, -8.542465e-09, 
    -8.520423e-09, -8.523539e-09, -8.529478e-09, -8.560006e-09, 
    -8.588713e-09, -8.61059e-09, -8.625225e-09, -8.639646e-09, -8.683296e-09, 
    -8.706406e-09, -8.758154e-09, -8.748817e-09, -8.764637e-09, 
    -8.779754e-09, -8.805133e-09, -8.800956e-09, -8.812137e-09, 
    -8.764221e-09, -8.796064e-09, -8.743497e-09, -8.757874e-09, 
    -8.643561e-09, -8.60003e-09, -8.581524e-09, -8.565331e-09, -8.525935e-09, 
    -8.55314e-09, -8.542415e-09, -8.567932e-09, -8.584147e-09, -8.576127e-09, 
    -8.625626e-09, -8.606381e-09, -8.707776e-09, -8.664098e-09, -8.77799e-09, 
    -8.750733e-09, -8.784524e-09, -8.767281e-09, -8.796825e-09, 
    -8.770236e-09, -8.816299e-09, -8.826329e-09, -8.819475e-09, 
    -8.845809e-09, -8.768762e-09, -8.798348e-09, -8.575903e-09, -8.57721e-09, 
    -8.583304e-09, -8.556518e-09, -8.55488e-09, -8.530338e-09, -8.552176e-09, 
    -8.561476e-09, -8.585087e-09, -8.599053e-09, -8.61233e-09, -8.641524e-09, 
    -8.674131e-09, -8.719732e-09, -8.7525e-09, -8.774466e-09, -8.760997e-09, 
    -8.772888e-09, -8.759595e-09, -8.753365e-09, -8.82257e-09, -8.783709e-09, 
    -8.84202e-09, -8.838795e-09, -8.812403e-09, -8.839158e-09, -8.578128e-09, 
    -8.570603e-09, -8.544472e-09, -8.564921e-09, -8.527666e-09, 
    -8.548518e-09, -8.560509e-09, -8.606781e-09, -8.616951e-09, 
    -8.626379e-09, -8.645001e-09, -8.668901e-09, -8.710831e-09, 
    -8.747318e-09, -8.780633e-09, -8.778192e-09, -8.779052e-09, 
    -8.786493e-09, -8.768059e-09, -8.78952e-09, -8.793122e-09, -8.783704e-09, 
    -8.838362e-09, -8.822746e-09, -8.838725e-09, -8.828558e-09, -8.57305e-09, 
    -8.585713e-09, -8.57887e-09, -8.591739e-09, -8.582672e-09, -8.622987e-09, 
    -8.635076e-09, -8.691647e-09, -8.66843e-09, -8.705382e-09, -8.672184e-09, 
    -8.678065e-09, -8.706585e-09, -8.673978e-09, -8.745306e-09, 
    -8.696944e-09, -8.786782e-09, -8.738479e-09, -8.78981e-09, -8.780489e-09, 
    -8.795922e-09, -8.809744e-09, -8.827135e-09, -8.859223e-09, 
    -8.851793e-09, -8.87863e-09, -8.604595e-09, -8.621022e-09, -8.619577e-09, 
    -8.63677e-09, -8.649486e-09, -8.677049e-09, -8.721261e-09, -8.704635e-09, 
    -8.735159e-09, -8.741287e-09, -8.694914e-09, -8.723385e-09, 
    -8.632018e-09, -8.646777e-09, -8.63799e-09, -8.60589e-09, -8.708464e-09, 
    -8.655818e-09, -8.753041e-09, -8.724516e-09, -8.807772e-09, 
    -8.766365e-09, -8.847702e-09, -8.882476e-09, -8.915213e-09, 
    -8.953468e-09, -8.629989e-09, -8.618827e-09, -8.638815e-09, 
    -8.666469e-09, -8.692135e-09, -8.726255e-09, -8.729748e-09, 
    -8.736141e-09, -8.752701e-09, -8.766624e-09, -8.73816e-09, -8.770114e-09, 
    -8.650197e-09, -8.713035e-09, -8.614606e-09, -8.64424e-09, -8.66484e-09, 
    -8.655804e-09, -8.702735e-09, -8.713797e-09, -8.75875e-09, -8.735512e-09, 
    -8.873892e-09, -8.812662e-09, -8.982603e-09, -8.935102e-09, 
    -8.614927e-09, -8.629952e-09, -8.682247e-09, -8.657365e-09, 
    -8.728534e-09, -8.746055e-09, -8.760299e-09, -8.778507e-09, 
    -8.780474e-09, -8.791263e-09, -8.773584e-09, -8.790565e-09, 
    -8.726329e-09, -8.755032e-09, -8.676271e-09, -8.695438e-09, 
    -8.686621e-09, -8.676948e-09, -8.706802e-09, -8.738608e-09, -8.73929e-09, 
    -8.749489e-09, -8.778227e-09, -8.728823e-09, -8.881791e-09, 
    -8.787311e-09, -8.646336e-09, -8.675277e-09, -8.679414e-09, 
    -8.668202e-09, -8.744298e-09, -8.716723e-09, -8.791e-09, -8.770924e-09, 
    -8.803818e-09, -8.787472e-09, -8.785067e-09, -8.764075e-09, 
    -8.751004e-09, -8.717987e-09, -8.691126e-09, -8.669828e-09, 
    -8.674781e-09, -8.698176e-09, -8.740554e-09, -8.780651e-09, 
    -8.771867e-09, -8.801319e-09, -8.723374e-09, -8.756055e-09, 
    -8.743422e-09, -8.776361e-09, -8.704193e-09, -8.765641e-09, 
    -8.688487e-09, -8.695252e-09, -8.716176e-09, -8.758269e-09, 
    -8.767586e-09, -8.77753e-09, -8.771394e-09, -8.741631e-09, -8.736755e-09, 
    -8.715668e-09, -8.709844e-09, -8.693779e-09, -8.680478e-09, -8.69263e-09, 
    -8.705393e-09, -8.741644e-09, -8.774315e-09, -8.809939e-09, -8.81866e-09, 
    -8.860285e-09, -8.826397e-09, -8.882317e-09, -8.834771e-09, 
    -8.917084e-09, -8.769206e-09, -8.833375e-09, -8.717129e-09, 
    -8.729651e-09, -8.752299e-09, -8.804253e-09, -8.776206e-09, 
    -8.809009e-09, -8.736564e-09, -8.698983e-09, -8.689262e-09, 
    -8.671123e-09, -8.689677e-09, -8.688168e-09, -8.705922e-09, 
    -8.700217e-09, -8.742847e-09, -8.719947e-09, -8.785007e-09, 
    -8.808751e-09, -8.875817e-09, -8.916937e-09, -8.958803e-09, 
    -8.977286e-09, -8.982912e-09, -8.985264e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.012621e-10, -1.017119e-10, -1.016245e-10, -1.019872e-10, -1.01786e-10, 
    -1.020236e-10, -1.013533e-10, -1.017297e-10, -1.014894e-10, 
    -1.013026e-10, -1.026914e-10, -1.020034e-10, -1.034062e-10, 
    -1.029674e-10, -1.0407e-10, -1.033379e-10, -1.042176e-10, -1.040489e-10, 
    -1.045568e-10, -1.044113e-10, -1.05061e-10, -1.04624e-10, -1.053979e-10, 
    -1.049566e-10, -1.050256e-10, -1.046096e-10, -1.021419e-10, 
    -1.026057e-10, -1.021144e-10, -1.021805e-10, -1.021509e-10, 
    -1.017901e-10, -1.016084e-10, -1.012277e-10, -1.012968e-10, 
    -1.015764e-10, -1.022103e-10, -1.019951e-10, -1.025375e-10, 
    -1.025252e-10, -1.031291e-10, -1.028568e-10, -1.03872e-10, -1.035834e-10, 
    -1.044174e-10, -1.042076e-10, -1.044075e-10, -1.043469e-10, 
    -1.044083e-10, -1.041007e-10, -1.042325e-10, -1.039618e-10, 
    -1.029078e-10, -1.032175e-10, -1.022939e-10, -1.017385e-10, 
    -1.013698e-10, -1.011081e-10, -1.011451e-10, -1.012156e-10, -1.01578e-10, 
    -1.019188e-10, -1.021785e-10, -1.023523e-10, -1.025235e-10, 
    -1.030417e-10, -1.03316e-10, -1.039303e-10, -1.038195e-10, -1.040073e-10, 
    -1.041868e-10, -1.044881e-10, -1.044385e-10, -1.045712e-10, 
    -1.040024e-10, -1.043804e-10, -1.037563e-10, -1.03927e-10, -1.025699e-10, 
    -1.020532e-10, -1.018335e-10, -1.016413e-10, -1.011736e-10, 
    -1.014965e-10, -1.013692e-10, -1.016721e-10, -1.018646e-10, 
    -1.017694e-10, -1.02357e-10, -1.021286e-10, -1.033323e-10, -1.028137e-10, 
    -1.041658e-10, -1.038422e-10, -1.042434e-10, -1.040387e-10, 
    -1.043894e-10, -1.040738e-10, -1.046206e-10, -1.047397e-10, 
    -1.046583e-10, -1.04971e-10, -1.040563e-10, -1.044075e-10, -1.017667e-10, 
    -1.017823e-10, -1.018546e-10, -1.015366e-10, -1.015172e-10, 
    -1.012258e-10, -1.014851e-10, -1.015955e-10, -1.018758e-10, 
    -1.020416e-10, -1.021992e-10, -1.025457e-10, -1.029328e-10, 
    -1.034742e-10, -1.038632e-10, -1.04124e-10, -1.039641e-10, -1.041053e-10, 
    -1.039474e-10, -1.038735e-10, -1.046951e-10, -1.042337e-10, -1.04926e-10, 
    -1.048877e-10, -1.045744e-10, -1.04892e-10, -1.017932e-10, -1.017038e-10, 
    -1.013936e-10, -1.016364e-10, -1.011941e-10, -1.014417e-10, -1.01584e-10, 
    -1.021333e-10, -1.02254e-10, -1.02366e-10, -1.02587e-10, -1.028708e-10, 
    -1.033685e-10, -1.038017e-10, -1.041972e-10, -1.041682e-10, 
    -1.041784e-10, -1.042668e-10, -1.040479e-10, -1.043027e-10, 
    -1.043455e-10, -1.042337e-10, -1.048826e-10, -1.046972e-10, 
    -1.048869e-10, -1.047662e-10, -1.017329e-10, -1.018832e-10, -1.01802e-10, 
    -1.019547e-10, -1.018471e-10, -1.023257e-10, -1.024692e-10, 
    -1.031408e-10, -1.028652e-10, -1.033038e-10, -1.029097e-10, 
    -1.029796e-10, -1.033181e-10, -1.02931e-10, -1.037778e-10, -1.032037e-10, 
    -1.042702e-10, -1.036968e-10, -1.043061e-10, -1.041955e-10, 
    -1.043787e-10, -1.045428e-10, -1.047493e-10, -1.051302e-10, -1.05042e-10, 
    -1.053606e-10, -1.021074e-10, -1.023024e-10, -1.022852e-10, 
    -1.024893e-10, -1.026403e-10, -1.029675e-10, -1.034923e-10, -1.03295e-10, 
    -1.036573e-10, -1.037301e-10, -1.031796e-10, -1.035176e-10, 
    -1.024329e-10, -1.026081e-10, -1.025038e-10, -1.021227e-10, 
    -1.033404e-10, -1.027154e-10, -1.038696e-10, -1.03531e-10, -1.045194e-10, 
    -1.040278e-10, -1.049934e-10, -1.054063e-10, -1.057949e-10, 
    -1.062491e-10, -1.024088e-10, -1.022763e-10, -1.025136e-10, 
    -1.028419e-10, -1.031466e-10, -1.035516e-10, -1.035931e-10, -1.03669e-10, 
    -1.038656e-10, -1.040309e-10, -1.03693e-10, -1.040723e-10, -1.026487e-10, 
    -1.033947e-10, -1.022262e-10, -1.02578e-10, -1.028225e-10, -1.027153e-10, 
    -1.032724e-10, -1.034037e-10, -1.039374e-10, -1.036615e-10, 
    -1.053044e-10, -1.045774e-10, -1.06595e-10, -1.060311e-10, -1.0223e-10, 
    -1.024084e-10, -1.030292e-10, -1.027338e-10, -1.035787e-10, 
    -1.037867e-10, -1.039558e-10, -1.04172e-10, -1.041953e-10, -1.043234e-10, 
    -1.041135e-10, -1.043151e-10, -1.035525e-10, -1.038933e-10, 
    -1.029582e-10, -1.031858e-10, -1.030811e-10, -1.029663e-10, 
    -1.033207e-10, -1.036983e-10, -1.037064e-10, -1.038275e-10, 
    -1.041686e-10, -1.035821e-10, -1.053982e-10, -1.042765e-10, 
    -1.026029e-10, -1.029465e-10, -1.029956e-10, -1.028625e-10, 
    -1.037658e-10, -1.034385e-10, -1.043203e-10, -1.040819e-10, 
    -1.044725e-10, -1.042784e-10, -1.042498e-10, -1.040006e-10, 
    -1.038455e-10, -1.034535e-10, -1.031346e-10, -1.028818e-10, 
    -1.029406e-10, -1.032183e-10, -1.037214e-10, -1.041974e-10, 
    -1.040931e-10, -1.044428e-10, -1.035174e-10, -1.039054e-10, 
    -1.037554e-10, -1.041465e-10, -1.032897e-10, -1.040192e-10, 
    -1.031033e-10, -1.031836e-10, -1.03432e-10, -1.039317e-10, -1.040423e-10, 
    -1.041604e-10, -1.040875e-10, -1.037342e-10, -1.036763e-10, -1.03426e-10, 
    -1.033568e-10, -1.031661e-10, -1.030082e-10, -1.031525e-10, -1.03304e-10, 
    -1.037343e-10, -1.041222e-10, -1.045451e-10, -1.046487e-10, 
    -1.051428e-10, -1.047405e-10, -1.054044e-10, -1.048399e-10, 
    -1.058172e-10, -1.040615e-10, -1.048234e-10, -1.034433e-10, -1.03592e-10, 
    -1.038608e-10, -1.044776e-10, -1.041447e-10, -1.045341e-10, -1.03674e-10, 
    -1.032279e-10, -1.031125e-10, -1.028971e-10, -1.031174e-10, 
    -1.030995e-10, -1.033103e-10, -1.032425e-10, -1.037486e-10, 
    -1.034768e-10, -1.042491e-10, -1.04531e-10, -1.053272e-10, -1.058154e-10, 
    -1.063125e-10, -1.065319e-10, -1.065987e-10, -1.066266e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.398598e-12, -8.435918e-12, -8.428663e-12, -8.458765e-12, -8.442067e-12, 
    -8.461778e-12, -8.406165e-12, -8.437398e-12, -8.417459e-12, 
    -8.401959e-12, -8.51719e-12, -8.460109e-12, -8.576502e-12, -8.540089e-12, 
    -8.631575e-12, -8.570836e-12, -8.643824e-12, -8.629824e-12, 
    -8.671967e-12, -8.659893e-12, -8.713798e-12, -8.67754e-12, -8.741748e-12, 
    -8.70514e-12, -8.710864e-12, -8.676343e-12, -8.471598e-12, -8.510082e-12, 
    -8.469316e-12, -8.474804e-12, -8.472342e-12, -8.442412e-12, 
    -8.427327e-12, -8.395747e-12, -8.40148e-12, -8.424677e-12, -8.477272e-12, 
    -8.459418e-12, -8.504419e-12, -8.503404e-12, -8.553509e-12, 
    -8.530916e-12, -8.615147e-12, -8.591206e-12, -8.660397e-12, 
    -8.642994e-12, -8.659579e-12, -8.654551e-12, -8.659645e-12, 
    -8.634123e-12, -8.645057e-12, -8.6226e-12, -8.535147e-12, -8.560845e-12, 
    -8.484206e-12, -8.43813e-12, -8.407534e-12, -8.385823e-12, -8.388893e-12, 
    -8.394743e-12, -8.424812e-12, -8.453088e-12, -8.474637e-12, 
    -8.489052e-12, -8.503257e-12, -8.546252e-12, -8.569016e-12, 
    -8.619988e-12, -8.61079e-12, -8.626373e-12, -8.641263e-12, -8.666262e-12, 
    -8.662147e-12, -8.673161e-12, -8.625964e-12, -8.65733e-12, -8.60555e-12, 
    -8.619712e-12, -8.507113e-12, -8.464235e-12, -8.446007e-12, 
    -8.430057e-12, -8.391252e-12, -8.418049e-12, -8.407485e-12, 
    -8.432619e-12, -8.448591e-12, -8.440692e-12, -8.489447e-12, 
    -8.470491e-12, -8.570364e-12, -8.527342e-12, -8.639526e-12, 
    -8.612678e-12, -8.645962e-12, -8.628978e-12, -8.658079e-12, 
    -8.631889e-12, -8.677261e-12, -8.687141e-12, -8.68039e-12, -8.706328e-12, 
    -8.630437e-12, -8.659578e-12, -8.440471e-12, -8.441758e-12, -8.44776e-12, 
    -8.421377e-12, -8.419763e-12, -8.39559e-12, -8.417099e-12, -8.42626e-12, 
    -8.449517e-12, -8.463273e-12, -8.476351e-12, -8.505106e-12, 
    -8.537224e-12, -8.582142e-12, -8.614418e-12, -8.636055e-12, 
    -8.622788e-12, -8.6345e-12, -8.621407e-12, -8.61527e-12, -8.683439e-12, 
    -8.645159e-12, -8.702598e-12, -8.69942e-12, -8.673423e-12, -8.699777e-12, 
    -8.442662e-12, -8.43525e-12, -8.409511e-12, -8.429654e-12, -8.392957e-12, 
    -8.413496e-12, -8.425307e-12, -8.470885e-12, -8.480903e-12, 
    -8.490189e-12, -8.508532e-12, -8.532073e-12, -8.573374e-12, 
    -8.609315e-12, -8.64213e-12, -8.639725e-12, -8.640572e-12, -8.647902e-12, 
    -8.629744e-12, -8.650883e-12, -8.65443e-12, -8.645155e-12, -8.698993e-12, 
    -8.683611e-12, -8.699351e-12, -8.689337e-12, -8.437659e-12, 
    -8.450134e-12, -8.443393e-12, -8.456068e-12, -8.447138e-12, 
    -8.486848e-12, -8.498755e-12, -8.554477e-12, -8.531609e-12, 
    -8.568007e-12, -8.535306e-12, -8.5411e-12, -8.569191e-12, -8.537074e-12, 
    -8.607332e-12, -8.559695e-12, -8.648186e-12, -8.600608e-12, 
    -8.651168e-12, -8.641988e-12, -8.65719e-12, -8.670804e-12, -8.687934e-12, 
    -8.719542e-12, -8.712223e-12, -8.738659e-12, -8.468732e-12, 
    -8.484912e-12, -8.483489e-12, -8.500423e-12, -8.512949e-12, 
    -8.540098e-12, -8.583647e-12, -8.567271e-12, -8.597337e-12, 
    -8.603373e-12, -8.557695e-12, -8.585739e-12, -8.495743e-12, -8.51028e-12, 
    -8.501626e-12, -8.470008e-12, -8.571042e-12, -8.519186e-12, 
    -8.614952e-12, -8.586854e-12, -8.668863e-12, -8.628075e-12, 
    -8.708194e-12, -8.742447e-12, -8.774695e-12, -8.812376e-12, 
    -8.493745e-12, -8.48275e-12, -8.502438e-12, -8.529678e-12, -8.554958e-12, 
    -8.588567e-12, -8.592007e-12, -8.598303e-12, -8.614616e-12, 
    -8.628331e-12, -8.600293e-12, -8.631769e-12, -8.51365e-12, -8.575545e-12, 
    -8.478592e-12, -8.507781e-12, -8.528072e-12, -8.519172e-12, 
    -8.565399e-12, -8.576295e-12, -8.620575e-12, -8.597685e-12, 
    -8.733991e-12, -8.673678e-12, -8.841075e-12, -8.794286e-12, 
    -8.478909e-12, -8.493707e-12, -8.545219e-12, -8.520709e-12, 
    -8.590812e-12, -8.608069e-12, -8.6221e-12, -8.640036e-12, -8.641973e-12, 
    -8.652599e-12, -8.635185e-12, -8.651912e-12, -8.588639e-12, 
    -8.616913e-12, -8.539332e-12, -8.558212e-12, -8.549527e-12, 
    -8.539999e-12, -8.569406e-12, -8.600734e-12, -8.601406e-12, 
    -8.611452e-12, -8.639759e-12, -8.591097e-12, -8.741772e-12, 
    -8.648708e-12, -8.509846e-12, -8.538353e-12, -8.542428e-12, 
    -8.531384e-12, -8.606339e-12, -8.579178e-12, -8.652341e-12, 
    -8.632566e-12, -8.664967e-12, -8.648866e-12, -8.646498e-12, 
    -8.625819e-12, -8.612945e-12, -8.580423e-12, -8.553964e-12, 
    -8.532987e-12, -8.537864e-12, -8.560909e-12, -8.602652e-12, 
    -8.642147e-12, -8.633495e-12, -8.662505e-12, -8.585728e-12, 
    -8.617919e-12, -8.605477e-12, -8.637922e-12, -8.566836e-12, 
    -8.627362e-12, -8.551365e-12, -8.558028e-12, -8.57864e-12, -8.620101e-12, 
    -8.629278e-12, -8.639073e-12, -8.633029e-12, -8.603711e-12, -8.59891e-12, 
    -8.578138e-12, -8.572402e-12, -8.556577e-12, -8.543476e-12, 
    -8.555446e-12, -8.568017e-12, -8.603725e-12, -8.635907e-12, 
    -8.670997e-12, -8.679587e-12, -8.720588e-12, -8.687208e-12, 
    -8.742291e-12, -8.695456e-12, -8.776537e-12, -8.630874e-12, 
    -8.694081e-12, -8.579578e-12, -8.591912e-12, -8.61422e-12, -8.665396e-12, 
    -8.637769e-12, -8.67008e-12, -8.598722e-12, -8.561703e-12, -8.552129e-12, 
    -8.534262e-12, -8.552537e-12, -8.55105e-12, -8.568539e-12, -8.562919e-12, 
    -8.60491e-12, -8.582354e-12, -8.646438e-12, -8.669826e-12, -8.735888e-12, 
    -8.776391e-12, -8.817631e-12, -8.835837e-12, -8.841379e-12, -8.843697e-12 ;

 SMIN_NH4 =
  0.0004358414, 0.0004376863, 0.0004373275, 0.0004388156, 0.0004379901, 
    0.0004389644, 0.0004362151, 0.0004377591, 0.0004367734, 0.000436007, 
    0.000441703, 0.0004388816, 0.0004446343, 0.0004428346, 0.0004473554, 
    0.0004443541, 0.0004479607, 0.0004472688, 0.000449351, 0.0004487544, 
    0.0004514176, 0.0004496262, 0.0004527982, 0.0004509897, 0.0004512725, 
    0.0004495668, 0.0004394498, 0.0004413521, 0.000439337, 0.0004396083, 
    0.0004394865, 0.0004380069, 0.0004372612, 0.0004356999, 0.0004359833, 
    0.00043713, 0.0004397299, 0.0004388473, 0.0004410715, 0.0004410213, 
    0.0004434976, 0.000442381, 0.0004465435, 0.0004453603, 0.0004487793, 
    0.0004479193, 0.0004487387, 0.0004484902, 0.0004487418, 0.0004474808, 
    0.0004480209, 0.0004469113, 0.0004425908, 0.0004438607, 0.0004400729, 
    0.0004377952, 0.0004362826, 0.0004352093, 0.0004353609, 0.0004356502, 
    0.0004371366, 0.0004385343, 0.0004395995, 0.0004403119, 0.0004410139, 
    0.000443139, 0.0004442639, 0.0004467826, 0.000446328, 0.000447098, 
    0.0004478337, 0.0004490688, 0.0004488655, 0.0004494096, 0.0004470774, 
    0.0004486273, 0.0004460687, 0.0004467684, 0.0004412051, 0.0004390856, 
    0.0004381845, 0.000437396, 0.0004354775, 0.0004368023, 0.00043628, 
    0.0004375224, 0.0004383119, 0.0004379214, 0.0004403313, 0.0004393943, 
    0.0004443304, 0.0004422042, 0.000447748, 0.0004464212, 0.0004480658, 
    0.0004472266, 0.0004486644, 0.0004473703, 0.000449612, 0.0004501002, 
    0.0004497665, 0.000451048, 0.0004472982, 0.0004487382, 0.0004379107, 
    0.0004379744, 0.0004382711, 0.0004369667, 0.0004368869, 0.0004356918, 
    0.0004367551, 0.000437208, 0.0004383576, 0.0004390375, 0.0004396838, 
    0.0004411052, 0.0004426925, 0.0004449122, 0.0004465072, 0.0004475762, 
    0.0004469206, 0.0004474993, 0.0004468523, 0.0004465489, 0.0004499171, 
    0.0004480258, 0.0004508635, 0.0004507065, 0.0004494221, 0.000450724, 
    0.000438019, 0.0004376525, 0.0004363801, 0.0004373757, 0.0004355615, 
    0.000436577, 0.0004371608, 0.0004394137, 0.0004399088, 0.0004403678, 
    0.0004412743, 0.0004424378, 0.0004444789, 0.0004462549, 0.0004478763, 
    0.0004477574, 0.0004477992, 0.0004481613, 0.0004472641, 0.0004483085, 
    0.0004484837, 0.0004480254, 0.0004506853, 0.0004499254, 0.0004507029, 
    0.0004502081, 0.0004377716, 0.0004383881, 0.0004380548, 0.0004386814, 
    0.0004382399, 0.0004402027, 0.0004407912, 0.0004435451, 0.0004424148, 
    0.0004442137, 0.0004425975, 0.0004428838, 0.0004442721, 0.0004426847, 
    0.0004461567, 0.0004438026, 0.0004481753, 0.0004458243, 0.0004483226, 
    0.0004478688, 0.0004486199, 0.0004492926, 0.0004501388, 0.0004517003, 
    0.0004513386, 0.0004526446, 0.0004393074, 0.0004401071, 0.0004400367, 
    0.0004408737, 0.0004414927, 0.0004428345, 0.0004449866, 0.0004441772, 
    0.000445663, 0.0004459613, 0.0004437038, 0.0004450897, 0.0004406419, 
    0.0004413603, 0.0004409325, 0.0004393696, 0.0004443632, 0.0004418003, 
    0.0004465329, 0.0004451443, 0.0004491965, 0.0004471812, 0.0004511395, 
    0.0004528317, 0.0004544245, 0.0004562857, 0.0004405436, 0.00044, 
    0.0004409731, 0.0004423195, 0.0004435687, 0.0004452297, 0.0004453996, 
    0.0004457106, 0.0004465166, 0.0004471943, 0.0004458088, 0.0004473641, 
    0.0004415268, 0.0004445856, 0.0004397938, 0.0004412366, 0.0004422394, 
    0.0004417995, 0.000444084, 0.0004446224, 0.0004468104, 0.0004456794, 
    0.0004524139, 0.0004494342, 0.000457703, 0.0004553921, 0.0004398101, 
    0.0004405415, 0.0004430874, 0.000441876, 0.0004453404, 0.0004461932, 
    0.0004468864, 0.0004477726, 0.0004478682, 0.0004483933, 0.0004475328, 
    0.0004483592, 0.0004452326, 0.0004466298, 0.0004427958, 0.0004437288, 
    0.0004432996, 0.0004428286, 0.0004442818, 0.00044583, 0.0004458631, 
    0.0004463595, 0.0004477582, 0.0004453534, 0.0004527981, 0.0004482001, 
    0.0004413391, 0.000442748, 0.0004429493, 0.0004424035, 0.0004461076, 
    0.0004447654, 0.0004483805, 0.0004474034, 0.0004490043, 0.0004482087, 
    0.0004480915, 0.0004470698, 0.0004464336, 0.0004448265, 0.0004435188, 
    0.000442482, 0.000442723, 0.0004438619, 0.0004459246, 0.0004478762, 
    0.0004474486, 0.0004488819, 0.0004450881, 0.0004466788, 0.0004460638, 
    0.0004476671, 0.0004441555, 0.0004471465, 0.0004433909, 0.0004437201, 
    0.0004447386, 0.0004467875, 0.0004472408, 0.0004477248, 0.000447426, 
    0.0004459774, 0.00044574, 0.0004447135, 0.00044443, 0.0004436479, 
    0.0004430003, 0.0004435919, 0.000444213, 0.0004459776, 0.0004475677, 
    0.0004493014, 0.0004497258, 0.0004517514, 0.0004501023, 0.0004528234, 
    0.0004505097, 0.000454515, 0.0004473198, 0.0004504429, 0.000444785, 
    0.0004453944, 0.0004464968, 0.0004490253, 0.0004476602, 0.0004492567, 
    0.0004457307, 0.0004439012, 0.000443428, 0.000442545, 0.0004434481, 
    0.0004433746, 0.0004442388, 0.000443961, 0.000446036, 0.0004449214, 
    0.0004480879, 0.0004492435, 0.0004525071, 0.0004545078, 0.0004565447, 
    0.0004574438, 0.0004577175, 0.0004578319 ;

 SMIN_NH4_vr =
  0.002870855, 0.002875837, 0.002874863, 0.002878877, 0.002876648, 
    0.00287927, 0.002871851, 0.002876013, 0.002873352, 0.002871278, 
    0.002886628, 0.002879032, 0.002894514, 0.002889671, 0.002901813, 
    0.002893751, 0.002903434, 0.002901574, 0.002907157, 0.002905554, 
    0.00291268, 0.002907887, 0.00291637, 0.002911532, 0.002912284, 
    0.002907713, 0.002880585, 0.002885706, 0.002880275, 0.002881007, 
    0.002880675, 0.00287668, 0.002874665, 0.002870447, 0.002871208, 
    0.002874304, 0.002881313, 0.00287893, 0.00288492, 0.002884786, 
    0.002891443, 0.00288844, 0.002899624, 0.002896443, 0.002905617, 
    0.002903306, 0.002905502, 0.002904831, 0.002905502, 0.00290212, 
    0.002903563, 0.002900586, 0.002889039, 0.00289245, 0.002882253, 
    0.002876104, 0.00287202, 0.002869122, 0.002869525, 0.002870306, 
    0.002874316, 0.002878084, 0.002880955, 0.00288287, 0.002884757, 
    0.002890473, 0.002893496, 0.002900258, 0.002899038, 0.002901099, 
    0.002903073, 0.00290638, 0.002905834, 0.002907287, 0.00290103, 
    0.002905187, 0.002898316, 0.002900195, 0.002885295, 0.002879586, 
    0.002877151, 0.002875021, 0.002869837, 0.002873415, 0.002872001, 
    0.002875352, 0.00287748, 0.002876423, 0.002882919, 0.002880389, 
    0.00289367, 0.002887953, 0.002902847, 0.002899282, 0.002903691, 
    0.00290144, 0.00290529, 0.00290182, 0.002907824, 0.002909132, 
    0.002908232, 0.002911665, 0.002901608, 0.00290547, 0.002876411, 
    0.002876583, 0.00287738, 0.002873854, 0.002873638, 0.002870406, 
    0.002873274, 0.002874497, 0.002877596, 0.002879424, 0.002881163, 
    0.002884993, 0.002889261, 0.002895225, 0.002899509, 0.002902374, 
    0.002900613, 0.002902162, 0.002900424, 0.002899605, 0.002908632, 
    0.002903564, 0.002911163, 0.002910743, 0.002907297, 0.002910781, 
    0.002876698, 0.002875705, 0.002872268, 0.002874952, 0.002870049, 
    0.002872791, 0.002874363, 0.002880436, 0.002881768, 0.002883005, 
    0.002885443, 0.00288857, 0.002894057, 0.002898824, 0.002903176, 
    0.002902852, 0.002902963, 0.002903929, 0.002901521, 0.002904318, 
    0.002904783, 0.002903556, 0.002910678, 0.002908643, 0.002910722, 
    0.002909392, 0.002876023, 0.002877681, 0.002876778, 0.002878468, 
    0.002877271, 0.002882562, 0.002884143, 0.002891551, 0.002888508, 
    0.002893346, 0.002888994, 0.002889764, 0.00289349, 0.002889221, 
    0.00289855, 0.002892219, 0.002903963, 0.002897645, 0.002904352, 
    0.002903131, 0.002905142, 0.002906945, 0.002909206, 0.002913386, 
    0.002912412, 0.002915907, 0.002880157, 0.002882306, 0.002882117, 
    0.002884367, 0.002886029, 0.002889642, 0.002895424, 0.002893245, 
    0.002897234, 0.002898035, 0.002891963, 0.002895687, 0.002883717, 
    0.002885646, 0.002884494, 0.002880278, 0.002893718, 0.002886819, 
    0.002899542, 0.002895809, 0.002906678, 0.002901273, 0.002911877, 
    0.002916402, 0.002920659, 0.00292562, 0.00288348, 0.002882011, 
    0.002884629, 0.002888252, 0.002891608, 0.002896073, 0.002896527, 
    0.002897357, 0.002899518, 0.002901338, 0.002897612, 0.002901785, 
    0.002886088, 0.002894316, 0.002881416, 0.002885301, 0.002887996, 
    0.002886813, 0.002892956, 0.002894399, 0.00290027, 0.002897235, 
    0.002915276, 0.0029073, 0.002929396, 0.002923231, 0.002881496, 
    0.002883462, 0.00289031, 0.002887052, 0.002896363, 0.002898654, 
    0.002900509, 0.002902886, 0.002903137, 0.002904545, 0.002902231, 
    0.002904449, 0.002896049, 0.002899803, 0.002889495, 0.002891999, 
    0.002890845, 0.002889573, 0.002893477, 0.002897636, 0.002897723, 
    0.00289905, 0.002902796, 0.002896343, 0.002916288, 0.002903971, 
    0.002885608, 0.002889392, 0.002889932, 0.002888465, 0.002898415, 
    0.00289481, 0.002904511, 0.002901886, 0.002906175, 0.002904043, 
    0.002903722, 0.002900982, 0.002899267, 0.00289495, 0.002891428, 
    0.002888641, 0.002889283, 0.002892346, 0.002897881, 0.002903121, 
    0.002901969, 0.00290581, 0.002895624, 0.002899896, 0.002898238, 
    0.002902543, 0.002893174, 0.002901202, 0.002891115, 0.002891996, 
    0.002894729, 0.002900231, 0.002901444, 0.002902742, 0.002901935, 
    0.002898045, 0.002897405, 0.002894643, 0.002893876, 0.002891775, 
    0.002890027, 0.002891618, 0.002893281, 0.002898023, 0.002902287, 
    0.002906932, 0.002908068, 0.002913482, 0.002909067, 0.002916341, 
    0.002910147, 0.002920858, 0.002901661, 0.002910033, 0.002894855, 
    0.002896488, 0.002899445, 0.002906223, 0.002902561, 0.00290684, 
    0.002897378, 0.002892455, 0.002891181, 0.002888806, 0.002891229, 
    0.002891032, 0.002893352, 0.002892601, 0.002898172, 0.002895179, 
    0.002903672, 0.00290677, 0.002915504, 0.002920846, 0.002926285, 
    0.002928678, 0.002929407, 0.002929708,
  0.001603353, 0.001609473, 0.001608284, 0.001613217, 0.001610482, 
    0.00161371, 0.001604595, 0.001609716, 0.001606448, 0.001603905, 
    0.001622778, 0.001613437, 0.001632473, 0.001626524, 0.001641459, 
    0.001631547, 0.001643457, 0.001641175, 0.001648043, 0.001646076, 
    0.00165485, 0.001648951, 0.001659396, 0.001653443, 0.001654374, 
    0.001648756, 0.001615319, 0.001621615, 0.001614945, 0.001615844, 
    0.001615441, 0.001610538, 0.001608064, 0.001602886, 0.001603827, 
    0.001607631, 0.001616248, 0.001613325, 0.001620692, 0.001620526, 
    0.001628718, 0.001625025, 0.001638781, 0.001634875, 0.001646158, 
    0.001643322, 0.001646025, 0.001645206, 0.001646036, 0.001641876, 
    0.001643658, 0.001639997, 0.001625717, 0.001629916, 0.001617383, 
    0.001609834, 0.00160482, 0.001601258, 0.001601761, 0.001602721, 
    0.001607653, 0.001612287, 0.001615817, 0.001618177, 0.001620502, 
    0.00162753, 0.00163125, 0.00163957, 0.001638071, 0.001640612, 0.00164304, 
    0.001647113, 0.001646443, 0.001648237, 0.001640546, 0.001645658, 
    0.001637216, 0.001639526, 0.001621129, 0.001614114, 0.001611126, 
    0.001608513, 0.001602149, 0.001606544, 0.001604811, 0.001608933, 
    0.001611551, 0.001610256, 0.001618242, 0.001615138, 0.001631471, 
    0.00162444, 0.001642757, 0.001638378, 0.001643806, 0.001641037, 
    0.00164578, 0.001641512, 0.001648905, 0.001650513, 0.001649414, 
    0.001653637, 0.001641275, 0.001646025, 0.00161022, 0.001610431, 
    0.001611415, 0.001607089, 0.001606825, 0.00160286, 0.001606389, 
    0.00160789, 0.001611703, 0.001613956, 0.001616098, 0.001620804, 
    0.001626056, 0.001633394, 0.001638662, 0.001642191, 0.001640028, 
    0.001641938, 0.001639802, 0.001638802, 0.00164991, 0.001643675, 
    0.00165303, 0.001652512, 0.00164828, 0.001652571, 0.001610579, 
    0.001609365, 0.001605144, 0.001608447, 0.001602428, 0.001605797, 
    0.001607734, 0.001615202, 0.001616843, 0.001618363, 0.001621364, 
    0.001625214, 0.001631963, 0.001637829, 0.001643182, 0.00164279, 
    0.001642928, 0.001644122, 0.001641162, 0.001644608, 0.001645186, 
    0.001643674, 0.001652443, 0.001649939, 0.001652501, 0.001650871, 
    0.00160976, 0.001611804, 0.001610699, 0.001612776, 0.001611312, 
    0.001617815, 0.001619764, 0.001628875, 0.001625138, 0.001631086, 
    0.001625743, 0.00162669, 0.001631278, 0.001626032, 0.001637505, 
    0.001629727, 0.001644169, 0.001636407, 0.001644655, 0.001643158, 
    0.001645636, 0.001647853, 0.001650643, 0.001655786, 0.001654595, 
    0.001658894, 0.00161485, 0.001617499, 0.001617266, 0.001620038, 
    0.001622087, 0.001626527, 0.00163364, 0.001630966, 0.001635876, 
    0.00163686, 0.001629402, 0.001633982, 0.001619271, 0.001621649, 
    0.001620234, 0.001615059, 0.001631581, 0.001623106, 0.001638749, 
    0.001634164, 0.001647537, 0.001640889, 0.00165394, 0.001659509, 
    0.00166475, 0.001670864, 0.001618945, 0.001617145, 0.001620368, 
    0.001624822, 0.001628955, 0.001634444, 0.001635006, 0.001636033, 
    0.001638695, 0.001640932, 0.001636357, 0.001641492, 0.001622199, 
    0.001632317, 0.001616464, 0.00162124, 0.00162456, 0.001623105, 
    0.001630661, 0.00163244, 0.001639666, 0.001635932, 0.001658134, 
    0.00164832, 0.001675518, 0.001667929, 0.001616516, 0.001618939, 
    0.001627363, 0.001623356, 0.00163481, 0.001637627, 0.001639916, 
    0.00164284, 0.001643156, 0.001644887, 0.001642049, 0.001644776, 
    0.001634455, 0.001639069, 0.001626401, 0.001629486, 0.001628068, 
    0.001626511, 0.001631315, 0.001636429, 0.001636539, 0.001638178, 
    0.001642791, 0.001634857, 0.001659397, 0.00164425, 0.00162158, 
    0.00162624, 0.001626907, 0.001625102, 0.001637344, 0.001632911, 
    0.001644845, 0.001641622, 0.001646903, 0.001644279, 0.001643893, 
    0.001640522, 0.001638422, 0.001633114, 0.001628792, 0.001625364, 
    0.001626162, 0.001629927, 0.001636742, 0.001643184, 0.001641773, 
    0.001646502, 0.001633981, 0.001639233, 0.001637203, 0.001642495, 
    0.001630895, 0.00164077, 0.001628368, 0.001629457, 0.001632823, 
    0.001639588, 0.001641086, 0.001642683, 0.001641698, 0.001636915, 
    0.001636132, 0.001632741, 0.001631804, 0.00162922, 0.001627079, 
    0.001629035, 0.001631088, 0.001636918, 0.001642166, 0.001647885, 
    0.001649284, 0.001655954, 0.001650523, 0.001659481, 0.001651863, 
    0.001665046, 0.001641344, 0.001651641, 0.001632976, 0.00163499, 
    0.001638629, 0.001646971, 0.00164247, 0.001647735, 0.001636101, 
    0.001630056, 0.001628493, 0.001625572, 0.001628559, 0.001628317, 
    0.001631174, 0.001630256, 0.001637111, 0.00163343, 0.001643883, 
    0.001647693, 0.001658444, 0.001665024, 0.001671718, 0.00167467, 
    0.001675568, 0.001675944,
  0.001504877, 0.001511566, 0.001510266, 0.001515659, 0.001512668, 
    0.001516199, 0.001506234, 0.001511832, 0.001508259, 0.00150548, 
    0.001526117, 0.0015159, 0.001536723, 0.001530214, 0.001546559, 
    0.00153571, 0.001548745, 0.001546247, 0.001553767, 0.001551613, 
    0.001561224, 0.00155476, 0.001566204, 0.001559681, 0.001560701, 
    0.001554547, 0.001517957, 0.001524845, 0.001517549, 0.001518531, 
    0.001518091, 0.00151273, 0.001510027, 0.001504366, 0.001505394, 
    0.001509552, 0.001518973, 0.001515777, 0.001523833, 0.001523651, 
    0.001532613, 0.001528573, 0.001543626, 0.00153935, 0.001551703, 
    0.001548597, 0.001551557, 0.00155066, 0.001551568, 0.001547014, 
    0.001548965, 0.001544957, 0.00152933, 0.001533924, 0.001520215, 
    0.001511962, 0.001506479, 0.001502586, 0.001503137, 0.001504186, 
    0.001509576, 0.001514643, 0.001518502, 0.001521083, 0.001523625, 
    0.001531315, 0.001535385, 0.00154449, 0.001542848, 0.00154563, 
    0.001548289, 0.001552749, 0.001552015, 0.001553979, 0.001545558, 
    0.001551155, 0.001541913, 0.001544441, 0.001524313, 0.001516639, 
    0.001513373, 0.001510516, 0.00150356, 0.001508364, 0.00150647, 
    0.001510976, 0.001513837, 0.001512422, 0.001521153, 0.001517759, 
    0.001535626, 0.001527934, 0.001547978, 0.001543185, 0.001549127, 
    0.001546096, 0.001551289, 0.001546615, 0.001554711, 0.001556472, 
    0.001555269, 0.001559893, 0.001546356, 0.001551557, 0.001512382, 
    0.001512613, 0.001513688, 0.001508961, 0.001508671, 0.001504338, 
    0.001508194, 0.001509836, 0.001514003, 0.001516467, 0.001518809, 
    0.001523956, 0.001529701, 0.001537731, 0.001543496, 0.001547359, 
    0.001544991, 0.001547082, 0.001544744, 0.001543648, 0.001555812, 
    0.001548984, 0.001559228, 0.001558662, 0.001554026, 0.001558725, 
    0.001512775, 0.001511447, 0.001506834, 0.001510444, 0.001503866, 
    0.001507548, 0.001509665, 0.00151783, 0.001519624, 0.001521286, 
    0.001524569, 0.00152878, 0.001536164, 0.001542585, 0.001548443, 
    0.001548014, 0.001548165, 0.001549473, 0.001546232, 0.001550005, 
    0.001550638, 0.001548983, 0.001558586, 0.001555843, 0.00155865, 
    0.001556864, 0.001511879, 0.001514113, 0.001512906, 0.001515176, 
    0.001513577, 0.001520687, 0.001522819, 0.001532786, 0.001528697, 
    0.001535204, 0.001529358, 0.001530394, 0.001535416, 0.001529675, 
    0.00154223, 0.001533719, 0.001549524, 0.001541029, 0.001550056, 
    0.001548418, 0.00155113, 0.001553559, 0.001556614, 0.001562248, 
    0.001560944, 0.001565654, 0.001517444, 0.001520341, 0.001520087, 
    0.001523118, 0.001525359, 0.001530215, 0.001538, 0.001535073, 
    0.001540446, 0.001541524, 0.001533362, 0.001538373, 0.00152228, 
    0.001524881, 0.001523333, 0.001517673, 0.001535747, 0.001526475, 
    0.001543591, 0.001538573, 0.001553213, 0.001545934, 0.001560225, 
    0.001566328, 0.00157207, 0.001578773, 0.001521922, 0.001519954, 
    0.001523478, 0.001528351, 0.001532872, 0.001538879, 0.001539493, 
    0.001540618, 0.001543531, 0.00154598, 0.001540973, 0.001546594, 
    0.001525483, 0.001536552, 0.00151921, 0.001524434, 0.001528064, 
    0.001526472, 0.001534739, 0.001536686, 0.001544595, 0.001540508, 
    0.001564821, 0.001554071, 0.001583876, 0.001575556, 0.001519267, 
    0.001521916, 0.001531131, 0.001526747, 0.00153928, 0.001542362, 
    0.001544868, 0.001548069, 0.001548415, 0.001550311, 0.001547204, 
    0.001550189, 0.001538892, 0.001543942, 0.001530078, 0.001533454, 
    0.001531901, 0.001530198, 0.001535455, 0.001541052, 0.001541172, 
    0.001542966, 0.001548019, 0.001539331, 0.001566207, 0.001549616, 
    0.001524804, 0.001529903, 0.001530632, 0.001528657, 0.001542053, 
    0.001537201, 0.001550265, 0.001546736, 0.001552518, 0.001549645, 
    0.001549223, 0.001545532, 0.001543233, 0.001537423, 0.001532695, 
    0.001528944, 0.001529816, 0.001533936, 0.001541394, 0.001548446, 
    0.001546902, 0.001552079, 0.001538372, 0.001544121, 0.001541899, 
    0.001547692, 0.001534995, 0.001545806, 0.00153223, 0.001533421, 
    0.001537105, 0.00154451, 0.001546149, 0.001547897, 0.001546819, 
    0.001541584, 0.001540726, 0.001537015, 0.00153599, 0.001533162, 
    0.001530819, 0.00153296, 0.001535206, 0.001541586, 0.001547332, 
    0.001553593, 0.001555125, 0.001562433, 0.001556484, 0.001566299, 
    0.001557953, 0.001572397, 0.001546433, 0.001557709, 0.001537273, 
    0.001539476, 0.00154346, 0.001552594, 0.001547665, 0.00155343, 
    0.001540693, 0.001534078, 0.001532366, 0.001529171, 0.001532439, 
    0.001532174, 0.0015353, 0.001534296, 0.001541798, 0.001537769, 
    0.001549212, 0.001553384, 0.00156516, 0.001572371, 0.001579708, 
    0.001582945, 0.00158393, 0.001584342,
  0.001428863, 0.00143567, 0.001434347, 0.001439837, 0.001436791, 
    0.001440386, 0.001430243, 0.00143594, 0.001432303, 0.001429476, 
    0.001450489, 0.001440082, 0.001461297, 0.001454662, 0.00147133, 
    0.001460265, 0.00147356, 0.001471011, 0.001478685, 0.001476487, 
    0.001486301, 0.0014797, 0.001491388, 0.001484725, 0.001485767, 
    0.001479482, 0.001442176, 0.001449193, 0.00144176, 0.001442761, 
    0.001442312, 0.001436854, 0.001434104, 0.001428343, 0.001429389, 
    0.00143362, 0.001443211, 0.001439956, 0.00144816, 0.001447975, 
    0.001457107, 0.00145299, 0.001468337, 0.001463976, 0.001476578, 
    0.001473409, 0.00147643, 0.001475514, 0.001476441, 0.001471794, 
    0.001473785, 0.001469695, 0.001453761, 0.001458444, 0.001444475, 
    0.001436074, 0.001430493, 0.001426533, 0.001427092, 0.00142816, 
    0.001433645, 0.001438801, 0.001442731, 0.001445359, 0.001447948, 
    0.001455785, 0.001459933, 0.001469219, 0.001467544, 0.001470382, 
    0.001473094, 0.001477646, 0.001476897, 0.001478903, 0.001470307, 
    0.00147602, 0.001466589, 0.001469169, 0.001448652, 0.001440834, 
    0.00143751, 0.001434601, 0.001427523, 0.001432411, 0.001430484, 
    0.001435068, 0.001437981, 0.001436541, 0.001445431, 0.001441975, 
    0.001460179, 0.001452339, 0.001472778, 0.001467888, 0.00147395, 
    0.001470856, 0.001476156, 0.001471387, 0.001479649, 0.001481448, 
    0.001480219, 0.001484941, 0.001471122, 0.001476429, 0.0014365, 
    0.001436735, 0.00143783, 0.001433018, 0.001432724, 0.001428314, 
    0.001432238, 0.001433909, 0.00143815, 0.001440658, 0.001443043, 
    0.001448285, 0.00145414, 0.001462325, 0.001468205, 0.001472145, 
    0.001469729, 0.001471862, 0.001469477, 0.00146836, 0.001480774, 
    0.001473804, 0.001484262, 0.001483683, 0.00147895, 0.001483748, 
    0.0014369, 0.001435548, 0.001430854, 0.001434528, 0.001427834, 
    0.001431581, 0.001433735, 0.001442047, 0.001443873, 0.001445566, 
    0.00144891, 0.001453201, 0.001460727, 0.001467275, 0.001473252, 
    0.001472814, 0.001472968, 0.001474303, 0.001470996, 0.001474846, 
    0.001475492, 0.001473803, 0.001483606, 0.001480805, 0.001483671, 
    0.001481847, 0.001435988, 0.001438263, 0.001437033, 0.001439345, 
    0.001437716, 0.001444957, 0.001447128, 0.001457284, 0.001453116, 
    0.001459749, 0.00145379, 0.001454846, 0.001459965, 0.001454112, 
    0.001466914, 0.001458235, 0.001474355, 0.001465689, 0.001474898, 
    0.001473226, 0.001475994, 0.001478473, 0.001481592, 0.001487346, 
    0.001486014, 0.001490825, 0.001441654, 0.001444604, 0.001444344, 
    0.001447432, 0.001449715, 0.001454663, 0.001462599, 0.001459615, 
    0.001465093, 0.001466193, 0.00145787, 0.00146298, 0.001446579, 
    0.001449229, 0.001447651, 0.001441887, 0.001460303, 0.001450852, 
    0.001468302, 0.001463183, 0.00147812, 0.001470692, 0.00148528, 
    0.001491515, 0.001497383, 0.001504238, 0.001446214, 0.00144421, 
    0.001447799, 0.001452764, 0.001457371, 0.001463495, 0.001464122, 
    0.001465269, 0.00146824, 0.001470739, 0.001465632, 0.001471365, 
    0.001449843, 0.001461123, 0.001443452, 0.001448773, 0.001452472, 
    0.001450849, 0.001459274, 0.001461259, 0.001469326, 0.001465156, 
    0.001489976, 0.001478997, 0.001509457, 0.001500947, 0.001443509, 
    0.001446207, 0.001455597, 0.00145113, 0.001463904, 0.001467048, 
    0.001469604, 0.00147287, 0.001473223, 0.001475158, 0.001471987, 
    0.001475033, 0.001463508, 0.001468659, 0.001454524, 0.001457964, 
    0.001456382, 0.001454645, 0.001460004, 0.001465712, 0.001465834, 
    0.001467664, 0.001472821, 0.001463956, 0.001491393, 0.00147445, 
    0.001449149, 0.001454346, 0.001455088, 0.001453075, 0.001466733, 
    0.001461785, 0.001475111, 0.00147151, 0.001477411, 0.001474479, 
    0.001474047, 0.001470281, 0.001467936, 0.001462011, 0.00145719, 
    0.001453367, 0.001454256, 0.001458456, 0.001466061, 0.001473255, 
    0.001471679, 0.001476962, 0.001462978, 0.001468842, 0.001466576, 
    0.001472485, 0.001459536, 0.001470563, 0.001456717, 0.001457931, 
    0.001461686, 0.00146924, 0.001470911, 0.001472695, 0.001471594, 
    0.001466254, 0.001465379, 0.001461595, 0.00146055, 0.001457666, 
    0.001455279, 0.00145746, 0.001459751, 0.001466257, 0.001472119, 
    0.001478509, 0.001480072, 0.001487537, 0.001481461, 0.001491487, 
    0.001482963, 0.001497719, 0.001471202, 0.001482712, 0.001461857, 
    0.001464105, 0.001468169, 0.001477489, 0.001472458, 0.001478342, 
    0.001465345, 0.001458601, 0.001456856, 0.0014536, 0.00145693, 
    0.001456659, 0.001459846, 0.001458822, 0.001466473, 0.001462363, 
    0.001474036, 0.001478295, 0.001490321, 0.001497692, 0.001505193, 
    0.001508505, 0.001509513, 0.001509934,
  0.001341426, 0.001347692, 0.001346474, 0.00135153, 0.001348725, 
    0.001352036, 0.001342696, 0.001347941, 0.001344592, 0.00134199, 
    0.001361351, 0.001351756, 0.001371329, 0.001365201, 0.001380602, 
    0.001370375, 0.001382666, 0.001380307, 0.001387408, 0.001385373, 
    0.001394464, 0.001388348, 0.001399179, 0.001393003, 0.001393969, 
    0.001388146, 0.001353686, 0.001360156, 0.001353302, 0.001354225, 
    0.001353811, 0.001348783, 0.00134625, 0.001340947, 0.00134191, 
    0.001345804, 0.00135464, 0.001351639, 0.001359202, 0.001359031, 
    0.001367459, 0.001363658, 0.001377834, 0.001373803, 0.001385458, 
    0.001382526, 0.00138532, 0.001384473, 0.001385332, 0.001381031, 
    0.001382873, 0.00137909, 0.00136437, 0.001368693, 0.001355805, 
    0.001348064, 0.001342926, 0.001339282, 0.001339797, 0.001340779, 
    0.001345827, 0.001350576, 0.001354196, 0.001356619, 0.001359007, 
    0.001366239, 0.001370069, 0.00137865, 0.001377101, 0.001379726, 
    0.001382234, 0.001386447, 0.001385753, 0.00138761, 0.001379656, 
    0.001384942, 0.001376218, 0.001378603, 0.001359657, 0.001352449, 
    0.001349387, 0.001346708, 0.001340193, 0.001344692, 0.001342918, 
    0.001347138, 0.00134982, 0.001348493, 0.001356685, 0.0013535, 
    0.001370296, 0.001363057, 0.001381941, 0.001377419, 0.001383026, 
    0.001380164, 0.001385068, 0.001380654, 0.001388301, 0.001389967, 
    0.001388829, 0.001393203, 0.00138041, 0.00138532, 0.001348456, 
    0.001348673, 0.001349681, 0.00134525, 0.001344979, 0.001340921, 
    0.001344532, 0.00134607, 0.001349976, 0.001352287, 0.001354484, 
    0.001359318, 0.001364719, 0.001372278, 0.001377712, 0.001381356, 
    0.001379121, 0.001381094, 0.001378889, 0.001377855, 0.001389343, 
    0.001382891, 0.001392573, 0.001392037, 0.001387654, 0.001392098, 
    0.001348825, 0.00134758, 0.001343258, 0.00134664, 0.001340479, 
    0.001343927, 0.00134591, 0.001353566, 0.001355249, 0.00135681, 
    0.001359893, 0.001363852, 0.001370802, 0.001376852, 0.00138238, 
    0.001381975, 0.001382117, 0.001383353, 0.001380293, 0.001383855, 
    0.001384453, 0.00138289, 0.001391966, 0.001389372, 0.001392026, 
    0.001390337, 0.001347984, 0.001350079, 0.001348947, 0.001351077, 
    0.001349577, 0.001356249, 0.001358251, 0.001367622, 0.001363775, 
    0.001369898, 0.001364396, 0.001365371, 0.001370099, 0.001364694, 
    0.001376519, 0.0013685, 0.001383401, 0.001375387, 0.001383903, 
    0.001382356, 0.001384917, 0.001387213, 0.001390101, 0.001395432, 
    0.001394197, 0.001398658, 0.001353204, 0.001355923, 0.001355684, 
    0.00135853, 0.001360636, 0.001365202, 0.001372531, 0.001369774, 
    0.001374835, 0.001375852, 0.001368163, 0.001372883, 0.001357744, 
    0.001360188, 0.001358733, 0.001353419, 0.00137041, 0.001361686, 
    0.001377802, 0.00137307, 0.001386885, 0.001380012, 0.001393518, 
    0.001399298, 0.001404741, 0.001411108, 0.001357408, 0.00135556, 
    0.001358869, 0.00136345, 0.001367702, 0.001373359, 0.001373938, 
    0.001374998, 0.001377745, 0.001380055, 0.001375334, 0.001380634, 
    0.001360756, 0.001371167, 0.001354861, 0.001359768, 0.00136318, 
    0.001361683, 0.001369459, 0.001371293, 0.001378749, 0.001374894, 
    0.001397871, 0.001387698, 0.001415958, 0.001408051, 0.001354914, 
    0.001357401, 0.001366064, 0.001361941, 0.001373737, 0.001376642, 
    0.001379005, 0.001382027, 0.001382353, 0.001384144, 0.00138121, 
    0.001384028, 0.001373371, 0.001378132, 0.001365073, 0.00136825, 
    0.001366788, 0.001365186, 0.001370133, 0.001375408, 0.00137552, 
    0.001377212, 0.001381983, 0.001373784, 0.001399186, 0.00138349, 
    0.001360115, 0.00136491, 0.001365594, 0.001363736, 0.001376351, 
    0.001371778, 0.001384101, 0.001380768, 0.001386228, 0.001383515, 
    0.001383116, 0.001379632, 0.001377464, 0.001371988, 0.001367535, 
    0.001364006, 0.001364826, 0.001368704, 0.001375731, 0.001382383, 
    0.001380925, 0.001385813, 0.001372881, 0.001378302, 0.001376206, 
    0.001381671, 0.001369701, 0.001379894, 0.001367098, 0.001368219, 
    0.001371688, 0.00137867, 0.001380214, 0.001381865, 0.001380846, 
    0.001375909, 0.0013751, 0.001371603, 0.001370638, 0.001367975, 
    0.00136577, 0.001367784, 0.0013699, 0.001375911, 0.001381332, 
    0.001387245, 0.001388693, 0.00139561, 0.001389979, 0.001399273, 
    0.001391372, 0.001405054, 0.001380485, 0.001391139, 0.001371845, 
    0.001373922, 0.001377679, 0.001386302, 0.001381645, 0.001387091, 
    0.001375068, 0.001368838, 0.001367226, 0.00136422, 0.001367295, 
    0.001367045, 0.001369987, 0.001369042, 0.00137611, 0.001372313, 
    0.001383106, 0.001387048, 0.00139819, 0.001405029, 0.001411995, 
    0.001415072, 0.001416009, 0.001416401,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.216114e-06, 1.22666e-06, 1.224606e-06, 1.233139e-06, 1.228402e-06, 
    1.233994e-06, 1.218248e-06, 1.227078e-06, 1.221437e-06, 1.21706e-06, 
    1.249786e-06, 1.233519e-06, 1.266805e-06, 1.256342e-06, 1.282712e-06, 
    1.265173e-06, 1.286264e-06, 1.282204e-06, 1.294443e-06, 1.290931e-06, 
    1.306651e-06, 1.296066e-06, 1.31484e-06, 1.304119e-06, 1.305793e-06, 
    1.295717e-06, 1.236785e-06, 1.247756e-06, 1.236137e-06, 1.237697e-06, 
    1.236997e-06, 1.228498e-06, 1.224227e-06, 1.215309e-06, 1.216925e-06, 
    1.223477e-06, 1.238399e-06, 1.233323e-06, 1.246137e-06, 1.245847e-06, 
    1.260192e-06, 1.253713e-06, 1.277955e-06, 1.27104e-06, 1.291077e-06, 
    1.286022e-06, 1.290839e-06, 1.289377e-06, 1.290858e-06, 1.283449e-06, 
    1.28662e-06, 1.280111e-06, 1.254927e-06, 1.262301e-06, 1.240373e-06, 
    1.227285e-06, 1.218634e-06, 1.212514e-06, 1.213378e-06, 1.215026e-06, 
    1.223515e-06, 1.231525e-06, 1.237648e-06, 1.241753e-06, 1.245804e-06, 
    1.258109e-06, 1.264649e-06, 1.279356e-06, 1.276695e-06, 1.281204e-06, 
    1.28552e-06, 1.292782e-06, 1.291585e-06, 1.29479e-06, 1.281084e-06, 
    1.290184e-06, 1.27518e-06, 1.279274e-06, 1.246907e-06, 1.234692e-06, 
    1.229518e-06, 1.224999e-06, 1.214042e-06, 1.221603e-06, 1.218619e-06, 
    1.225724e-06, 1.230249e-06, 1.22801e-06, 1.241865e-06, 1.236469e-06, 
    1.265037e-06, 1.252689e-06, 1.285016e-06, 1.277241e-06, 1.286883e-06, 
    1.281958e-06, 1.290402e-06, 1.282801e-06, 1.295984e-06, 1.298864e-06, 
    1.296895e-06, 1.304465e-06, 1.282379e-06, 1.290837e-06, 1.227948e-06, 
    1.228313e-06, 1.230014e-06, 1.222543e-06, 1.222087e-06, 1.215264e-06, 
    1.221334e-06, 1.223924e-06, 1.230512e-06, 1.234417e-06, 1.238135e-06, 
    1.246332e-06, 1.255519e-06, 1.268427e-06, 1.277744e-06, 1.284009e-06, 
    1.280165e-06, 1.283558e-06, 1.279765e-06, 1.277989e-06, 1.297784e-06, 
    1.286649e-06, 1.303375e-06, 1.302446e-06, 1.294865e-06, 1.30255e-06, 
    1.228569e-06, 1.226469e-06, 1.219191e-06, 1.224884e-06, 1.214522e-06, 
    1.220316e-06, 1.223654e-06, 1.236581e-06, 1.239431e-06, 1.242076e-06, 
    1.24731e-06, 1.254043e-06, 1.265902e-06, 1.276268e-06, 1.285771e-06, 
    1.285073e-06, 1.285318e-06, 1.287445e-06, 1.282179e-06, 1.288311e-06, 
    1.289341e-06, 1.286647e-06, 1.302321e-06, 1.297833e-06, 1.302426e-06, 
    1.299502e-06, 1.227151e-06, 1.230687e-06, 1.228775e-06, 1.232371e-06, 
    1.229837e-06, 1.241124e-06, 1.244519e-06, 1.260469e-06, 1.25391e-06, 
    1.264358e-06, 1.254969e-06, 1.25663e-06, 1.264698e-06, 1.255475e-06, 
    1.275694e-06, 1.261967e-06, 1.287528e-06, 1.273752e-06, 1.288393e-06, 
    1.285728e-06, 1.290142e-06, 1.294102e-06, 1.299093e-06, 1.308329e-06, 
    1.306187e-06, 1.313931e-06, 1.235968e-06, 1.240573e-06, 1.240167e-06, 
    1.244995e-06, 1.248572e-06, 1.256343e-06, 1.268861e-06, 1.264146e-06, 
    1.272809e-06, 1.274551e-06, 1.261393e-06, 1.269463e-06, 1.243659e-06, 
    1.247808e-06, 1.245337e-06, 1.236329e-06, 1.26523e-06, 1.250353e-06, 
    1.277896e-06, 1.269783e-06, 1.293537e-06, 1.281694e-06, 1.305009e-06, 
    1.315043e-06, 1.324525e-06, 1.335649e-06, 1.24309e-06, 1.239957e-06, 
    1.24557e-06, 1.253357e-06, 1.260607e-06, 1.270279e-06, 1.27127e-06, 
    1.273087e-06, 1.2778e-06, 1.28177e-06, 1.273661e-06, 1.282765e-06, 
    1.248771e-06, 1.266525e-06, 1.238771e-06, 1.247094e-06, 1.252896e-06, 
    1.250349e-06, 1.263606e-06, 1.266741e-06, 1.279522e-06, 1.272907e-06, 
    1.312562e-06, 1.294938e-06, 1.344154e-06, 1.330302e-06, 1.238863e-06, 
    1.243079e-06, 1.257811e-06, 1.25079e-06, 1.270926e-06, 1.275908e-06, 
    1.279966e-06, 1.285162e-06, 1.285724e-06, 1.288809e-06, 1.283755e-06, 
    1.288609e-06, 1.270298e-06, 1.278464e-06, 1.256122e-06, 1.26154e-06, 
    1.259046e-06, 1.256312e-06, 1.264757e-06, 1.273787e-06, 1.273981e-06, 
    1.276883e-06, 1.28508e-06, 1.271005e-06, 1.314844e-06, 1.287676e-06, 
    1.247685e-06, 1.255842e-06, 1.25701e-06, 1.253845e-06, 1.275407e-06, 
    1.267572e-06, 1.288734e-06, 1.282996e-06, 1.292404e-06, 1.287725e-06, 
    1.287036e-06, 1.281041e-06, 1.277316e-06, 1.26793e-06, 1.260319e-06, 
    1.254303e-06, 1.2557e-06, 1.262314e-06, 1.27434e-06, 1.285773e-06, 
    1.283264e-06, 1.291686e-06, 1.269457e-06, 1.278753e-06, 1.275155e-06, 
    1.284546e-06, 1.26402e-06, 1.281489e-06, 1.259575e-06, 1.261488e-06, 
    1.267416e-06, 1.279386e-06, 1.282043e-06, 1.284883e-06, 1.28313e-06, 
    1.274647e-06, 1.273261e-06, 1.267271e-06, 1.26562e-06, 1.26107e-06, 
    1.257309e-06, 1.260745e-06, 1.264358e-06, 1.27465e-06, 1.283963e-06, 
    1.294157e-06, 1.296658e-06, 1.308634e-06, 1.29888e-06, 1.314996e-06, 
    1.301286e-06, 1.325066e-06, 1.282506e-06, 1.300888e-06, 1.267687e-06, 
    1.271242e-06, 1.277685e-06, 1.292529e-06, 1.284504e-06, 1.293891e-06, 
    1.273206e-06, 1.262543e-06, 1.259792e-06, 1.254668e-06, 1.259909e-06, 
    1.259482e-06, 1.264508e-06, 1.262891e-06, 1.274992e-06, 1.268485e-06, 
    1.287017e-06, 1.293816e-06, 1.313117e-06, 1.325023e-06, 1.337203e-06, 
    1.342598e-06, 1.344242e-06, 1.34493e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  7.708913e-06, 7.743616e-06, 7.736852e-06, 7.764858e-06, 7.749315e-06, 
    7.76764e-06, 7.71591e-06, 7.744933e-06, 7.726395e-06, 7.711974e-06, 
    7.81919e-06, 7.766045e-06, 7.874544e-06, 7.840557e-06, 7.925979e-06, 
    7.869225e-06, 7.937429e-06, 7.924335e-06, 7.963758e-06, 7.952446e-06, 
    8.002879e-06, 7.968952e-06, 8.029067e-06, 7.994768e-06, 8.000115e-06, 
    7.96779e-06, 7.776805e-06, 7.812624e-06, 7.774664e-06, 7.779771e-06, 
    7.777473e-06, 7.749596e-06, 7.735551e-06, 7.706197e-06, 7.711514e-06, 
    7.733072e-06, 7.782009e-06, 7.765381e-06, 7.807289e-06, 7.806344e-06, 
    7.853047e-06, 7.831974e-06, 7.910604e-06, 7.888225e-06, 7.952908e-06, 
    7.936614e-06, 7.952124e-06, 7.947408e-06, 7.952161e-06, 7.928288e-06, 
    7.938496e-06, 7.917502e-06, 7.836014e-06, 7.859977e-06, 7.788513e-06, 
    7.745589e-06, 7.717145e-06, 7.696976e-06, 7.699809e-06, 7.705244e-06, 
    7.733182e-06, 7.759483e-06, 7.779544e-06, 7.792958e-06, 7.806184e-06, 
    7.846247e-06, 7.867493e-06, 7.915102e-06, 7.906513e-06, 7.921057e-06, 
    7.934985e-06, 7.958357e-06, 7.954505e-06, 7.964796e-06, 7.920639e-06, 
    7.94997e-06, 7.901547e-06, 7.914779e-06, 7.809815e-06, 7.769902e-06, 
    7.752911e-06, 7.738076e-06, 7.701995e-06, 7.726899e-06, 7.717068e-06, 
    7.740434e-06, 7.755288e-06, 7.747928e-06, 7.793315e-06, 7.775647e-06, 
    7.868741e-06, 7.828606e-06, 7.93337e-06, 7.908257e-06, 7.939368e-06, 
    7.923488e-06, 7.950682e-06, 7.926193e-06, 7.968619e-06, 7.977865e-06, 
    7.971528e-06, 7.995824e-06, 7.924783e-06, 7.952036e-06, 7.747768e-06, 
    7.748968e-06, 7.754544e-06, 7.729979e-06, 7.728478e-06, 7.705999e-06, 
    7.725982e-06, 7.734498e-06, 7.756132e-06, 7.768919e-06, 7.781086e-06, 
    7.807877e-06, 7.837803e-06, 7.879716e-06, 7.909874e-06, 7.930092e-06, 
    7.917685e-06, 7.928622e-06, 7.916376e-06, 7.910629e-06, 7.974373e-06, 
    7.938556e-06, 7.992304e-06, 7.989331e-06, 7.964974e-06, 7.989642e-06, 
    7.749793e-06, 7.742887e-06, 7.718943e-06, 7.737664e-06, 7.703537e-06, 
    7.722624e-06, 7.73359e-06, 7.775992e-06, 7.785321e-06, 7.793969e-06, 
    7.811055e-06, 7.832989e-06, 7.871521e-06, 7.905081e-06, 7.935764e-06, 
    7.933503e-06, 7.934291e-06, 7.941131e-06, 7.924147e-06, 7.943903e-06, 
    7.947207e-06, 7.938536e-06, 7.988908e-06, 7.974507e-06, 7.989234e-06, 
    7.979844e-06, 7.74512e-06, 7.756711e-06, 7.750428e-06, 7.762223e-06, 
    7.753893e-06, 7.790858e-06, 7.801938e-06, 7.853889e-06, 7.832555e-06, 
    7.866513e-06, 7.83599e-06, 7.841392e-06, 7.867572e-06, 7.83762e-06, 
    7.903194e-06, 7.858687e-06, 7.941388e-06, 7.896871e-06, 7.944162e-06, 
    7.935563e-06, 7.949772e-06, 7.96251e-06, 7.978529e-06, 8.008126e-06, 
    8.001255e-06, 8.02603e-06, 7.774015e-06, 7.789064e-06, 7.787743e-06, 
    7.803507e-06, 7.815167e-06, 7.84049e-06, 7.881123e-06, 7.865823e-06, 
    7.893892e-06, 7.899531e-06, 7.856861e-06, 7.883034e-06, 7.799071e-06, 
    7.812597e-06, 7.804539e-06, 7.775071e-06, 7.869263e-06, 7.820868e-06, 
    7.910272e-06, 7.884008e-06, 7.960668e-06, 7.922508e-06, 7.997474e-06, 
    8.029555e-06, 8.059807e-06, 8.095139e-06, 7.797288e-06, 7.787037e-06, 
    7.80537e-06, 7.830751e-06, 7.854327e-06, 7.885707e-06, 7.888913e-06, 
    7.894781e-06, 7.910015e-06, 7.922837e-06, 7.89661e-06, 7.926029e-06, 
    7.815709e-06, 7.873468e-06, 7.78305e-06, 7.810236e-06, 7.829143e-06, 
    7.820851e-06, 7.863972e-06, 7.87413e-06, 7.915478e-06, 7.894098e-06, 
    8.021601e-06, 7.965125e-06, 8.122089e-06, 8.078146e-06, 7.783448e-06, 
    7.797224e-06, 7.845229e-06, 7.822377e-06, 7.887784e-06, 7.903906e-06, 
    7.917007e-06, 7.93377e-06, 7.935569e-06, 7.945508e-06, 7.929207e-06, 
    7.944851e-06, 7.885685e-06, 7.912107e-06, 7.839658e-06, 7.857256e-06, 
    7.849153e-06, 7.840251e-06, 7.867681e-06, 7.896927e-06, 7.897557e-06, 
    7.906925e-06, 7.93334e-06, 7.887897e-06, 8.028837e-06, 7.941685e-06, 
    7.812254e-06, 7.838805e-06, 7.842609e-06, 7.832314e-06, 7.902265e-06, 
    7.876895e-06, 7.945267e-06, 7.926762e-06, 7.957059e-06, 7.941996e-06, 
    7.939761e-06, 7.920428e-06, 7.908374e-06, 7.877989e-06, 7.853273e-06, 
    7.833712e-06, 7.838243e-06, 7.859739e-06, 7.898697e-06, 7.935624e-06, 
    7.927519e-06, 7.954652e-06, 7.882866e-06, 7.912938e-06, 7.901289e-06, 
    7.931628e-06, 7.86538e-06, 7.921886e-06, 7.850938e-06, 7.857142e-06, 
    7.876368e-06, 7.915092e-06, 7.923671e-06, 7.932826e-06, 7.927162e-06, 
    7.899751e-06, 7.895258e-06, 7.875849e-06, 7.870478e-06, 7.855715e-06, 
    7.843471e-06, 7.854639e-06, 7.866349e-06, 7.899704e-06, 7.929771e-06, 
    7.962586e-06, 7.970628e-06, 8.00898e-06, 7.97772e-06, 8.029278e-06, 
    7.985392e-06, 8.061394e-06, 7.925162e-06, 7.984304e-06, 7.87725e-06, 
    7.888757e-06, 7.909582e-06, 7.957424e-06, 7.931586e-06, 7.961802e-06, 
    7.895078e-06, 7.860486e-06, 7.851554e-06, 7.834886e-06, 7.85192e-06, 
    7.850535e-06, 7.866847e-06, 7.861589e-06, 7.900788e-06, 7.879723e-06, 
    7.939591e-06, 7.961469e-06, 8.023331e-06, 8.061292e-06, 8.100009e-06, 
    8.117095e-06, 8.122299e-06, 8.124465e-06,
  4.017422e-06, 4.048206e-06, 4.042216e-06, 4.067095e-06, 4.05329e-06, 
    4.069589e-06, 4.023659e-06, 4.049428e-06, 4.032971e-06, 4.020194e-06, 
    4.115537e-06, 4.068208e-06, 4.164955e-06, 4.1346e-06, 4.211023e-06, 
    4.160221e-06, 4.221297e-06, 4.209562e-06, 4.244937e-06, 4.234792e-06, 
    4.280145e-06, 4.249623e-06, 4.303738e-06, 4.272852e-06, 4.277676e-06, 
    4.248616e-06, 4.077722e-06, 4.10963e-06, 4.075833e-06, 4.080377e-06, 
    4.078339e-06, 4.053572e-06, 4.041109e-06, 4.015078e-06, 4.0198e-06, 
    4.038924e-06, 4.08242e-06, 4.06764e-06, 4.104945e-06, 4.104101e-06, 
    4.14578e-06, 4.126967e-06, 4.197268e-06, 4.177242e-06, 4.235215e-06, 
    4.220606e-06, 4.234527e-06, 4.230305e-06, 4.234582e-06, 4.213165e-06, 
    4.222336e-06, 4.20351e-06, 4.130487e-06, 4.151894e-06, 4.088169e-06, 
    4.050026e-06, 4.024786e-06, 4.006908e-06, 4.009434e-06, 4.014249e-06, 
    4.039036e-06, 4.062402e-06, 4.080242e-06, 4.092191e-06, 4.10398e-06, 
    4.139723e-06, 4.158705e-06, 4.201318e-06, 4.193621e-06, 4.206667e-06, 
    4.219154e-06, 4.240141e-06, 4.236685e-06, 4.245939e-06, 4.206328e-06, 
    4.232636e-06, 4.189239e-06, 4.20109e-06, 4.107162e-06, 4.071626e-06, 
    4.056538e-06, 4.043367e-06, 4.011375e-06, 4.033456e-06, 4.024745e-06, 
    4.045485e-06, 4.058682e-06, 4.052155e-06, 4.092518e-06, 4.076806e-06, 
    4.159831e-06, 4.12399e-06, 4.217697e-06, 4.195201e-06, 4.223096e-06, 
    4.208855e-06, 4.233266e-06, 4.211294e-06, 4.249388e-06, 4.257697e-06, 
    4.252017e-06, 4.273858e-06, 4.210076e-06, 4.234525e-06, 4.05197e-06, 
    4.053034e-06, 4.057997e-06, 4.036201e-06, 4.03487e-06, 4.014947e-06, 
    4.032675e-06, 4.040232e-06, 4.05945e-06, 4.07083e-06, 4.08166e-06, 
    4.105513e-06, 4.132212e-06, 4.169666e-06, 4.196658e-06, 4.214787e-06, 
    4.203669e-06, 4.213484e-06, 4.202511e-06, 4.197373e-06, 4.254581e-06, 
    4.22242e-06, 4.270714e-06, 4.268037e-06, 4.246158e-06, 4.268339e-06, 
    4.053783e-06, 4.047658e-06, 4.026417e-06, 4.043036e-06, 4.01278e-06, 
    4.029702e-06, 4.039443e-06, 4.077129e-06, 4.085433e-06, 4.093132e-06, 
    4.108359e-06, 4.127929e-06, 4.162346e-06, 4.192384e-06, 4.219882e-06, 
    4.217865e-06, 4.218575e-06, 4.224724e-06, 4.209496e-06, 4.227226e-06, 
    4.230202e-06, 4.222419e-06, 4.267678e-06, 4.25473e-06, 4.26798e-06, 
    4.259548e-06, 4.049649e-06, 4.059959e-06, 4.054386e-06, 4.064867e-06, 
    4.05748e-06, 4.090357e-06, 4.100234e-06, 4.146581e-06, 4.127543e-06, 
    4.157866e-06, 4.130621e-06, 4.135442e-06, 4.158846e-06, 4.132093e-06, 
    4.190721e-06, 4.150929e-06, 4.224963e-06, 4.185092e-06, 4.227466e-06, 
    4.219763e-06, 4.232521e-06, 4.243958e-06, 4.258367e-06, 4.284995e-06, 
    4.278824e-06, 4.301132e-06, 4.07535e-06, 4.088754e-06, 4.087578e-06, 
    4.101626e-06, 4.112027e-06, 4.134611e-06, 4.170925e-06, 4.157257e-06, 
    4.182369e-06, 4.187415e-06, 4.149272e-06, 4.172671e-06, 4.097739e-06, 
    4.109805e-06, 4.102623e-06, 4.076404e-06, 4.160398e-06, 4.117207e-06, 
    4.197103e-06, 4.173605e-06, 4.242326e-06, 4.208092e-06, 4.275428e-06, 
    4.304323e-06, 4.331608e-06, 4.363548e-06, 4.096083e-06, 4.086965e-06, 
    4.1033e-06, 4.125932e-06, 4.146988e-06, 4.175036e-06, 4.177913e-06, 
    4.183175e-06, 4.196825e-06, 4.208312e-06, 4.184835e-06, 4.211194e-06, 
    4.112596e-06, 4.164158e-06, 4.083517e-06, 4.107729e-06, 4.124598e-06, 
    4.1172e-06, 4.155697e-06, 4.164789e-06, 4.20181e-06, 4.182659e-06, 
    4.297181e-06, 4.246368e-06, 4.387941e-06, 4.348201e-06, 4.083781e-06, 
    4.096054e-06, 4.138871e-06, 4.118478e-06, 4.176914e-06, 4.191344e-06, 
    4.203093e-06, 4.218122e-06, 4.219749e-06, 4.228666e-06, 4.214058e-06, 
    4.22809e-06, 4.175096e-06, 4.198747e-06, 4.133974e-06, 4.149701e-06, 
    4.142464e-06, 4.134529e-06, 4.159038e-06, 4.185203e-06, 4.185771e-06, 
    4.194173e-06, 4.217871e-06, 4.177151e-06, 4.303741e-06, 4.225381e-06, 
    4.109452e-06, 4.133151e-06, 4.136549e-06, 4.127358e-06, 4.189896e-06, 
    4.167194e-06, 4.228449e-06, 4.211862e-06, 4.239055e-06, 4.225533e-06, 
    4.223545e-06, 4.206207e-06, 4.195425e-06, 4.168232e-06, 4.146159e-06, 
    4.128692e-06, 4.132751e-06, 4.151948e-06, 4.186808e-06, 4.219893e-06, 
    4.212636e-06, 4.236986e-06, 4.172666e-06, 4.199587e-06, 4.189172e-06, 
    4.216351e-06, 4.156892e-06, 4.207482e-06, 4.143996e-06, 4.149549e-06, 
    4.166744e-06, 4.20141e-06, 4.209106e-06, 4.217315e-06, 4.21225e-06, 
    4.187696e-06, 4.183681e-06, 4.166327e-06, 4.161537e-06, 4.14834e-06, 
    4.137424e-06, 4.147395e-06, 4.157876e-06, 4.187709e-06, 4.214659e-06, 
    4.24412e-06, 4.251344e-06, 4.285867e-06, 4.257745e-06, 4.304177e-06, 
    4.264674e-06, 4.333152e-06, 4.210432e-06, 4.263529e-06, 4.167529e-06, 
    4.177833e-06, 4.196487e-06, 4.239407e-06, 4.216223e-06, 4.243345e-06, 
    4.183525e-06, 4.152607e-06, 4.144631e-06, 4.129751e-06, 4.144972e-06, 
    4.143733e-06, 4.158316e-06, 4.153628e-06, 4.188701e-06, 4.169848e-06, 
    4.223493e-06, 4.243132e-06, 4.298789e-06, 4.333038e-06, 4.368017e-06, 
    4.383489e-06, 4.388203e-06, 4.390174e-06,
  3.798637e-06, 3.832563e-06, 3.825959e-06, 3.853395e-06, 3.838166e-06, 
    3.856147e-06, 3.805506e-06, 3.833911e-06, 3.815768e-06, 3.801688e-06, 
    3.906881e-06, 3.854622e-06, 3.961507e-06, 3.927936e-06, 4.012506e-06, 
    3.956272e-06, 4.023888e-06, 4.010884e-06, 4.050089e-06, 4.03884e-06, 
    4.089155e-06, 4.055285e-06, 4.115349e-06, 4.081058e-06, 4.086412e-06, 
    4.054169e-06, 3.865118e-06, 3.900357e-06, 3.863034e-06, 3.868049e-06, 
    3.865799e-06, 3.838479e-06, 3.824741e-06, 3.796052e-06, 3.801254e-06, 
    3.822331e-06, 3.870306e-06, 3.853993e-06, 3.895169e-06, 3.894238e-06, 
    3.940295e-06, 3.9195e-06, 3.997267e-06, 3.975098e-06, 4.03931e-06, 
    4.023119e-06, 4.038548e-06, 4.033867e-06, 4.038609e-06, 4.014875e-06, 
    4.025036e-06, 4.00418e-06, 3.92339e-06, 3.947058e-06, 3.87665e-06, 
    3.834575e-06, 3.806749e-06, 3.787055e-06, 3.789836e-06, 3.795141e-06, 
    3.822454e-06, 3.848216e-06, 3.867898e-06, 3.881088e-06, 3.894104e-06, 
    3.933606e-06, 3.954594e-06, 4.001754e-06, 3.993229e-06, 4.007679e-06, 
    4.02151e-06, 4.044772e-06, 4.04094e-06, 4.051201e-06, 4.007301e-06, 
    4.036453e-06, 3.988376e-06, 4.0015e-06, 3.897632e-06, 3.858392e-06, 
    3.841754e-06, 3.827227e-06, 3.791975e-06, 3.816303e-06, 3.806705e-06, 
    3.829561e-06, 3.844114e-06, 3.836913e-06, 3.881449e-06, 3.864107e-06, 
    3.955839e-06, 3.916212e-06, 4.019896e-06, 3.994979e-06, 4.025878e-06, 
    4.010099e-06, 4.037151e-06, 4.012801e-06, 4.055024e-06, 4.064242e-06, 
    4.057942e-06, 4.082171e-06, 4.011453e-06, 4.038547e-06, 3.836711e-06, 
    3.837885e-06, 3.843357e-06, 3.819329e-06, 3.817862e-06, 3.795909e-06, 
    3.815441e-06, 3.823771e-06, 3.844959e-06, 3.857513e-06, 3.869464e-06, 
    3.895799e-06, 3.9253e-06, 3.966717e-06, 3.996592e-06, 4.016671e-06, 
    4.004354e-06, 4.015227e-06, 4.003073e-06, 3.997382e-06, 4.060786e-06, 
    4.02513e-06, 4.078683e-06, 4.075712e-06, 4.051445e-06, 4.076046e-06, 
    3.838709e-06, 3.831956e-06, 3.808545e-06, 3.826861e-06, 3.793522e-06, 
    3.812166e-06, 3.822904e-06, 3.864466e-06, 3.873628e-06, 3.882127e-06, 
    3.898941e-06, 3.920563e-06, 3.958618e-06, 3.991861e-06, 4.022316e-06, 
    4.020081e-06, 4.020868e-06, 4.027682e-06, 4.01081e-06, 4.030455e-06, 
    4.033755e-06, 4.025128e-06, 4.075314e-06, 4.060949e-06, 4.075649e-06, 
    4.066294e-06, 3.834151e-06, 3.845521e-06, 3.839375e-06, 3.850935e-06, 
    3.842788e-06, 3.879067e-06, 3.889973e-06, 3.941186e-06, 3.920136e-06, 
    3.953664e-06, 3.923537e-06, 3.928867e-06, 3.954754e-06, 3.925164e-06, 
    3.990023e-06, 3.945995e-06, 4.027947e-06, 3.983794e-06, 4.03072e-06, 
    4.022184e-06, 4.036324e-06, 4.049004e-06, 4.064984e-06, 4.094535e-06, 
    4.087684e-06, 4.112453e-06, 3.8625e-06, 3.877296e-06, 3.875995e-06, 
    3.891505e-06, 3.902994e-06, 3.927947e-06, 3.968109e-06, 3.952986e-06, 
    3.980771e-06, 3.986359e-06, 3.944155e-06, 3.970042e-06, 3.887215e-06, 
    3.900542e-06, 3.892606e-06, 3.863665e-06, 3.956465e-06, 3.908719e-06, 
    3.997086e-06, 3.971074e-06, 4.047195e-06, 4.009258e-06, 4.083915e-06, 
    4.116003e-06, 4.146314e-06, 4.181841e-06, 3.885385e-06, 3.875319e-06, 
    3.893353e-06, 3.918359e-06, 3.941631e-06, 3.972657e-06, 3.97584e-06, 
    3.981665e-06, 3.996775e-06, 4.009498e-06, 3.983505e-06, 4.01269e-06, 
    3.903631e-06, 3.960623e-06, 3.871514e-06, 3.89825e-06, 3.916884e-06, 
    3.908708e-06, 3.95126e-06, 3.961318e-06, 4.0023e-06, 3.981093e-06, 
    4.108071e-06, 4.051681e-06, 4.208986e-06, 4.164768e-06, 3.871804e-06, 
    3.885351e-06, 3.932658e-06, 3.910119e-06, 3.974734e-06, 3.990708e-06, 
    4.003717e-06, 4.020368e-06, 4.022169e-06, 4.032051e-06, 4.015863e-06, 
    4.031412e-06, 3.972724e-06, 3.998905e-06, 3.927242e-06, 3.94463e-06, 
    3.936628e-06, 3.927856e-06, 3.954956e-06, 3.983913e-06, 3.984537e-06, 
    3.993842e-06, 4.020104e-06, 3.974997e-06, 4.115365e-06, 4.028423e-06, 
    3.900147e-06, 3.926338e-06, 3.93009e-06, 3.91993e-06, 3.989105e-06, 
    3.96398e-06, 4.031811e-06, 4.01343e-06, 4.043567e-06, 4.028579e-06, 
    4.026376e-06, 4.007167e-06, 3.995227e-06, 3.96513e-06, 3.940715e-06, 
    3.921404e-06, 3.925891e-06, 3.947117e-06, 3.985689e-06, 4.02233e-06, 
    4.014291e-06, 4.041273e-06, 3.970034e-06, 3.999837e-06, 3.988305e-06, 
    4.018405e-06, 3.952584e-06, 4.008591e-06, 3.938321e-06, 3.944462e-06, 
    3.963482e-06, 4.001859e-06, 4.010377e-06, 4.019474e-06, 4.013861e-06, 
    3.986671e-06, 3.982226e-06, 3.96302e-06, 3.957722e-06, 3.943125e-06, 
    3.931055e-06, 3.942081e-06, 3.953674e-06, 3.986684e-06, 4.016532e-06, 
    4.049184e-06, 4.057194e-06, 4.09551e-06, 4.064302e-06, 4.115851e-06, 
    4.071998e-06, 4.148042e-06, 4.011854e-06, 4.07072e-06, 3.96435e-06, 
    3.975751e-06, 3.996407e-06, 4.043962e-06, 4.018263e-06, 4.048327e-06, 
    3.982052e-06, 3.947848e-06, 3.939024e-06, 3.922576e-06, 3.9394e-06, 
    3.938031e-06, 3.954157e-06, 3.948972e-06, 3.987782e-06, 3.966915e-06, 
    4.026319e-06, 4.048091e-06, 4.109852e-06, 4.147909e-06, 4.186808e-06, 
    4.204028e-06, 4.209276e-06, 4.21147e-06,
  3.865609e-06, 3.902637e-06, 3.895425e-06, 3.925389e-06, 3.908754e-06, 
    3.928395e-06, 3.873102e-06, 3.90411e-06, 3.884301e-06, 3.868936e-06, 
    3.983859e-06, 3.926729e-06, 4.043637e-06, 4.006885e-06, 4.09952e-06, 
    4.037907e-06, 4.111999e-06, 4.097738e-06, 4.140738e-06, 4.128397e-06, 
    4.183635e-06, 4.146441e-06, 4.212411e-06, 4.174738e-06, 4.18062e-06, 
    4.145216e-06, 3.938195e-06, 3.976724e-06, 3.935917e-06, 3.941399e-06, 
    3.938939e-06, 3.909097e-06, 3.8941e-06, 3.862787e-06, 3.868462e-06, 
    3.891466e-06, 3.943865e-06, 3.92604e-06, 3.971041e-06, 3.970023e-06, 
    4.020411e-06, 3.997653e-06, 4.082811e-06, 4.058519e-06, 4.128912e-06, 
    4.111153e-06, 4.128077e-06, 4.122942e-06, 4.128144e-06, 4.102114e-06, 
    4.113256e-06, 4.090388e-06, 4.00191e-06, 4.027814e-06, 3.950797e-06, 
    3.904838e-06, 3.874459e-06, 3.852973e-06, 3.856007e-06, 3.861794e-06, 
    3.891601e-06, 3.919729e-06, 3.941231e-06, 3.955647e-06, 3.969876e-06, 
    4.013096e-06, 4.036067e-06, 4.087731e-06, 4.078385e-06, 4.094226e-06, 
    4.109389e-06, 4.134905e-06, 4.1307e-06, 4.141961e-06, 4.093808e-06, 
    4.125779e-06, 4.073066e-06, 4.08745e-06, 3.973745e-06, 3.930845e-06, 
    3.912677e-06, 3.896811e-06, 3.85834e-06, 3.884887e-06, 3.874412e-06, 
    3.899357e-06, 3.915249e-06, 3.907385e-06, 3.956041e-06, 3.93709e-06, 
    4.03743e-06, 3.994059e-06, 4.107618e-06, 4.080303e-06, 4.114179e-06, 
    4.096876e-06, 4.126545e-06, 4.099838e-06, 4.146156e-06, 4.156275e-06, 
    4.149359e-06, 4.175959e-06, 4.09836e-06, 4.128076e-06, 3.907165e-06, 
    3.908447e-06, 3.914422e-06, 3.88819e-06, 3.886588e-06, 3.862631e-06, 
    3.883945e-06, 3.893038e-06, 3.916171e-06, 3.929885e-06, 3.942944e-06, 
    3.97173e-06, 4.004001e-06, 4.049341e-06, 4.082071e-06, 4.104081e-06, 
    4.090578e-06, 4.102498e-06, 4.089174e-06, 4.082936e-06, 4.152482e-06, 
    4.11336e-06, 4.172128e-06, 4.168865e-06, 4.142229e-06, 4.169232e-06, 
    3.909347e-06, 3.901972e-06, 3.876419e-06, 3.896409e-06, 3.860026e-06, 
    3.880371e-06, 3.892093e-06, 3.937485e-06, 3.947493e-06, 3.956784e-06, 
    3.975165e-06, 3.998816e-06, 4.040472e-06, 4.076888e-06, 4.110271e-06, 
    4.107821e-06, 4.108684e-06, 4.116157e-06, 4.097656e-06, 4.119199e-06, 
    4.12282e-06, 4.113356e-06, 4.168428e-06, 4.152658e-06, 4.168796e-06, 
    4.158524e-06, 3.904369e-06, 3.916786e-06, 3.910074e-06, 3.9227e-06, 
    3.913803e-06, 3.953441e-06, 3.965365e-06, 4.021388e-06, 3.99835e-06, 
    4.035047e-06, 4.00207e-06, 4.007904e-06, 4.036246e-06, 4.003849e-06, 
    4.074875e-06, 4.026654e-06, 4.116448e-06, 4.068052e-06, 4.11949e-06, 
    4.110127e-06, 4.125636e-06, 4.13955e-06, 4.157087e-06, 4.18954e-06, 
    4.182015e-06, 4.209226e-06, 3.935333e-06, 3.951504e-06, 3.95008e-06, 
    3.967036e-06, 3.979599e-06, 4.006895e-06, 4.050865e-06, 4.034303e-06, 
    4.064734e-06, 4.070856e-06, 4.024635e-06, 4.052983e-06, 3.962346e-06, 
    3.976921e-06, 3.96824e-06, 3.936608e-06, 4.038116e-06, 3.985863e-06, 
    4.082613e-06, 4.054111e-06, 4.137564e-06, 4.095957e-06, 4.177874e-06, 
    4.213133e-06, 4.246452e-06, 4.285548e-06, 3.960345e-06, 3.949341e-06, 
    3.969055e-06, 3.996408e-06, 4.021872e-06, 4.055847e-06, 4.059331e-06, 
    4.065714e-06, 4.082271e-06, 4.096217e-06, 4.067733e-06, 4.099717e-06, 
    3.980304e-06, 4.042667e-06, 3.945184e-06, 3.974415e-06, 3.994794e-06, 
    3.985848e-06, 4.032412e-06, 4.043425e-06, 4.088329e-06, 4.065087e-06, 
    4.204417e-06, 4.142491e-06, 4.315435e-06, 4.266758e-06, 3.9455e-06, 
    3.960307e-06, 4.012054e-06, 3.987392e-06, 4.05812e-06, 4.075623e-06, 
    4.089879e-06, 4.108137e-06, 4.110112e-06, 4.120951e-06, 4.103196e-06, 
    4.120249e-06, 4.055919e-06, 4.084606e-06, 4.006123e-06, 4.025156e-06, 
    4.016395e-06, 4.006795e-06, 4.03646e-06, 4.06818e-06, 4.06886e-06, 
    4.079058e-06, 4.10786e-06, 4.058409e-06, 4.21244e-06, 4.116982e-06, 
    3.976485e-06, 4.005139e-06, 4.009241e-06, 3.998124e-06, 4.073866e-06, 
    4.046341e-06, 4.120686e-06, 4.100529e-06, 4.133582e-06, 4.117141e-06, 
    4.114725e-06, 4.093662e-06, 4.080574e-06, 4.047602e-06, 4.02087e-06, 
    3.999735e-06, 4.004645e-06, 4.027878e-06, 4.070125e-06, 4.110289e-06, 
    4.101475e-06, 4.131065e-06, 4.052972e-06, 4.085629e-06, 4.072991e-06, 
    4.105983e-06, 4.033863e-06, 4.095235e-06, 4.018249e-06, 4.02497e-06, 
    4.045796e-06, 4.087847e-06, 4.097181e-06, 4.107157e-06, 4.101e-06, 
    4.0712e-06, 4.066329e-06, 4.04529e-06, 4.039489e-06, 4.023506e-06, 
    4.010296e-06, 4.022364e-06, 4.035057e-06, 4.071213e-06, 4.103931e-06, 
    4.139747e-06, 4.148537e-06, 4.190618e-06, 4.156345e-06, 4.212975e-06, 
    4.164804e-06, 4.248363e-06, 4.098807e-06, 4.163392e-06, 4.046746e-06, 
    4.059234e-06, 4.081871e-06, 4.134021e-06, 4.105828e-06, 4.13881e-06, 
    4.066138e-06, 4.02868e-06, 4.019018e-06, 4.001019e-06, 4.01943e-06, 
    4.017931e-06, 4.035584e-06, 4.029907e-06, 4.072416e-06, 4.049555e-06, 
    4.114664e-06, 4.13855e-06, 4.20637e-06, 4.248211e-06, 4.291011e-06, 
    4.309972e-06, 4.315752e-06, 4.318169e-06,
  4.108354e-06, 4.14695e-06, 4.139431e-06, 4.170682e-06, 4.153329e-06, 
    4.173817e-06, 4.116162e-06, 4.148488e-06, 4.127834e-06, 4.111819e-06, 
    4.231721e-06, 4.172079e-06, 4.294188e-06, 4.255769e-06, 4.352662e-06, 
    4.288198e-06, 4.365729e-06, 4.350793e-06, 4.395833e-06, 4.382902e-06, 
    4.440811e-06, 4.401808e-06, 4.471002e-06, 4.431477e-06, 4.437647e-06, 
    4.400526e-06, 4.184041e-06, 4.224269e-06, 4.181664e-06, 4.187385e-06, 
    4.184817e-06, 4.153687e-06, 4.138052e-06, 4.105411e-06, 4.111326e-06, 
    4.135304e-06, 4.189959e-06, 4.171358e-06, 4.218326e-06, 4.217262e-06, 
    4.269903e-06, 4.246122e-06, 4.335169e-06, 4.30975e-06, 4.383441e-06, 
    4.36484e-06, 4.382567e-06, 4.377187e-06, 4.382637e-06, 4.355375e-06, 
    4.367043e-06, 4.343099e-06, 4.25057e-06, 4.277643e-06, 4.197193e-06, 
    4.149249e-06, 4.117576e-06, 4.095187e-06, 4.098348e-06, 4.104378e-06, 
    4.135445e-06, 4.164775e-06, 4.187209e-06, 4.202254e-06, 4.217109e-06, 
    4.262264e-06, 4.286273e-06, 4.34032e-06, 4.330536e-06, 4.347118e-06, 
    4.362992e-06, 4.389721e-06, 4.385315e-06, 4.397115e-06, 4.346679e-06, 
    4.380161e-06, 4.324969e-06, 4.340024e-06, 4.221159e-06, 4.176372e-06, 
    4.157424e-06, 4.140876e-06, 4.10078e-06, 4.128445e-06, 4.117527e-06, 
    4.143529e-06, 4.160102e-06, 4.1519e-06, 4.202666e-06, 4.182887e-06, 
    4.287698e-06, 4.242368e-06, 4.361139e-06, 4.332543e-06, 4.368009e-06, 
    4.34989e-06, 4.380963e-06, 4.352992e-06, 4.401511e-06, 4.412118e-06, 
    4.404868e-06, 4.432755e-06, 4.351445e-06, 4.382567e-06, 4.151671e-06, 
    4.153008e-06, 4.159239e-06, 4.131889e-06, 4.130218e-06, 4.105249e-06, 
    4.127462e-06, 4.136942e-06, 4.161063e-06, 4.17537e-06, 4.188996e-06, 
    4.219046e-06, 4.252756e-06, 4.300153e-06, 4.334393e-06, 4.357434e-06, 
    4.343297e-06, 4.355777e-06, 4.341828e-06, 4.335298e-06, 4.408143e-06, 
    4.367153e-06, 4.428738e-06, 4.425317e-06, 4.397396e-06, 4.425702e-06, 
    4.153947e-06, 4.146255e-06, 4.119619e-06, 4.140456e-06, 4.102536e-06, 
    4.123737e-06, 4.135958e-06, 4.183301e-06, 4.193744e-06, 4.203442e-06, 
    4.222633e-06, 4.247337e-06, 4.290877e-06, 4.32897e-06, 4.363917e-06, 
    4.36135e-06, 4.362254e-06, 4.370082e-06, 4.350708e-06, 4.373267e-06, 
    4.377061e-06, 4.367147e-06, 4.424859e-06, 4.408325e-06, 4.425244e-06, 
    4.414474e-06, 4.148755e-06, 4.161705e-06, 4.154704e-06, 4.167875e-06, 
    4.158594e-06, 4.199955e-06, 4.212402e-06, 4.270928e-06, 4.24685e-06, 
    4.285205e-06, 4.250737e-06, 4.256833e-06, 4.286463e-06, 4.252595e-06, 
    4.326866e-06, 4.276433e-06, 4.370386e-06, 4.31973e-06, 4.373572e-06, 
    4.363765e-06, 4.380009e-06, 4.394588e-06, 4.412968e-06, 4.447003e-06, 
    4.439108e-06, 4.467658e-06, 4.181054e-06, 4.197932e-06, 4.196443e-06, 
    4.214144e-06, 4.227263e-06, 4.255777e-06, 4.301745e-06, 4.284425e-06, 
    4.316252e-06, 4.322658e-06, 4.274317e-06, 4.303961e-06, 4.209249e-06, 
    4.224469e-06, 4.215402e-06, 4.182385e-06, 4.288414e-06, 4.233808e-06, 
    4.334961e-06, 4.30514e-06, 4.392507e-06, 4.348932e-06, 4.434766e-06, 
    4.471763e-06, 4.506743e-06, 4.547832e-06, 4.207159e-06, 4.195672e-06, 
    4.216252e-06, 4.244823e-06, 4.271431e-06, 4.306956e-06, 4.3106e-06, 
    4.317278e-06, 4.334603e-06, 4.3492e-06, 4.319392e-06, 4.352864e-06, 
    4.228007e-06, 4.293172e-06, 4.191335e-06, 4.221852e-06, 4.243136e-06, 
    4.233791e-06, 4.282448e-06, 4.293964e-06, 4.340945e-06, 4.316621e-06, 
    4.462616e-06, 4.397673e-06, 4.579261e-06, 4.52808e-06, 4.191663e-06, 
    4.207119e-06, 4.26117e-06, 4.235402e-06, 4.309333e-06, 4.327646e-06, 
    4.342566e-06, 4.361683e-06, 4.363749e-06, 4.375102e-06, 4.356507e-06, 
    4.374366e-06, 4.307032e-06, 4.337046e-06, 4.25497e-06, 4.274863e-06, 
    4.265704e-06, 4.255673e-06, 4.28668e-06, 4.31986e-06, 4.320569e-06, 
    4.331242e-06, 4.361402e-06, 4.309634e-06, 4.471042e-06, 4.370954e-06, 
    4.22401e-06, 4.253946e-06, 4.25823e-06, 4.246612e-06, 4.325808e-06, 
    4.297014e-06, 4.374825e-06, 4.353715e-06, 4.388334e-06, 4.371112e-06, 
    4.368581e-06, 4.346526e-06, 4.332827e-06, 4.298332e-06, 4.270384e-06, 
    4.248296e-06, 4.253426e-06, 4.27771e-06, 4.321895e-06, 4.363937e-06, 
    4.354707e-06, 4.385698e-06, 4.303948e-06, 4.338119e-06, 4.324894e-06, 
    4.359426e-06, 4.283966e-06, 4.348182e-06, 4.267642e-06, 4.274668e-06, 
    4.296444e-06, 4.340443e-06, 4.35021e-06, 4.360656e-06, 4.354208e-06, 
    4.323019e-06, 4.317921e-06, 4.295913e-06, 4.289849e-06, 4.273138e-06, 
    4.259331e-06, 4.271945e-06, 4.285216e-06, 4.323032e-06, 4.357279e-06, 
    4.394796e-06, 4.404005e-06, 4.448138e-06, 4.412196e-06, 4.471604e-06, 
    4.421071e-06, 4.508759e-06, 4.351918e-06, 4.419584e-06, 4.297436e-06, 
    4.310498e-06, 4.334187e-06, 4.388799e-06, 4.359264e-06, 4.393815e-06, 
    4.317721e-06, 4.27855e-06, 4.268446e-06, 4.249637e-06, 4.268877e-06, 
    4.26731e-06, 4.285764e-06, 4.279829e-06, 4.32429e-06, 4.300374e-06, 
    4.368518e-06, 4.393542e-06, 4.464662e-06, 4.508594e-06, 4.553571e-06, 
    4.573513e-06, 4.579593e-06, 4.582137e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.778234, 5.778215, 5.778219, 5.778203, 5.778212, 5.778202, 5.778231, 
    5.778214, 5.778225, 5.778233, 5.778173, 5.778203, 5.778142, 5.778162, 
    5.778114, 5.778146, 5.778108, 5.778115, 5.778093, 5.7781, 5.778072, 
    5.77809, 5.778057, 5.778076, 5.778073, 5.778091, 5.778197, 5.778177, 
    5.778198, 5.778195, 5.778196, 5.778212, 5.77822, 5.778236, 5.778233, 
    5.778221, 5.778194, 5.778203, 5.77818, 5.778181, 5.778154, 5.778166, 
    5.778123, 5.778135, 5.778099, 5.778108, 5.7781, 5.778102, 5.7781, 
    5.778113, 5.778107, 5.778119, 5.778164, 5.778151, 5.778191, 5.778214, 
    5.77823, 5.778241, 5.77824, 5.778237, 5.778221, 5.778206, 5.778195, 
    5.778188, 5.778181, 5.778158, 5.778147, 5.77812, 5.778125, 5.778117, 
    5.778109, 5.778096, 5.778099, 5.778093, 5.778117, 5.778101, 5.778128, 
    5.778121, 5.778179, 5.778201, 5.77821, 5.778218, 5.778238, 5.778224, 
    5.77823, 5.778217, 5.778209, 5.778213, 5.778188, 5.778197, 5.778146, 
    5.778168, 5.77811, 5.778124, 5.778107, 5.778116, 5.7781, 5.778114, 
    5.77809, 5.778085, 5.778089, 5.778076, 5.778115, 5.7781, 5.778213, 
    5.778213, 5.778209, 5.778223, 5.778224, 5.778236, 5.778225, 5.77822, 
    5.778208, 5.778201, 5.778194, 5.77818, 5.778163, 5.77814, 5.778123, 
    5.778112, 5.778119, 5.778113, 5.77812, 5.778122, 5.778088, 5.778107, 
    5.778078, 5.778079, 5.778092, 5.778079, 5.778212, 5.778216, 5.778229, 
    5.778219, 5.778238, 5.778227, 5.778221, 5.778197, 5.778192, 5.778187, 
    5.778178, 5.778166, 5.778144, 5.778126, 5.778109, 5.77811, 5.77811, 
    5.778106, 5.778115, 5.778104, 5.778102, 5.778107, 5.77808, 5.778087, 
    5.778079, 5.778084, 5.778214, 5.778208, 5.778212, 5.778205, 5.77821, 
    5.778189, 5.778183, 5.778154, 5.778166, 5.778147, 5.778164, 5.778161, 
    5.778146, 5.778163, 5.778127, 5.778152, 5.778106, 5.77813, 5.778104, 
    5.778109, 5.778101, 5.778094, 5.778085, 5.778069, 5.778072, 5.778059, 
    5.778198, 5.77819, 5.778191, 5.778182, 5.778175, 5.778162, 5.778139, 
    5.778147, 5.778132, 5.778129, 5.778152, 5.778138, 5.778184, 5.778177, 
    5.778182, 5.778198, 5.778145, 5.778172, 5.778123, 5.778137, 5.778095, 
    5.778116, 5.778075, 5.778057, 5.77804, 5.778021, 5.778185, 5.778191, 
    5.778181, 5.778167, 5.778154, 5.778136, 5.778135, 5.778131, 5.778123, 
    5.778116, 5.778131, 5.778114, 5.778175, 5.778143, 5.778193, 5.778178, 
    5.778168, 5.778172, 5.778149, 5.778143, 5.77812, 5.778132, 5.778061, 
    5.778092, 5.778006, 5.77803, 5.778193, 5.778185, 5.778159, 5.778172, 
    5.778135, 5.778126, 5.778119, 5.77811, 5.778109, 5.778103, 5.778112, 
    5.778104, 5.778136, 5.778122, 5.778162, 5.778152, 5.778157, 5.778162, 
    5.778146, 5.77813, 5.77813, 5.778125, 5.77811, 5.778135, 5.778057, 
    5.778105, 5.778177, 5.778162, 5.77816, 5.778166, 5.778127, 5.778141, 
    5.778103, 5.778114, 5.778097, 5.778105, 5.778107, 5.778117, 5.778124, 
    5.778141, 5.778154, 5.778165, 5.778162, 5.778151, 5.778129, 5.778109, 
    5.778113, 5.778098, 5.778138, 5.778121, 5.778128, 5.778111, 5.778148, 
    5.778116, 5.778156, 5.778152, 5.778141, 5.77812, 5.778115, 5.778111, 
    5.778113, 5.778129, 5.778131, 5.778142, 5.778145, 5.778153, 5.77816, 
    5.778153, 5.778147, 5.778129, 5.778112, 5.778094, 5.77809, 5.778068, 
    5.778085, 5.778057, 5.778081, 5.778039, 5.778115, 5.778082, 5.778141, 
    5.778135, 5.778123, 5.778097, 5.778111, 5.778094, 5.778131, 5.778151, 
    5.778155, 5.778164, 5.778155, 5.778156, 5.778147, 5.77815, 5.778128, 
    5.77814, 5.778107, 5.778094, 5.77806, 5.778039, 5.778018, 5.778008, 
    5.778006, 5.778005 ;

 SOIL1C_TO_SOIL2C =
  3.09861e-08, 3.112362e-08, 3.109689e-08, 3.12078e-08, 3.114627e-08, 
    3.12189e-08, 3.101398e-08, 3.112907e-08, 3.10556e-08, 3.099848e-08, 
    3.142307e-08, 3.121275e-08, 3.164162e-08, 3.150745e-08, 3.184453e-08, 
    3.162074e-08, 3.188966e-08, 3.183808e-08, 3.199334e-08, 3.194886e-08, 
    3.214746e-08, 3.201388e-08, 3.225043e-08, 3.211556e-08, 3.213665e-08, 
    3.200947e-08, 3.125508e-08, 3.139689e-08, 3.124668e-08, 3.12669e-08, 
    3.125783e-08, 3.114754e-08, 3.109196e-08, 3.09756e-08, 3.099672e-08, 
    3.108219e-08, 3.127599e-08, 3.121021e-08, 3.137602e-08, 3.137228e-08, 
    3.15569e-08, 3.147365e-08, 3.1784e-08, 3.169579e-08, 3.195072e-08, 
    3.18866e-08, 3.19477e-08, 3.192918e-08, 3.194794e-08, 3.185391e-08, 
    3.18942e-08, 3.181146e-08, 3.148924e-08, 3.158393e-08, 3.130154e-08, 
    3.113177e-08, 3.101903e-08, 3.093903e-08, 3.095034e-08, 3.09719e-08, 
    3.10827e-08, 3.118688e-08, 3.126629e-08, 3.13194e-08, 3.137174e-08, 
    3.153016e-08, 3.161403e-08, 3.180183e-08, 3.176795e-08, 3.182536e-08, 
    3.188022e-08, 3.197232e-08, 3.195717e-08, 3.199774e-08, 3.182385e-08, 
    3.193941e-08, 3.174864e-08, 3.180082e-08, 3.138594e-08, 3.122796e-08, 
    3.116079e-08, 3.110202e-08, 3.095903e-08, 3.105777e-08, 3.101885e-08, 
    3.111146e-08, 3.117031e-08, 3.114121e-08, 3.132086e-08, 3.125101e-08, 
    3.1619e-08, 3.146048e-08, 3.187382e-08, 3.17749e-08, 3.189754e-08, 
    3.183496e-08, 3.194218e-08, 3.184568e-08, 3.201285e-08, 3.204925e-08, 
    3.202437e-08, 3.211994e-08, 3.184033e-08, 3.19477e-08, 3.114039e-08, 
    3.114513e-08, 3.116725e-08, 3.107004e-08, 3.106409e-08, 3.097502e-08, 
    3.105428e-08, 3.108803e-08, 3.117372e-08, 3.122441e-08, 3.12726e-08, 
    3.137855e-08, 3.149689e-08, 3.16624e-08, 3.178132e-08, 3.186103e-08, 
    3.181215e-08, 3.18553e-08, 3.180706e-08, 3.178445e-08, 3.203561e-08, 
    3.189458e-08, 3.21062e-08, 3.209449e-08, 3.199871e-08, 3.209581e-08, 
    3.114847e-08, 3.112115e-08, 3.102631e-08, 3.110053e-08, 3.096531e-08, 
    3.1041e-08, 3.108452e-08, 3.125246e-08, 3.128937e-08, 3.132359e-08, 
    3.139117e-08, 3.147791e-08, 3.163009e-08, 3.176251e-08, 3.188341e-08, 
    3.187456e-08, 3.187768e-08, 3.190468e-08, 3.183778e-08, 3.191566e-08, 
    3.192874e-08, 3.189456e-08, 3.209292e-08, 3.203624e-08, 3.209423e-08, 
    3.205734e-08, 3.113004e-08, 3.1176e-08, 3.115116e-08, 3.119786e-08, 
    3.116496e-08, 3.131128e-08, 3.135515e-08, 3.156046e-08, 3.14762e-08, 
    3.161031e-08, 3.148983e-08, 3.151117e-08, 3.161468e-08, 3.149634e-08, 
    3.17552e-08, 3.157969e-08, 3.190573e-08, 3.173043e-08, 3.191672e-08, 
    3.188289e-08, 3.19389e-08, 3.198906e-08, 3.205217e-08, 3.216862e-08, 
    3.214166e-08, 3.223905e-08, 3.124453e-08, 3.130415e-08, 3.12989e-08, 
    3.13613e-08, 3.140745e-08, 3.150749e-08, 3.166794e-08, 3.16076e-08, 
    3.171838e-08, 3.174062e-08, 3.157232e-08, 3.167565e-08, 3.134405e-08, 
    3.139762e-08, 3.136573e-08, 3.124923e-08, 3.16215e-08, 3.143043e-08, 
    3.178328e-08, 3.167976e-08, 3.198191e-08, 3.183163e-08, 3.212681e-08, 
    3.225301e-08, 3.237181e-08, 3.251063e-08, 3.133669e-08, 3.129618e-08, 
    3.136872e-08, 3.146909e-08, 3.156223e-08, 3.168607e-08, 3.169874e-08, 
    3.172194e-08, 3.178204e-08, 3.183257e-08, 3.172927e-08, 3.184524e-08, 
    3.141003e-08, 3.163809e-08, 3.128086e-08, 3.138841e-08, 3.146317e-08, 
    3.143038e-08, 3.160071e-08, 3.164085e-08, 3.1804e-08, 3.171966e-08, 
    3.222186e-08, 3.199965e-08, 3.261636e-08, 3.244399e-08, 3.128202e-08, 
    3.133655e-08, 3.152635e-08, 3.143604e-08, 3.169434e-08, 3.175792e-08, 
    3.180962e-08, 3.18757e-08, 3.188283e-08, 3.192199e-08, 3.185783e-08, 
    3.191946e-08, 3.168633e-08, 3.179051e-08, 3.150466e-08, 3.157422e-08, 
    3.154222e-08, 3.150712e-08, 3.161547e-08, 3.17309e-08, 3.173337e-08, 
    3.177039e-08, 3.187468e-08, 3.169539e-08, 3.225052e-08, 3.190765e-08, 
    3.139602e-08, 3.150106e-08, 3.151607e-08, 3.147538e-08, 3.175155e-08, 
    3.165147e-08, 3.192104e-08, 3.184818e-08, 3.196756e-08, 3.190824e-08, 
    3.189951e-08, 3.182332e-08, 3.177589e-08, 3.165606e-08, 3.155857e-08, 
    3.148128e-08, 3.149925e-08, 3.158416e-08, 3.173796e-08, 3.188348e-08, 
    3.18516e-08, 3.195848e-08, 3.167561e-08, 3.179421e-08, 3.174837e-08, 
    3.186791e-08, 3.1606e-08, 3.1829e-08, 3.1549e-08, 3.157355e-08, 
    3.164949e-08, 3.180225e-08, 3.183606e-08, 3.187215e-08, 3.184988e-08, 
    3.174187e-08, 3.172417e-08, 3.164764e-08, 3.162651e-08, 3.15682e-08, 
    3.151993e-08, 3.156403e-08, 3.161035e-08, 3.174192e-08, 3.186049e-08, 
    3.198977e-08, 3.202142e-08, 3.217248e-08, 3.20495e-08, 3.225243e-08, 
    3.207989e-08, 3.23786e-08, 3.184194e-08, 3.207482e-08, 3.165295e-08, 
    3.169839e-08, 3.178059e-08, 3.196913e-08, 3.186735e-08, 3.198639e-08, 
    3.172348e-08, 3.158709e-08, 3.155181e-08, 3.148598e-08, 3.155331e-08, 
    3.154784e-08, 3.161227e-08, 3.159157e-08, 3.174628e-08, 3.166318e-08, 
    3.189929e-08, 3.198545e-08, 3.222884e-08, 3.237806e-08, 3.252999e-08, 
    3.259706e-08, 3.261748e-08, 3.262602e-08 ;

 SOIL1C_TO_SOIL3C =
  3.675195e-10, 3.691511e-10, 3.688339e-10, 3.7015e-10, 3.694199e-10, 
    3.702817e-10, 3.678503e-10, 3.692158e-10, 3.683441e-10, 3.676664e-10, 
    3.727043e-10, 3.702087e-10, 3.752973e-10, 3.737054e-10, 3.77705e-10, 
    3.750496e-10, 3.782405e-10, 3.776285e-10, 3.794708e-10, 3.78943e-10, 
    3.812996e-10, 3.797145e-10, 3.825215e-10, 3.809211e-10, 3.811714e-10, 
    3.796622e-10, 3.70711e-10, 3.723935e-10, 3.706113e-10, 3.708512e-10, 
    3.707435e-10, 3.69435e-10, 3.687755e-10, 3.673948e-10, 3.676455e-10, 
    3.686596e-10, 3.709591e-10, 3.701785e-10, 3.72146e-10, 3.721015e-10, 
    3.742921e-10, 3.733044e-10, 3.769868e-10, 3.759401e-10, 3.789651e-10, 
    3.782042e-10, 3.789293e-10, 3.787095e-10, 3.789322e-10, 3.778164e-10, 
    3.782944e-10, 3.773127e-10, 3.734893e-10, 3.746128e-10, 3.712622e-10, 
    3.692478e-10, 3.679101e-10, 3.66961e-10, 3.670952e-10, 3.673509e-10, 
    3.686656e-10, 3.699017e-10, 3.708439e-10, 3.714741e-10, 3.720952e-10, 
    3.739748e-10, 3.7497e-10, 3.771984e-10, 3.767963e-10, 3.774776e-10, 
    3.781286e-10, 3.792214e-10, 3.790416e-10, 3.795231e-10, 3.774597e-10, 
    3.788309e-10, 3.765673e-10, 3.771864e-10, 3.722637e-10, 3.703891e-10, 
    3.695922e-10, 3.688949e-10, 3.671983e-10, 3.683699e-10, 3.67908e-10, 
    3.690069e-10, 3.697051e-10, 3.693598e-10, 3.714914e-10, 3.706626e-10, 
    3.75029e-10, 3.731481e-10, 3.780526e-10, 3.768789e-10, 3.78334e-10, 
    3.775915e-10, 3.788637e-10, 3.777187e-10, 3.797023e-10, 3.801342e-10, 
    3.798391e-10, 3.809731e-10, 3.776552e-10, 3.789293e-10, 3.693501e-10, 
    3.694064e-10, 3.696688e-10, 3.685154e-10, 3.684448e-10, 3.673879e-10, 
    3.683284e-10, 3.687289e-10, 3.697457e-10, 3.703471e-10, 3.709188e-10, 
    3.72176e-10, 3.735801e-10, 3.755439e-10, 3.769549e-10, 3.779008e-10, 
    3.773209e-10, 3.778329e-10, 3.772605e-10, 3.769922e-10, 3.799724e-10, 
    3.782989e-10, 3.808099e-10, 3.80671e-10, 3.795345e-10, 3.806866e-10, 
    3.69446e-10, 3.691219e-10, 3.679966e-10, 3.688772e-10, 3.672729e-10, 
    3.681708e-10, 3.686872e-10, 3.706799e-10, 3.711178e-10, 3.715238e-10, 
    3.723257e-10, 3.733549e-10, 3.751606e-10, 3.767318e-10, 3.781664e-10, 
    3.780613e-10, 3.780983e-10, 3.784188e-10, 3.77625e-10, 3.785491e-10, 
    3.787042e-10, 3.782987e-10, 3.806524e-10, 3.799799e-10, 3.806681e-10, 
    3.802302e-10, 3.692273e-10, 3.697726e-10, 3.694779e-10, 3.700321e-10, 
    3.696417e-10, 3.713777e-10, 3.718983e-10, 3.743344e-10, 3.733347e-10, 
    3.749259e-10, 3.734963e-10, 3.737496e-10, 3.749777e-10, 3.735736e-10, 
    3.766451e-10, 3.745625e-10, 3.784312e-10, 3.763512e-10, 3.785616e-10, 
    3.781603e-10, 3.788248e-10, 3.7942e-10, 3.801689e-10, 3.815507e-10, 
    3.812307e-10, 3.823865e-10, 3.705857e-10, 3.712931e-10, 3.712309e-10, 
    3.719713e-10, 3.725188e-10, 3.737058e-10, 3.756097e-10, 3.748938e-10, 
    3.762082e-10, 3.764721e-10, 3.744751e-10, 3.757012e-10, 3.717666e-10, 
    3.724022e-10, 3.720238e-10, 3.706415e-10, 3.750586e-10, 3.727915e-10, 
    3.769783e-10, 3.757499e-10, 3.793351e-10, 3.77552e-10, 3.810546e-10, 
    3.82552e-10, 3.839618e-10, 3.856091e-10, 3.716793e-10, 3.711986e-10, 
    3.720594e-10, 3.732502e-10, 3.743554e-10, 3.758248e-10, 3.759752e-10, 
    3.762504e-10, 3.769636e-10, 3.775632e-10, 3.763375e-10, 3.777135e-10, 
    3.725495e-10, 3.752555e-10, 3.710168e-10, 3.722929e-10, 3.7318e-10, 
    3.72791e-10, 3.748119e-10, 3.752883e-10, 3.772241e-10, 3.762234e-10, 
    3.821824e-10, 3.795457e-10, 3.868637e-10, 3.848183e-10, 3.710306e-10, 
    3.716776e-10, 3.739297e-10, 3.728581e-10, 3.759229e-10, 3.766774e-10, 
    3.772908e-10, 3.780749e-10, 3.781596e-10, 3.786242e-10, 3.778629e-10, 
    3.785941e-10, 3.758279e-10, 3.77064e-10, 3.736723e-10, 3.744977e-10, 
    3.74118e-10, 3.737015e-10, 3.749871e-10, 3.763567e-10, 3.763861e-10, 
    3.768253e-10, 3.780628e-10, 3.759354e-10, 3.825226e-10, 3.78454e-10, 
    3.723832e-10, 3.736295e-10, 3.738077e-10, 3.733248e-10, 3.766017e-10, 
    3.754143e-10, 3.786128e-10, 3.777484e-10, 3.791649e-10, 3.78461e-10, 
    3.783574e-10, 3.774534e-10, 3.768905e-10, 3.754687e-10, 3.74312e-10, 
    3.733949e-10, 3.736081e-10, 3.746156e-10, 3.764405e-10, 3.781672e-10, 
    3.777889e-10, 3.790572e-10, 3.757007e-10, 3.77108e-10, 3.76564e-10, 
    3.779825e-10, 3.748747e-10, 3.775208e-10, 3.741984e-10, 3.744897e-10, 
    3.753907e-10, 3.772034e-10, 3.776046e-10, 3.780328e-10, 3.777686e-10, 
    3.764869e-10, 3.762769e-10, 3.753689e-10, 3.751181e-10, 3.744263e-10, 
    3.738534e-10, 3.743768e-10, 3.749264e-10, 3.764875e-10, 3.778944e-10, 
    3.794285e-10, 3.79804e-10, 3.815964e-10, 3.801372e-10, 3.825452e-10, 
    3.804977e-10, 3.840424e-10, 3.776744e-10, 3.804377e-10, 3.754318e-10, 
    3.75971e-10, 3.769463e-10, 3.791836e-10, 3.779758e-10, 3.793884e-10, 
    3.762687e-10, 3.746503e-10, 3.742317e-10, 3.734506e-10, 3.742496e-10, 
    3.741846e-10, 3.749492e-10, 3.747035e-10, 3.765393e-10, 3.755532e-10, 
    3.783548e-10, 3.793773e-10, 3.822653e-10, 3.84036e-10, 3.858388e-10, 
    3.866348e-10, 3.86877e-10, 3.869783e-10 ;

 SOIL1C_vr =
  19.98094, 19.98089, 19.9809, 19.98086, 19.98088, 19.98086, 19.98093, 
    19.98089, 19.98092, 19.98094, 19.98078, 19.98086, 19.9807, 19.98075, 
    19.98062, 19.9807, 19.9806, 19.98062, 19.98056, 19.98058, 19.9805, 
    19.98055, 19.98047, 19.98052, 19.98051, 19.98056, 19.98084, 19.98079, 
    19.98084, 19.98084, 19.98084, 19.98088, 19.9809, 19.98095, 19.98094, 
    19.98091, 19.98083, 19.98086, 19.9808, 19.9808, 19.98073, 19.98076, 
    19.98064, 19.98067, 19.98058, 19.9806, 19.98058, 19.98059, 19.98058, 
    19.98062, 19.9806, 19.98063, 19.98075, 19.98072, 19.98082, 19.98089, 
    19.98093, 19.98096, 19.98096, 19.98095, 19.98091, 19.98087, 19.98084, 
    19.98082, 19.9808, 19.98074, 19.98071, 19.98063, 19.98065, 19.98063, 
    19.98061, 19.98057, 19.98058, 19.98056, 19.98063, 19.98058, 19.98066, 
    19.98063, 19.98079, 19.98085, 19.98088, 19.9809, 19.98095, 19.98092, 
    19.98093, 19.9809, 19.98087, 19.98088, 19.98082, 19.98084, 19.9807, 
    19.98076, 19.98061, 19.98065, 19.9806, 19.98062, 19.98058, 19.98062, 
    19.98056, 19.98054, 19.98055, 19.98052, 19.98062, 19.98058, 19.98088, 
    19.98088, 19.98088, 19.98091, 19.98092, 19.98095, 19.98092, 19.98091, 
    19.98087, 19.98085, 19.98083, 19.98079, 19.98075, 19.98069, 19.98064, 
    19.98061, 19.98063, 19.98062, 19.98063, 19.98064, 19.98055, 19.9806, 
    19.98052, 19.98053, 19.98056, 19.98052, 19.98088, 19.98089, 19.98093, 
    19.9809, 19.98095, 19.98092, 19.98091, 19.98084, 19.98083, 19.98082, 
    19.98079, 19.98076, 19.9807, 19.98065, 19.9806, 19.98061, 19.98061, 
    19.9806, 19.98062, 19.98059, 19.98059, 19.9806, 19.98053, 19.98055, 
    19.98053, 19.98054, 19.98089, 19.98087, 19.98088, 19.98086, 19.98088, 
    19.98082, 19.9808, 19.98073, 19.98076, 19.98071, 19.98075, 19.98075, 
    19.98071, 19.98075, 19.98065, 19.98072, 19.9806, 19.98066, 19.98059, 
    19.9806, 19.98058, 19.98056, 19.98054, 19.9805, 19.98051, 19.98047, 
    19.98085, 19.98082, 19.98083, 19.9808, 19.98078, 19.98075, 19.98069, 
    19.98071, 19.98067, 19.98066, 19.98072, 19.98068, 19.98081, 19.98079, 
    19.9808, 19.98084, 19.9807, 19.98078, 19.98064, 19.98068, 19.98057, 
    19.98062, 19.98051, 19.98046, 19.98042, 19.98037, 19.98081, 19.98083, 
    19.9808, 19.98076, 19.98073, 19.98068, 19.98067, 19.98067, 19.98064, 
    19.98062, 19.98066, 19.98062, 19.98078, 19.9807, 19.98083, 19.98079, 
    19.98076, 19.98078, 19.98071, 19.9807, 19.98063, 19.98067, 19.98048, 
    19.98056, 19.98033, 19.98039, 19.98083, 19.98081, 19.98074, 19.98077, 
    19.98068, 19.98065, 19.98063, 19.98061, 19.9806, 19.98059, 19.98061, 
    19.98059, 19.98068, 19.98064, 19.98075, 19.98072, 19.98073, 19.98075, 
    19.98071, 19.98066, 19.98066, 19.98065, 19.98061, 19.98067, 19.98047, 
    19.98059, 19.98079, 19.98075, 19.98074, 19.98076, 19.98065, 19.98069, 
    19.98059, 19.98062, 19.98057, 19.98059, 19.9806, 19.98063, 19.98064, 
    19.98069, 19.98073, 19.98076, 19.98075, 19.98072, 19.98066, 19.9806, 
    19.98062, 19.98058, 19.98068, 19.98064, 19.98066, 19.98061, 19.98071, 
    19.98063, 19.98073, 19.98072, 19.98069, 19.98063, 19.98062, 19.98061, 
    19.98062, 19.98066, 19.98067, 19.98069, 19.9807, 19.98072, 19.98074, 
    19.98072, 19.98071, 19.98066, 19.98061, 19.98056, 19.98055, 19.9805, 
    19.98054, 19.98046, 19.98053, 19.98042, 19.98062, 19.98053, 19.98069, 
    19.98067, 19.98064, 19.98057, 19.98061, 19.98057, 19.98067, 19.98072, 
    19.98073, 19.98075, 19.98073, 19.98073, 19.98071, 19.98071, 19.98066, 
    19.98069, 19.9806, 19.98057, 19.98047, 19.98042, 19.98036, 19.98034, 
    19.98033, 19.98033,
  19.98318, 19.98312, 19.98313, 19.98308, 19.9831, 19.98307, 19.98317, 
    19.98311, 19.98315, 19.98317, 19.98298, 19.98307, 19.98287, 19.98294, 
    19.98278, 19.98288, 19.98276, 19.98278, 19.98271, 19.98273, 19.98264, 
    19.9827, 19.98259, 19.98265, 19.98264, 19.9827, 19.98305, 19.98299, 
    19.98306, 19.98305, 19.98305, 19.9831, 19.98313, 19.98318, 19.98318, 
    19.98314, 19.98304, 19.98307, 19.983, 19.983, 19.98291, 19.98295, 
    19.98281, 19.98285, 19.98273, 19.98276, 19.98273, 19.98274, 19.98273, 
    19.98277, 19.98276, 19.98279, 19.98294, 19.9829, 19.98303, 19.98311, 
    19.98316, 19.9832, 19.9832, 19.98319, 19.98314, 19.98309, 19.98305, 
    19.98302, 19.983, 19.98293, 19.98289, 19.9828, 19.98281, 19.98279, 
    19.98276, 19.98272, 19.98273, 19.98271, 19.98279, 19.98273, 19.98282, 
    19.9828, 19.98299, 19.98307, 19.9831, 19.98313, 19.98319, 19.98315, 
    19.98316, 19.98312, 19.98309, 19.98311, 19.98302, 19.98306, 19.98288, 
    19.98296, 19.98277, 19.98281, 19.98275, 19.98278, 19.98273, 19.98278, 
    19.9827, 19.98268, 19.98269, 19.98265, 19.98278, 19.98273, 19.98311, 
    19.9831, 19.9831, 19.98314, 19.98314, 19.98318, 19.98315, 19.98313, 
    19.98309, 19.98307, 19.98305, 19.983, 19.98294, 19.98286, 19.98281, 
    19.98277, 19.98279, 19.98277, 19.9828, 19.98281, 19.98269, 19.98276, 
    19.98266, 19.98266, 19.98271, 19.98266, 19.9831, 19.98312, 19.98316, 
    19.98313, 19.98319, 19.98315, 19.98313, 19.98306, 19.98304, 19.98302, 
    19.98299, 19.98295, 19.98288, 19.98282, 19.98276, 19.98277, 19.98276, 
    19.98275, 19.98278, 19.98275, 19.98274, 19.98276, 19.98266, 19.98269, 
    19.98266, 19.98268, 19.98311, 19.98309, 19.9831, 19.98308, 19.9831, 
    19.98303, 19.98301, 19.98291, 19.98295, 19.98289, 19.98294, 19.98293, 
    19.98289, 19.98294, 19.98282, 19.9829, 19.98275, 19.98283, 19.98275, 
    19.98276, 19.98273, 19.98271, 19.98268, 19.98263, 19.98264, 19.9826, 
    19.98306, 19.98303, 19.98303, 19.983, 19.98298, 19.98294, 19.98286, 
    19.98289, 19.98284, 19.98283, 19.98291, 19.98286, 19.98301, 19.98299, 
    19.983, 19.98306, 19.98288, 19.98297, 19.98281, 19.98286, 19.98272, 
    19.98278, 19.98265, 19.98259, 19.98253, 19.98247, 19.98302, 19.98303, 
    19.983, 19.98295, 19.98291, 19.98285, 19.98285, 19.98284, 19.98281, 
    19.98278, 19.98283, 19.98278, 19.98298, 19.98288, 19.98304, 19.98299, 
    19.98296, 19.98297, 19.98289, 19.98287, 19.9828, 19.98284, 19.9826, 
    19.98271, 19.98242, 19.9825, 19.98304, 19.98302, 19.98293, 19.98297, 
    19.98285, 19.98282, 19.9828, 19.98277, 19.98276, 19.98274, 19.98277, 
    19.98274, 19.98285, 19.98281, 19.98294, 19.9829, 19.98292, 19.98294, 
    19.98289, 19.98283, 19.98283, 19.98281, 19.98277, 19.98285, 19.98259, 
    19.98275, 19.98299, 19.98294, 19.98293, 19.98295, 19.98282, 19.98287, 
    19.98274, 19.98278, 19.98272, 19.98275, 19.98275, 19.98279, 19.98281, 
    19.98287, 19.98291, 19.98295, 19.98294, 19.9829, 19.98283, 19.98276, 
    19.98278, 19.98273, 19.98286, 19.9828, 19.98282, 19.98277, 19.98289, 
    19.98279, 19.98292, 19.98291, 19.98287, 19.9828, 19.98278, 19.98277, 
    19.98278, 19.98283, 19.98284, 19.98287, 19.98288, 19.98291, 19.98293, 
    19.98291, 19.98289, 19.98283, 19.98277, 19.98271, 19.9827, 19.98263, 
    19.98268, 19.98259, 19.98267, 19.98253, 19.98278, 19.98267, 19.98287, 
    19.98285, 19.98281, 19.98272, 19.98277, 19.98271, 19.98284, 19.9829, 
    19.98292, 19.98295, 19.98291, 19.98292, 19.98289, 19.9829, 19.98282, 
    19.98286, 19.98275, 19.98271, 19.9826, 19.98253, 19.98246, 19.98243, 
    19.98242, 19.98242,
  19.98421, 19.98414, 19.98416, 19.9841, 19.98413, 19.98409, 19.9842, 
    19.98414, 19.98418, 19.98421, 19.98399, 19.9841, 19.98388, 19.98395, 
    19.98377, 19.98389, 19.98375, 19.98378, 19.9837, 19.98372, 19.98362, 
    19.98369, 19.98357, 19.98364, 19.98363, 19.98369, 19.98408, 19.984, 
    19.98408, 19.98407, 19.98407, 19.98413, 19.98416, 19.98422, 19.98421, 
    19.98416, 19.98406, 19.9841, 19.98401, 19.98401, 19.98392, 19.98396, 
    19.9838, 19.98385, 19.98372, 19.98375, 19.98372, 19.98373, 19.98372, 
    19.98377, 19.98375, 19.98379, 19.98396, 19.98391, 19.98405, 19.98414, 
    19.9842, 19.98424, 19.98423, 19.98422, 19.98416, 19.98411, 19.98407, 
    19.98404, 19.98402, 19.98393, 19.98389, 19.9838, 19.98381, 19.98378, 
    19.98376, 19.98371, 19.98372, 19.9837, 19.98379, 19.98373, 19.98382, 
    19.9838, 19.98401, 19.98409, 19.98412, 19.98415, 19.98423, 19.98418, 
    19.9842, 19.98415, 19.98412, 19.98413, 19.98404, 19.98408, 19.98389, 
    19.98397, 19.98376, 19.98381, 19.98375, 19.98378, 19.98372, 19.98377, 
    19.98369, 19.98367, 19.98368, 19.98363, 19.98378, 19.98372, 19.98413, 
    19.98413, 19.98412, 19.98417, 19.98417, 19.98422, 19.98418, 19.98416, 
    19.98412, 19.98409, 19.98407, 19.98401, 19.98395, 19.98387, 19.98381, 
    19.98377, 19.98379, 19.98377, 19.98379, 19.9838, 19.98368, 19.98375, 
    19.98364, 19.98365, 19.9837, 19.98365, 19.98413, 19.98414, 19.98419, 
    19.98415, 19.98422, 19.98418, 19.98416, 19.98408, 19.98406, 19.98404, 
    19.984, 19.98396, 19.98388, 19.98382, 19.98376, 19.98376, 19.98376, 
    19.98374, 19.98378, 19.98374, 19.98373, 19.98375, 19.98365, 19.98368, 
    19.98365, 19.98367, 19.98414, 19.98412, 19.98413, 19.9841, 19.98412, 
    19.98405, 19.98402, 19.98392, 19.98396, 19.98389, 19.98396, 19.98394, 
    19.98389, 19.98395, 19.98382, 19.98391, 19.98374, 19.98383, 19.98374, 
    19.98376, 19.98373, 19.9837, 19.98367, 19.98361, 19.98362, 19.98357, 
    19.98408, 19.98405, 19.98405, 19.98402, 19.984, 19.98395, 19.98386, 
    19.98389, 19.98384, 19.98383, 19.98391, 19.98386, 19.98403, 19.984, 
    19.98402, 19.98408, 19.98389, 19.98399, 19.9838, 19.98386, 19.9837, 
    19.98378, 19.98363, 19.98357, 19.98351, 19.98343, 19.98403, 19.98405, 
    19.98402, 19.98396, 19.98392, 19.98385, 19.98385, 19.98384, 19.98381, 
    19.98378, 19.98383, 19.98377, 19.984, 19.98388, 19.98406, 19.98401, 
    19.98397, 19.98399, 19.9839, 19.98388, 19.9838, 19.98384, 19.98358, 
    19.9837, 19.98338, 19.98347, 19.98406, 19.98403, 19.98394, 19.98398, 
    19.98385, 19.98382, 19.98379, 19.98376, 19.98376, 19.98373, 19.98377, 
    19.98374, 19.98385, 19.9838, 19.98395, 19.98391, 19.98393, 19.98395, 
    19.98389, 19.98383, 19.98383, 19.98381, 19.98376, 19.98385, 19.98357, 
    19.98374, 19.984, 19.98395, 19.98394, 19.98396, 19.98382, 19.98387, 
    19.98374, 19.98377, 19.98371, 19.98374, 19.98375, 19.98379, 19.98381, 
    19.98387, 19.98392, 19.98396, 19.98395, 19.98391, 19.98383, 19.98376, 
    19.98377, 19.98372, 19.98386, 19.9838, 19.98382, 19.98376, 19.9839, 
    19.98378, 19.98392, 19.98391, 19.98387, 19.9838, 19.98378, 19.98376, 
    19.98377, 19.98383, 19.98384, 19.98388, 19.98388, 19.98392, 19.98394, 
    19.98392, 19.98389, 19.98383, 19.98377, 19.9837, 19.98368, 19.98361, 
    19.98367, 19.98357, 19.98365, 19.9835, 19.98378, 19.98366, 19.98387, 
    19.98385, 19.98381, 19.98371, 19.98376, 19.9837, 19.98384, 19.98391, 
    19.98392, 19.98396, 19.98392, 19.98392, 19.98389, 19.9839, 19.98382, 
    19.98387, 19.98375, 19.9837, 19.98358, 19.9835, 19.98343, 19.98339, 
    19.98338, 19.98338,
  19.98501, 19.98494, 19.98495, 19.98489, 19.98492, 19.98489, 19.98499, 
    19.98493, 19.98497, 19.985, 19.98478, 19.98489, 19.98467, 19.98474, 
    19.98456, 19.98468, 19.98454, 19.98456, 19.98448, 19.98451, 19.9844, 
    19.98447, 19.98435, 19.98442, 19.98441, 19.98447, 19.98487, 19.98479, 
    19.98487, 19.98486, 19.98487, 19.98492, 19.98495, 19.98501, 19.985, 
    19.98496, 19.98486, 19.98489, 19.9848, 19.98481, 19.98471, 19.98475, 
    19.98459, 19.98464, 19.9845, 19.98454, 19.98451, 19.98452, 19.98451, 
    19.98456, 19.98454, 19.98458, 19.98475, 19.9847, 19.98484, 19.98493, 
    19.98499, 19.98503, 19.98503, 19.98501, 19.98496, 19.9849, 19.98486, 
    19.98483, 19.98481, 19.98472, 19.98468, 19.98458, 19.9846, 19.98457, 
    19.98454, 19.98449, 19.9845, 19.98448, 19.98457, 19.98451, 19.98461, 
    19.98458, 19.9848, 19.98488, 19.98492, 19.98495, 19.98502, 19.98497, 
    19.98499, 19.98494, 19.98491, 19.98493, 19.98483, 19.98487, 19.98468, 
    19.98476, 19.98454, 19.9846, 19.98453, 19.98457, 19.98451, 19.98456, 
    19.98447, 19.98445, 19.98447, 19.98442, 19.98456, 19.98451, 19.98493, 
    19.98492, 19.98491, 19.98496, 19.98497, 19.98501, 19.98497, 19.98495, 
    19.98491, 19.98488, 19.98486, 19.9848, 19.98474, 19.98466, 19.98459, 
    19.98455, 19.98458, 19.98455, 19.98458, 19.98459, 19.98446, 19.98454, 
    19.98442, 19.98443, 19.98448, 19.98443, 19.98492, 19.98494, 19.98499, 
    19.98495, 19.98502, 19.98498, 19.98496, 19.98487, 19.98485, 19.98483, 
    19.9848, 19.98475, 19.98467, 19.9846, 19.98454, 19.98454, 19.98454, 
    19.98453, 19.98456, 19.98452, 19.98452, 19.98454, 19.98443, 19.98446, 
    19.98443, 19.98445, 19.98493, 19.98491, 19.98492, 19.9849, 19.98491, 
    19.98484, 19.98482, 19.98471, 19.98475, 19.98468, 19.98475, 19.98473, 
    19.98468, 19.98474, 19.98461, 19.9847, 19.98453, 19.98462, 19.98452, 
    19.98454, 19.98451, 19.98449, 19.98445, 19.98439, 19.98441, 19.98436, 
    19.98487, 19.98484, 19.98484, 19.98481, 19.98479, 19.98474, 19.98465, 
    19.98468, 19.98463, 19.98462, 19.9847, 19.98465, 19.98482, 19.98479, 
    19.98481, 19.98487, 19.98468, 19.98478, 19.98459, 19.98465, 19.98449, 
    19.98457, 19.98441, 19.98435, 19.98429, 19.98421, 19.98483, 19.98485, 
    19.98481, 19.98476, 19.98471, 19.98464, 19.98464, 19.98462, 19.98459, 
    19.98457, 19.98462, 19.98456, 19.98479, 19.98467, 19.98485, 19.9848, 
    19.98476, 19.98478, 19.98469, 19.98467, 19.98458, 19.98462, 19.98436, 
    19.98448, 19.98416, 19.98425, 19.98485, 19.98483, 19.98473, 19.98477, 
    19.98464, 19.98461, 19.98458, 19.98454, 19.98454, 19.98452, 19.98455, 
    19.98452, 19.98464, 19.98459, 19.98474, 19.9847, 19.98472, 19.98474, 
    19.98468, 19.98462, 19.98462, 19.9846, 19.98454, 19.98464, 19.98435, 
    19.98453, 19.98479, 19.98474, 19.98473, 19.98475, 19.98461, 19.98466, 
    19.98452, 19.98456, 19.9845, 19.98453, 19.98453, 19.98457, 19.9846, 
    19.98466, 19.98471, 19.98475, 19.98474, 19.9847, 19.98462, 19.98454, 
    19.98456, 19.9845, 19.98465, 19.98459, 19.98461, 19.98455, 19.98468, 
    19.98457, 19.98471, 19.9847, 19.98466, 19.98458, 19.98457, 19.98455, 
    19.98456, 19.98461, 19.98462, 19.98466, 19.98467, 19.9847, 19.98473, 
    19.98471, 19.98468, 19.98461, 19.98455, 19.98449, 19.98447, 19.98439, 
    19.98445, 19.98435, 19.98444, 19.98428, 19.98456, 19.98444, 19.98466, 
    19.98464, 19.98459, 19.9845, 19.98455, 19.98449, 19.98462, 19.9847, 
    19.98471, 19.98475, 19.98471, 19.98471, 19.98468, 19.98469, 19.98461, 
    19.98466, 19.98453, 19.98449, 19.98436, 19.98428, 19.9842, 19.98417, 
    19.98416, 19.98415,
  19.9861, 19.98604, 19.98605, 19.986, 19.98603, 19.98599, 19.98609, 
    19.98603, 19.98607, 19.9861, 19.9859, 19.98599, 19.98579, 19.98586, 
    19.98569, 19.9858, 19.98567, 19.9857, 19.98562, 19.98565, 19.98555, 
    19.98561, 19.9855, 19.98557, 19.98556, 19.98562, 19.98598, 19.98591, 
    19.98598, 19.98597, 19.98597, 19.98602, 19.98605, 19.98611, 19.9861, 
    19.98606, 19.98596, 19.986, 19.98592, 19.98592, 19.98583, 19.98587, 
    19.98572, 19.98577, 19.98564, 19.98567, 19.98565, 19.98565, 19.98565, 
    19.98569, 19.98567, 19.98571, 19.98586, 19.98582, 19.98595, 19.98603, 
    19.98609, 19.98612, 19.98612, 19.98611, 19.98606, 19.98601, 19.98597, 
    19.98594, 19.98592, 19.98584, 19.9858, 19.98572, 19.98573, 19.9857, 
    19.98568, 19.98563, 19.98564, 19.98562, 19.9857, 19.98565, 19.98574, 
    19.98572, 19.98591, 19.98599, 19.98602, 19.98605, 19.98611, 19.98607, 
    19.98609, 19.98604, 19.98602, 19.98603, 19.98594, 19.98598, 19.9858, 
    19.98588, 19.98568, 19.98573, 19.98567, 19.9857, 19.98565, 19.98569, 
    19.98561, 19.9856, 19.98561, 19.98556, 19.9857, 19.98565, 19.98603, 
    19.98603, 19.98602, 19.98606, 19.98606, 19.98611, 19.98607, 19.98605, 
    19.98601, 19.98599, 19.98597, 19.98592, 19.98586, 19.98578, 19.98573, 
    19.98569, 19.98571, 19.98569, 19.98571, 19.98572, 19.9856, 19.98567, 
    19.98557, 19.98558, 19.98562, 19.98557, 19.98602, 19.98604, 19.98608, 
    19.98605, 19.98611, 19.98608, 19.98606, 19.98598, 19.98596, 19.98594, 
    19.98591, 19.98587, 19.9858, 19.98573, 19.98568, 19.98568, 19.98568, 
    19.98567, 19.9857, 19.98566, 19.98565, 19.98567, 19.98558, 19.9856, 
    19.98558, 19.98559, 19.98603, 19.98601, 19.98602, 19.986, 19.98602, 
    19.98595, 19.98593, 19.98583, 19.98587, 19.98581, 19.98586, 19.98585, 
    19.9858, 19.98586, 19.98574, 19.98582, 19.98567, 19.98575, 19.98566, 
    19.98568, 19.98565, 19.98563, 19.9856, 19.98554, 19.98555, 19.98551, 
    19.98598, 19.98595, 19.98595, 19.98592, 19.9859, 19.98586, 19.98578, 
    19.98581, 19.98575, 19.98574, 19.98582, 19.98577, 19.98593, 19.98591, 
    19.98592, 19.98598, 19.9858, 19.98589, 19.98572, 19.98577, 19.98563, 
    19.9857, 19.98556, 19.9855, 19.98544, 19.98538, 19.98594, 19.98595, 
    19.98592, 19.98587, 19.98583, 19.98577, 19.98576, 19.98575, 19.98572, 
    19.9857, 19.98575, 19.98569, 19.9859, 19.98579, 19.98596, 19.98591, 
    19.98588, 19.98589, 19.98581, 19.98579, 19.98571, 19.98575, 19.98552, 
    19.98562, 19.98533, 19.98541, 19.98596, 19.98594, 19.98585, 19.98589, 
    19.98577, 19.98573, 19.98571, 19.98568, 19.98568, 19.98566, 19.98569, 
    19.98566, 19.98577, 19.98572, 19.98586, 19.98582, 19.98584, 19.98586, 
    19.9858, 19.98575, 19.98575, 19.98573, 19.98568, 19.98577, 19.9855, 
    19.98566, 19.98591, 19.98586, 19.98585, 19.98587, 19.98574, 19.98579, 
    19.98566, 19.98569, 19.98564, 19.98566, 19.98567, 19.9857, 19.98573, 
    19.98578, 19.98583, 19.98587, 19.98586, 19.98582, 19.98574, 19.98568, 
    19.98569, 19.98564, 19.98577, 19.98572, 19.98574, 19.98568, 19.98581, 
    19.9857, 19.98583, 19.98582, 19.98579, 19.98571, 19.9857, 19.98568, 
    19.98569, 19.98574, 19.98575, 19.98579, 19.9858, 19.98583, 19.98585, 
    19.98583, 19.98581, 19.98574, 19.98569, 19.98563, 19.98561, 19.98554, 
    19.9856, 19.9855, 19.98558, 19.98544, 19.9857, 19.98558, 19.98579, 
    19.98576, 19.98573, 19.98564, 19.98568, 19.98563, 19.98575, 19.98582, 
    19.98583, 19.98586, 19.98583, 19.98584, 19.98581, 19.98582, 19.98574, 
    19.98578, 19.98567, 19.98563, 19.98551, 19.98544, 19.98537, 19.98534, 
    19.98533, 19.98532,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222793, 0.7222769, 0.7222774, 0.7222754, 0.7222765, 0.7222753, 
    0.7222788, 0.7222768, 0.7222781, 0.7222791, 0.7222717, 0.7222754, 
    0.7222678, 0.7222702, 0.7222643, 0.7222682, 0.7222635, 0.7222644, 
    0.7222617, 0.7222624, 0.722259, 0.7222613, 0.7222571, 0.7222595, 
    0.7222592, 0.7222614, 0.7222746, 0.7222722, 0.7222748, 0.7222744, 
    0.7222745, 0.7222765, 0.7222775, 0.7222795, 0.7222791, 0.7222776, 
    0.7222742, 0.7222754, 0.7222725, 0.7222726, 0.7222693, 0.7222708, 
    0.7222654, 0.7222669, 0.7222624, 0.7222635, 0.7222624, 0.7222628, 
    0.7222624, 0.7222641, 0.7222634, 0.7222648, 0.7222705, 0.7222688, 
    0.7222738, 0.7222768, 0.7222788, 0.7222801, 0.72228, 0.7222796, 
    0.7222776, 0.7222758, 0.7222744, 0.7222735, 0.7222726, 0.7222698, 
    0.7222683, 0.722265, 0.7222656, 0.7222646, 0.7222636, 0.722262, 
    0.7222623, 0.7222616, 0.7222646, 0.7222626, 0.722266, 0.7222651, 
    0.7222723, 0.7222751, 0.7222763, 0.7222773, 0.7222798, 0.7222781, 
    0.7222788, 0.7222772, 0.7222761, 0.7222766, 0.7222735, 0.7222747, 
    0.7222682, 0.722271, 0.7222638, 0.7222655, 0.7222633, 0.7222645, 
    0.7222626, 0.7222642, 0.7222613, 0.7222607, 0.7222611, 0.7222595, 
    0.7222643, 0.7222624, 0.7222766, 0.7222766, 0.7222762, 0.7222779, 
    0.7222779, 0.7222795, 0.7222781, 0.7222775, 0.722276, 0.7222751, 
    0.7222743, 0.7222725, 0.7222704, 0.7222674, 0.7222654, 0.722264, 
    0.7222648, 0.7222641, 0.7222649, 0.7222653, 0.722261, 0.7222634, 
    0.7222597, 0.7222599, 0.7222615, 0.7222599, 0.7222765, 0.722277, 
    0.7222787, 0.7222773, 0.7222797, 0.7222784, 0.7222776, 0.7222747, 
    0.722274, 0.7222734, 0.7222722, 0.7222707, 0.722268, 0.7222657, 
    0.7222636, 0.7222638, 0.7222637, 0.7222632, 0.7222644, 0.722263, 
    0.7222628, 0.7222634, 0.7222599, 0.7222609, 0.7222599, 0.7222605, 
    0.7222768, 0.722276, 0.7222764, 0.7222756, 0.7222762, 0.7222736, 
    0.7222729, 0.7222692, 0.7222707, 0.7222684, 0.7222705, 0.7222701, 
    0.7222683, 0.7222704, 0.7222658, 0.7222689, 0.7222632, 0.7222663, 
    0.722263, 0.7222636, 0.7222626, 0.7222617, 0.7222607, 0.7222586, 
    0.722259, 0.7222574, 0.7222748, 0.7222738, 0.7222738, 0.7222728, 
    0.7222719, 0.7222702, 0.7222674, 0.7222684, 0.7222665, 0.7222661, 
    0.7222691, 0.7222672, 0.7222731, 0.7222721, 0.7222727, 0.7222747, 
    0.7222682, 0.7222716, 0.7222654, 0.7222672, 0.7222618, 0.7222645, 
    0.7222593, 0.7222571, 0.7222551, 0.7222526, 0.7222732, 0.7222739, 
    0.7222726, 0.7222708, 0.7222692, 0.722267, 0.7222669, 0.7222664, 
    0.7222654, 0.7222645, 0.7222663, 0.7222643, 0.7222719, 0.7222679, 
    0.7222742, 0.7222723, 0.722271, 0.7222716, 0.7222686, 0.7222679, 
    0.722265, 0.7222665, 0.7222577, 0.7222615, 0.7222508, 0.7222537, 
    0.7222741, 0.7222732, 0.7222698, 0.7222714, 0.7222669, 0.7222658, 
    0.7222649, 0.7222638, 0.7222636, 0.7222629, 0.7222641, 0.722263, 
    0.722267, 0.7222652, 0.7222703, 0.722269, 0.7222696, 0.7222702, 
    0.7222683, 0.7222663, 0.7222662, 0.7222656, 0.7222638, 0.7222669, 
    0.7222571, 0.7222632, 0.7222722, 0.7222703, 0.72227, 0.7222707, 
    0.7222659, 0.7222677, 0.7222629, 0.7222642, 0.7222621, 0.7222632, 
    0.7222633, 0.7222646, 0.7222655, 0.7222676, 0.7222693, 0.7222707, 
    0.7222703, 0.7222688, 0.7222661, 0.7222636, 0.7222642, 0.7222623, 
    0.7222672, 0.7222652, 0.722266, 0.7222639, 0.7222685, 0.7222645, 
    0.7222695, 0.7222691, 0.7222677, 0.722265, 0.7222644, 0.7222638, 
    0.7222642, 0.7222661, 0.7222664, 0.7222677, 0.7222681, 0.7222691, 
    0.72227, 0.7222692, 0.7222684, 0.7222661, 0.722264, 0.7222617, 0.7222612, 
    0.7222585, 0.7222607, 0.7222571, 0.7222601, 0.7222549, 0.7222643, 
    0.7222602, 0.7222676, 0.7222669, 0.7222654, 0.7222621, 0.7222639, 
    0.7222618, 0.7222664, 0.7222688, 0.7222694, 0.7222705, 0.7222694, 
    0.7222695, 0.7222683, 0.7222687, 0.722266, 0.7222674, 0.7222633, 
    0.7222618, 0.7222576, 0.7222549, 0.7222522, 0.7222511, 0.7222507, 
    0.7222506 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  -2.006177e-36, 1.541976e-20, 2.055969e-20, -1.027984e-20, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -2.055969e-20, 3.083953e-20, 1.027984e-20, -3.083953e-20, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 2.055969e-20, 2.569961e-20, -1.541976e-20, 
    -1.541976e-20, 1.027984e-20, 0, 3.083953e-20, -1.541976e-20, 
    -4.625929e-20, 1.541976e-20, 2.569961e-20, -1.541976e-20, 1.027984e-20, 
    3.083953e-20, 1.027984e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    -3.597945e-20, 1.541976e-20, -2.055969e-20, 2.055969e-20, 2.055969e-20, 
    2.006177e-36, 1.541976e-20, 1.027984e-20, 4.111937e-20, 5.139921e-21, 
    1.027984e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.541976e-20, 1.541976e-20, 
    -5.139921e-21, 2.006177e-36, -2.006177e-36, 3.083953e-20, -5.139921e-21, 
    -3.083953e-20, 2.055969e-20, -2.055969e-20, -2.569961e-20, 0, 
    -2.569961e-20, 5.139921e-21, 0, -2.055969e-20, -2.569961e-20, 
    -1.027984e-20, 1.541976e-20, -1.027984e-20, -2.006177e-36, -5.139921e-20, 
    2.006177e-36, -1.541976e-20, -1.541976e-20, -1.027984e-20, 4.111937e-20, 
    2.569961e-20, -2.569961e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -2.569961e-20, 1.027984e-20, -1.541976e-20, -1.541976e-20, -5.139921e-21, 
    1.541976e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, 2.055969e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, 1.027984e-20, 2.569961e-20, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, -5.139921e-20, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -5.139921e-21, -2.569961e-20, 0, -5.139921e-21, 
    -3.597945e-20, 1.541976e-20, 1.541976e-20, -2.055969e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, -1.027984e-20, 2.006177e-36, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 
    2.569961e-20, 0, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -2.569961e-20, 1.027984e-20, 
    -5.653913e-20, 4.625929e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, -3.083953e-20, 1.027984e-20, -2.006177e-36, 
    -1.541976e-20, 2.055969e-20, -1.541976e-20, -2.055969e-20, 1.027984e-20, 
    -3.083953e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, -1.541976e-20, 
    1.541976e-20, -2.055969e-20, -2.569961e-20, 5.139921e-21, -5.139921e-21, 
    -2.569961e-20, 1.027984e-20, 3.083953e-20, 3.083953e-20, 5.139921e-21, 
    -2.569961e-20, -2.055969e-20, 0, 1.027984e-20, 2.569961e-20, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, -2.055969e-20, -2.006177e-36, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 0, 0, 1.541976e-20, -5.139921e-21, 0, 
    1.541976e-20, 2.006177e-36, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.055969e-20, -1.027984e-20, 1.027984e-20, -2.055969e-20, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.006177e-36, 1.541976e-20, 2.569961e-20, 
    -2.055969e-20, 5.139921e-21, 1.541976e-20, 3.083953e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -1.541976e-20, 2.569961e-20, -1.027984e-20, 
    5.139921e-21, -2.569961e-20, -1.027984e-20, -1.027984e-20, -2.055969e-20, 
    -1.541976e-20, 2.055969e-20, -1.541976e-20, -2.569961e-20, 1.027984e-20, 
    1.541976e-20, -1.027984e-20, -5.139921e-21, -3.083953e-20, 4.111937e-20, 
    -2.055969e-20, -1.027984e-20, 2.569961e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -3.083953e-20, -2.006177e-36, 2.055969e-20, 
    -1.027984e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, 5.139921e-21, 2.055969e-20, -2.055969e-20, 3.597945e-20, 
    -5.139921e-21, -3.083953e-20, 2.569961e-20, 5.139921e-21, -2.569961e-20, 
    4.111937e-20, 5.139921e-21, 4.111937e-20, -1.541976e-20, -5.139921e-21, 
    3.083953e-20, -1.027984e-20, 5.139921e-21, 2.006177e-36, 2.569961e-20, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, 2.569961e-20, -1.027984e-20, 
    4.625929e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 0, 3.597945e-20, 
    -1.027984e-20, -1.541976e-20, -2.569961e-20, 0, -5.139921e-21, 
    -1.541976e-20, -1.541976e-20, 1.541976e-20, 1.541976e-20, -1.541976e-20, 
    -5.139921e-21, -2.569961e-20, -5.139921e-21, 2.569961e-20, -2.055969e-20, 
    2.569961e-20, 2.055969e-20, -1.027984e-20, 2.055969e-20, -1.541976e-20, 
    2.055969e-20, 2.055969e-20, -1.027984e-20, 2.006177e-36, -2.569961e-20, 
    -3.597945e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, 
    2.569961e-20, -1.541976e-20, 0, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    -3.083953e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    2.055969e-20, -1.027984e-20, -2.569961e-20, -1.027984e-20, -1.027984e-20, 
    -4.625929e-20, 0, -2.055969e-20, -1.541976e-20, -2.569961e-20,
  1.541976e-20, 2.006177e-36, -2.569961e-20, 0, 0, -1.541976e-20, 
    5.139921e-21, 1.027984e-20, -2.006177e-36, 2.006177e-36, -5.139921e-21, 
    -3.083953e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -2.055969e-20, 1.541976e-20, 0, 5.139921e-21, 0, -1.027984e-20, 
    -2.055969e-20, -2.006177e-36, -1.027984e-20, -1.541976e-20, 1.027984e-20, 
    -2.006177e-36, -2.569961e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, 0, 2.569961e-20, 1.027984e-20, -2.569961e-20, 2.569961e-20, 
    3.083953e-20, 2.055969e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 2.055969e-20, 2.569961e-20, 2.055969e-20, 
    -5.139921e-21, 5.139921e-21, 2.569961e-20, -5.139921e-21, 0, 
    1.027984e-20, 0, 1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -4.111937e-20, -2.569961e-20, 1.027984e-20, -2.055969e-20, 
    -5.139921e-21, 2.055969e-20, 5.139921e-21, 5.139921e-21, 0, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    0, 1.541976e-20, 1.541976e-20, 1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -5.139921e-21, 1.541976e-20, 1.027984e-20, -5.139921e-21, -3.083953e-20, 
    -1.027984e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, -1.541976e-20, 
    -1.541976e-20, 0, -1.027984e-20, 0, -5.139921e-21, -2.006177e-36, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 2.055969e-20, 
    3.083953e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -1.027984e-20, 0, -3.083953e-20, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 2.055969e-20, 3.597945e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 1.027984e-20, 0, 5.139921e-21, 
    -1.027984e-20, 1.541976e-20, -5.139921e-21, -2.055969e-20, 0, 
    1.027984e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, 
    5.139921e-21, -2.569961e-20, -1.541976e-20, 2.055969e-20, -1.027984e-20, 
    5.139921e-21, 3.083953e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    0, -5.139921e-21, 1.541976e-20, -1.027984e-20, -2.055969e-20, 
    5.139921e-21, 1.541976e-20, 0, -5.139921e-21, 2.055969e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    2.569961e-20, 1.027984e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, 
    1.541976e-20, 0, -5.139921e-21, -2.055969e-20, 2.055969e-20, 
    -1.541976e-20, 3.083953e-20, -2.006177e-36, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, 2.569961e-20, -2.006177e-36, 
    -1.027984e-20, -3.597945e-20, -2.055969e-20, 0, 1.541976e-20, 
    -2.569961e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, 5.139921e-21, -2.006177e-36, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, 2.569961e-20, 3.597945e-20, 1.027984e-20, -1.027984e-20, 
    3.083953e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -2.006177e-36, -2.055969e-20, -5.139921e-21, -1.541976e-20, 2.055969e-20, 
    2.055969e-20, -1.541976e-20, -1.541976e-20, 2.569961e-20, -3.597945e-20, 
    0, 5.139921e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -1.541976e-20, 0, -2.569961e-20, 
    -1.541976e-20, -1.541976e-20, -5.139921e-21, -2.055969e-20, 5.139921e-21, 
    2.055969e-20, 5.139921e-21, 5.139921e-21, -1.541976e-20, 5.139921e-21, 0, 
    -1.027984e-20, -2.055969e-20, 5.139921e-21, 5.139921e-21, -2.006177e-36, 
    -1.027984e-20, -2.055969e-20, 1.541976e-20, 1.027984e-20, -3.083953e-20, 
    -1.541976e-20, 2.569961e-20, 3.083953e-20, 1.027984e-20, -2.006177e-36, 
    1.541976e-20, 1.541976e-20, 0, 0, -2.055969e-20, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, -2.006177e-36, 2.569961e-20, 2.006177e-36, 
    -1.541976e-20, 0, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, 0, 0, -2.055969e-20, -2.055969e-20, -2.055969e-20, 
    1.541976e-20, 0, -2.055969e-20, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, 5.139921e-21, -2.055969e-20, 2.006177e-36, -5.139921e-21, 
    2.569961e-20, -2.569961e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 
    -2.006177e-36, 0, -3.083953e-20, -1.027984e-20, 2.569961e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, 2.569961e-20, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, 0, 2.055969e-20,
  1.027984e-20, -3.083953e-20, -5.139921e-21, -1.541976e-20, 1.541976e-20, 
    2.055969e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 3.083953e-20, -1.541976e-20, 2.055969e-20, 3.083953e-20, 
    5.139921e-21, -3.597945e-20, 5.139921e-21, 5.139921e-21, 2.006177e-36, 
    -1.027984e-20, -4.111937e-20, 1.541976e-20, 2.006177e-36, 5.139921e-21, 
    -2.006177e-36, 5.139921e-21, -1.541976e-20, -1.027984e-20, 0, 
    1.027984e-20, -2.006177e-36, -5.139921e-21, 1.541976e-20, 0, 
    -5.139921e-21, -1.541976e-20, 3.083953e-20, -5.139921e-21, 1.027984e-20, 
    -2.055969e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -4.111937e-20, 3.083953e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, -2.055969e-20, 2.055969e-20, -2.055969e-20, 
    -5.139921e-21, 5.653913e-20, -5.139921e-21, -2.055969e-20, 1.027984e-20, 
    1.027984e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 2.055969e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -2.569961e-20, -2.055969e-20, 3.083953e-20, -2.569961e-20, -2.055969e-20, 
    -1.541976e-20, 1.541976e-20, -1.541976e-20, -1.541976e-20, -2.569961e-20, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, -2.569961e-20, 
    0, 5.139921e-21, -5.139921e-21, 2.055969e-20, 5.139921e-21, 5.139921e-21, 
    1.541976e-20, -3.083953e-20, 2.569961e-20, 5.139921e-21, 1.541976e-20, 0, 
    5.139921e-21, -5.139921e-21, -2.006177e-36, -2.055969e-20, 0, 
    -2.006177e-36, 2.055969e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, 2.055969e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, -3.597945e-20, -1.541976e-20, 1.541976e-20, 2.055969e-20, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, 
    -2.006177e-36, -2.569961e-20, -5.139921e-21, -2.055969e-20, 
    -2.055969e-20, 2.055969e-20, -5.139921e-21, -2.006177e-36, 1.541976e-20, 
    1.027984e-20, -1.027984e-20, 3.083953e-20, 4.111937e-20, 3.083953e-20, 
    1.027984e-20, 5.139921e-21, 4.625929e-20, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    4.111937e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, -2.055969e-20, -3.083953e-20, 
    -1.541976e-20, 3.083953e-20, -1.541976e-20, 2.055969e-20, 2.055969e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -2.006177e-36, 2.006177e-36, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 2.055969e-20, 
    -1.027984e-20, -2.006177e-36, -1.027984e-20, 3.083953e-20, -1.027984e-20, 
    -2.055969e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, -5.653913e-20, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, -2.055969e-20, 
    -1.541976e-20, 2.569961e-20, -5.139921e-21, 2.055969e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, -4.111937e-20, 2.006177e-36, -4.111937e-20, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 2.569961e-20, 1.541976e-20, 
    -5.139921e-21, 0, -2.006177e-36, -5.139921e-21, 2.569961e-20, 
    1.027984e-20, -5.139921e-21, 2.055969e-20, -2.055969e-20, 2.055969e-20, 
    3.597945e-20, -5.139921e-21, -2.055969e-20, 1.027984e-20, 1.027984e-20, 
    -2.055969e-20, 1.541976e-20, -2.006177e-36, 5.139921e-21, 2.006177e-36, 
    1.027984e-20, 1.027984e-20, 0, 1.027984e-20, -2.006177e-36, 5.139921e-21, 
    2.006177e-36, 3.083953e-20, 3.083953e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-20, -5.139921e-21, 5.139921e-21, 4.625929e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 0, -2.569961e-20, 2.055969e-20, 
    5.139921e-21, -2.055969e-20, 3.597945e-20, -2.006177e-36, 2.569961e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, -2.006177e-36, 4.111937e-20, 
    1.541976e-20, -1.027984e-20, -2.006177e-36, 2.055969e-20, 3.083953e-20, 
    -1.027984e-20, -2.055969e-20, -2.055969e-20, -1.541976e-20, 1.027984e-20, 
    2.006177e-36, -5.139921e-21, -2.006177e-36, -2.006177e-36, 1.541976e-20, 
    -2.569961e-20, -5.139921e-21, 1.027984e-20, 0, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 2.055969e-20, -2.006177e-36, 5.139921e-21, 
    -2.569961e-20, 5.139921e-21, -2.569961e-20, -5.139921e-21, -2.006177e-36, 
    -2.055969e-20, 2.569961e-20, -2.055969e-20, 5.139921e-21, -2.055969e-20, 
    2.006177e-36, 4.625929e-20, -5.139921e-21, 1.541976e-20, 3.083953e-20, 
    -2.569961e-20, -2.055969e-20, -1.541976e-20, 1.027984e-20, 0, 
    2.569961e-20, 1.541976e-20, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    3.597945e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, 1.027984e-20, 
    2.569961e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, -2.006177e-36, 
    5.139921e-21,
  -2.006177e-36, 2.569961e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 2.055969e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -1.541976e-20, -3.083953e-20, 2.055969e-20, 2.569961e-20, -2.569961e-20, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    1.027984e-20, 0, 0, 2.055969e-20, 5.139921e-21, 2.055969e-20, 
    -1.027984e-20, -5.139921e-21, 1.541976e-20, 2.055969e-20, 5.139921e-21, 
    2.569961e-20, -3.597945e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -2.006177e-36, 2.569961e-20, -1.027984e-20, 1.027984e-20, -3.083953e-20, 
    -2.569961e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -3.597945e-20, 3.597945e-20, 1.027984e-20, 2.006177e-36, 2.055969e-20, 
    -1.541976e-20, 2.055969e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, -1.027984e-20, -2.055969e-20, 3.083953e-20, 4.111937e-20, 
    3.083953e-20, 5.139921e-21, 2.006177e-36, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, -3.597945e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, -2.055969e-20, -2.569961e-20, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, 2.055969e-20, -1.541976e-20, 
    -1.541976e-20, 4.625929e-20, -1.541976e-20, 1.541976e-20, 2.055969e-20, 
    -1.027984e-20, 0, 1.541976e-20, -1.541976e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, -1.027984e-20, -1.541976e-20, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, 2.055969e-20, 2.569961e-20, 2.569961e-20, 
    2.055969e-20, -3.597945e-20, 5.139921e-21, 2.569961e-20, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 2.006177e-36, 2.055969e-20, 
    -1.027984e-20, 0, 3.083953e-20, -1.027984e-20, 2.055969e-20, 
    2.055969e-20, -1.541976e-20, -1.541976e-20, -2.569961e-20, 0, 
    1.027984e-20, 5.139921e-21, -3.083953e-20, 2.006177e-36, -5.139921e-21, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    5.139921e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, -2.006177e-36, 
    -2.006177e-36, 5.139921e-21, 1.027984e-20, 5.139921e-21, 3.083953e-20, 
    -3.597945e-20, -1.027984e-20, -2.055969e-20, 2.055969e-20, 1.541976e-20, 
    -2.006177e-36, 2.055969e-20, -2.055969e-20, 5.139921e-21, -3.597945e-20, 
    -1.541976e-20, -2.569961e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 3.597945e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    0, -1.541976e-20, 2.569961e-20, -3.597945e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -4.625929e-20, 1.027984e-20, -1.027984e-20, 
    0, -1.541976e-20, 5.139921e-21, -3.597945e-20, 1.027984e-20, 
    1.027984e-20, 4.111937e-20, 3.083953e-20, -2.055969e-20, 3.083953e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, -3.083953e-20, -4.111937e-20, 
    -5.139921e-21, -5.139921e-21, 2.055969e-20, 2.569961e-20, -2.006177e-36, 
    -5.139921e-21, 2.055969e-20, -3.083953e-20, -1.027984e-20, 1.541976e-20, 
    1.027984e-20, 2.569961e-20, -1.027984e-20, 3.597945e-20, -1.541976e-20, 
    2.569961e-20, 5.139921e-21, 2.006177e-36, -3.083953e-20, 0, 
    -1.027984e-20, 0, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -3.597945e-20, -3.083953e-20, 1.541976e-20, 2.055969e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, -1.541976e-20, 2.055969e-20, 
    -2.055969e-20, -5.139921e-21, 4.111937e-20, 0, -1.541976e-20, 0, 
    -2.055969e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, -2.006177e-36, 
    2.569961e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, -1.541976e-20, 
    -2.055969e-20, -1.541976e-20, -2.569961e-20, 0, -1.541976e-20, 
    1.541976e-20, 1.027984e-20, 0, 5.139921e-21, 1.027984e-20, 0, 
    -1.541976e-20, 0, -1.027984e-20, -2.055969e-20, -1.027984e-20, 
    2.569961e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, -5.653913e-20, 
    -5.139921e-21, 2.006177e-36, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -4.111937e-20, -1.027984e-20, -5.139921e-21, 2.006177e-36, -4.111937e-20, 
    -2.569961e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -2.055969e-20, -2.055969e-20, 1.027984e-20, -4.111937e-20, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, 3.083953e-20, 3.083953e-20, 
    -1.541976e-20, -1.541976e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    -3.597945e-20, -5.139921e-21, 2.055969e-20, -1.027984e-20, -5.139921e-21, 
    2.055969e-20, -4.625929e-20, 1.541976e-20, 1.027984e-20, -3.083953e-20, 
    -1.541976e-20, -1.541976e-20, -1.541976e-20, -2.006177e-36, 
    -2.006177e-36, 5.139921e-21, 2.055969e-20, 5.139921e-21, 2.569961e-20, 
    -2.569961e-20, 0, 2.006177e-36, 1.027984e-20, -2.055969e-20, 
    -2.055969e-20, -2.569961e-20, 0, -1.541976e-20, -5.139921e-21, 
    2.006177e-36, -1.027984e-20, 1.541976e-20, -2.569961e-20, 1.027984e-20, 
    1.541976e-20, -1.027984e-20, -1.541976e-20, -1.541976e-20, 5.139921e-21, 
    2.055969e-20, -1.541976e-20, -3.597945e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21,
  -3.083953e-20, -1.541976e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    0, 2.006177e-36, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, 2.006177e-36, 5.139921e-21, 3.597945e-20, 2.569961e-20, 
    1.541976e-20, 5.139921e-21, 2.055969e-20, 2.055969e-20, -3.597945e-20, 
    -1.541976e-20, -2.055969e-20, 2.055969e-20, -4.625929e-20, 1.027984e-20, 
    1.541976e-20, 2.006177e-36, 1.541976e-20, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, -1.541976e-20, -1.541976e-20, 2.055969e-20, 2.055969e-20, 
    -5.139921e-21, 2.569961e-20, -3.083953e-20, -2.569961e-20, -1.541976e-20, 
    -4.111937e-20, -1.541976e-20, -3.083953e-20, -2.569961e-20, 
    -1.027984e-20, 1.541976e-20, -2.055969e-20, 0, 2.569961e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -1.541976e-20, 2.055969e-20, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, -2.006177e-36, 
    -1.541976e-20, 1.027984e-20, -1.541976e-20, -1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 0, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, -2.055969e-20, -5.139921e-21, 1.541976e-20, -2.569961e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 2.569961e-20, 3.083953e-20, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, -2.055969e-20, 
    -2.006177e-36, 5.139921e-21, 1.541976e-20, 1.541976e-20, -2.569961e-20, 
    1.027984e-20, 5.139921e-21, -2.055969e-20, -4.111937e-20, -2.055969e-20, 
    1.027984e-20, -2.006177e-36, -2.569961e-20, 0, 0, -1.541976e-20, 
    2.055969e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 0, 5.139921e-21, 
    2.006177e-36, 5.139921e-21, -5.139921e-21, 3.597945e-20, 1.027984e-20, 
    -5.139921e-21, 2.055969e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    2.006177e-36, -2.055969e-20, 2.055969e-20, -1.027984e-20, -1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 2.006177e-36, 1.027984e-20, 0, 
    2.055969e-20, -1.027984e-20, 1.027984e-20, -2.055969e-20, -1.541976e-20, 
    2.055969e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, -2.055969e-20, 
    1.541976e-20, 1.541976e-20, -5.139921e-21, 3.083953e-20, -2.569961e-20, 
    5.139921e-21, -2.055969e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    0, 5.139921e-21, 0, -2.569961e-20, 2.055969e-20, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, -2.055969e-20, 2.055969e-20, 2.055969e-20, 
    -3.083953e-20, -1.027984e-20, 2.055969e-20, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.006177e-36, -2.055969e-20, -2.569961e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-20, 2.569961e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, 1.027984e-20, 3.597945e-20, 
    -1.027984e-20, -2.055969e-20, 0, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, -1.541976e-20, 3.597945e-20, 5.139921e-21, 2.055969e-20, 
    0, 1.027984e-20, 1.541976e-20, 0, -2.006177e-36, 1.027984e-20, 
    -1.541976e-20, 2.055969e-20, -1.541976e-20, -3.597945e-20, 1.541976e-20, 
    1.541976e-20, 0, 0, 2.055969e-20, 5.139921e-21, 0, -1.541976e-20, 
    -4.111937e-20, -1.541976e-20, -4.625929e-20, 5.139921e-21, 5.139921e-21, 
    0, 2.569961e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -2.006177e-36, 3.597945e-20, -2.569961e-20, 1.027984e-20, 2.055969e-20, 
    0, -2.569961e-20, -1.541976e-20, -1.541976e-20, 2.055969e-20, 
    -1.541976e-20, 1.541976e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 
    -1.027984e-20, -1.541976e-20, -2.055969e-20, 1.541976e-20, 0, 
    2.055969e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.055969e-20, -1.541976e-20, 
    -2.569961e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, -2.006177e-36, 
    2.569961e-20, -3.083953e-20, 2.569961e-20, 3.083953e-20, 1.027984e-20, 
    5.139921e-21, -2.569961e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 2.569961e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    2.006177e-36, 1.027984e-20, -5.139921e-21, 2.569961e-20, 2.055969e-20, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    -2.055969e-20, 4.111937e-20, -2.055969e-20, 0, -5.139921e-21, 
    -5.139921e-21, 3.597945e-20, 1.541976e-20, 2.055969e-20, -3.083953e-20, 
    -1.027984e-20, -2.055969e-20, 0, -1.027984e-20, -2.006177e-36, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -5.139921e-21, 3.083953e-20, -5.139921e-21, -3.597945e-20, 2.055969e-20, 
    0, -1.027984e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, -4.111937e-20, 2.055969e-20, 
    -5.139921e-21, 2.055969e-20, -5.139921e-21, -2.006177e-36, 1.027984e-20, 
    -3.083953e-20, -2.006177e-36, 0, -3.083953e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 2.569961e-20, 5.139921e-21,
  8.598834e-29, 8.598806e-29, 8.598811e-29, 8.598789e-29, 8.598802e-29, 
    8.598787e-29, 8.598828e-29, 8.598805e-29, 8.59882e-29, 8.598832e-29, 
    8.598745e-29, 8.598788e-29, 8.598701e-29, 8.598728e-29, 8.598659e-29, 
    8.598705e-29, 8.598649e-29, 8.59866e-29, 8.598628e-29, 8.598637e-29, 
    8.598597e-29, 8.598624e-29, 8.598576e-29, 8.598604e-29, 8.598599e-29, 
    8.598625e-29, 8.598779e-29, 8.598751e-29, 8.598781e-29, 8.598777e-29, 
    8.598779e-29, 8.598801e-29, 8.598813e-29, 8.598836e-29, 8.598832e-29, 
    8.598814e-29, 8.598775e-29, 8.598788e-29, 8.598755e-29, 8.598755e-29, 
    8.598717e-29, 8.598735e-29, 8.598671e-29, 8.598689e-29, 8.598637e-29, 
    8.59865e-29, 8.598638e-29, 8.598642e-29, 8.598638e-29, 8.598657e-29, 
    8.598649e-29, 8.598666e-29, 8.598731e-29, 8.598712e-29, 8.59877e-29, 
    8.598805e-29, 8.598828e-29, 8.598844e-29, 8.598841e-29, 8.598837e-29, 
    8.598814e-29, 8.598793e-29, 8.598777e-29, 8.598766e-29, 8.598755e-29, 
    8.598723e-29, 8.598706e-29, 8.598668e-29, 8.598675e-29, 8.598663e-29, 
    8.598652e-29, 8.598633e-29, 8.598636e-29, 8.598628e-29, 8.598663e-29, 
    8.59864e-29, 8.598678e-29, 8.598668e-29, 8.598752e-29, 8.598785e-29, 
    8.598799e-29, 8.598811e-29, 8.59884e-29, 8.59882e-29, 8.598828e-29, 
    8.598808e-29, 8.598796e-29, 8.598802e-29, 8.598766e-29, 8.59878e-29, 
    8.598705e-29, 8.598737e-29, 8.598653e-29, 8.598673e-29, 8.598648e-29, 
    8.598661e-29, 8.598639e-29, 8.598658e-29, 8.598625e-29, 8.598617e-29, 
    8.598622e-29, 8.598603e-29, 8.59866e-29, 8.598638e-29, 8.598803e-29, 
    8.598802e-29, 8.598797e-29, 8.598817e-29, 8.598818e-29, 8.598837e-29, 
    8.59882e-29, 8.598813e-29, 8.598796e-29, 8.598785e-29, 8.598776e-29, 
    8.598754e-29, 8.59873e-29, 8.598696e-29, 8.598672e-29, 8.598655e-29, 
    8.598666e-29, 8.598657e-29, 8.598666e-29, 8.598671e-29, 8.59862e-29, 
    8.598649e-29, 8.598606e-29, 8.598608e-29, 8.598627e-29, 8.598607e-29, 
    8.598801e-29, 8.598807e-29, 8.598826e-29, 8.598811e-29, 8.598838e-29, 
    8.598823e-29, 8.598814e-29, 8.59878e-29, 8.598772e-29, 8.598766e-29, 
    8.598752e-29, 8.598734e-29, 8.598703e-29, 8.598676e-29, 8.598651e-29, 
    8.598653e-29, 8.598652e-29, 8.598646e-29, 8.59866e-29, 8.598645e-29, 
    8.598642e-29, 8.598649e-29, 8.598608e-29, 8.59862e-29, 8.598608e-29, 
    8.598615e-29, 8.598805e-29, 8.598796e-29, 8.598801e-29, 8.598791e-29, 
    8.598798e-29, 8.598768e-29, 8.598759e-29, 8.598717e-29, 8.598734e-29, 
    8.598707e-29, 8.598731e-29, 8.598727e-29, 8.598706e-29, 8.59873e-29, 
    8.598677e-29, 8.598713e-29, 8.598646e-29, 8.598683e-29, 8.598644e-29, 
    8.598651e-29, 8.59864e-29, 8.59863e-29, 8.598616e-29, 8.598593e-29, 
    8.598598e-29, 8.598578e-29, 8.598781e-29, 8.598769e-29, 8.59877e-29, 
    8.598758e-29, 8.598748e-29, 8.598728e-29, 8.598695e-29, 8.598707e-29, 
    8.598685e-29, 8.59868e-29, 8.598714e-29, 8.598693e-29, 8.598761e-29, 
    8.59875e-29, 8.598757e-29, 8.598781e-29, 8.598704e-29, 8.598743e-29, 
    8.598672e-29, 8.598693e-29, 8.598631e-29, 8.598662e-29, 8.598601e-29, 
    8.598575e-29, 8.598551e-29, 8.598522e-29, 8.598763e-29, 8.598771e-29, 
    8.598756e-29, 8.598736e-29, 8.598717e-29, 8.598692e-29, 8.598689e-29, 
    8.598684e-29, 8.598672e-29, 8.598662e-29, 8.598683e-29, 8.598659e-29, 
    8.598748e-29, 8.598701e-29, 8.598774e-29, 8.598752e-29, 8.598737e-29, 
    8.598743e-29, 8.598709e-29, 8.598701e-29, 8.598668e-29, 8.598684e-29, 
    8.598581e-29, 8.598627e-29, 8.598501e-29, 8.598536e-29, 8.598774e-29, 
    8.598763e-29, 8.598724e-29, 8.598742e-29, 8.59869e-29, 8.598677e-29, 
    8.598666e-29, 8.598652e-29, 8.598651e-29, 8.598643e-29, 8.598656e-29, 
    8.598643e-29, 8.598691e-29, 8.59867e-29, 8.598728e-29, 8.598714e-29, 
    8.59872e-29, 8.598728e-29, 8.598706e-29, 8.598682e-29, 8.598682e-29, 
    8.598674e-29, 8.598652e-29, 8.598689e-29, 8.598576e-29, 8.598646e-29, 
    8.598751e-29, 8.598729e-29, 8.598726e-29, 8.598734e-29, 8.598678e-29, 
    8.598698e-29, 8.598643e-29, 8.598658e-29, 8.598634e-29, 8.598646e-29, 
    8.598648e-29, 8.598663e-29, 8.598673e-29, 8.598698e-29, 8.598717e-29, 
    8.598733e-29, 8.59873e-29, 8.598712e-29, 8.598681e-29, 8.598651e-29, 
    8.598657e-29, 8.598636e-29, 8.598693e-29, 8.598669e-29, 8.598678e-29, 
    8.598654e-29, 8.598708e-29, 8.598662e-29, 8.598719e-29, 8.598714e-29, 
    8.598699e-29, 8.598668e-29, 8.598661e-29, 8.598653e-29, 8.598658e-29, 
    8.59868e-29, 8.598684e-29, 8.598699e-29, 8.598704e-29, 8.598716e-29, 
    8.598725e-29, 8.598716e-29, 8.598707e-29, 8.59868e-29, 8.598655e-29, 
    8.598629e-29, 8.598623e-29, 8.598592e-29, 8.598617e-29, 8.598575e-29, 
    8.598611e-29, 8.59855e-29, 8.59866e-29, 8.598612e-29, 8.598698e-29, 
    8.598689e-29, 8.598672e-29, 8.598633e-29, 8.598654e-29, 8.59863e-29, 
    8.598684e-29, 8.598711e-29, 8.598719e-29, 8.598732e-29, 8.598719e-29, 
    8.598719e-29, 8.598707e-29, 8.598711e-29, 8.598679e-29, 8.598696e-29, 
    8.598648e-29, 8.59863e-29, 8.59858e-29, 8.59855e-29, 8.598518e-29, 
    8.598505e-29, 8.598501e-29, 8.598499e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.135031e-08, 1.14007e-08, 1.139091e-08, 1.143155e-08, 1.1409e-08, 
    1.143562e-08, 1.136053e-08, 1.14027e-08, 1.137578e-08, 1.135485e-08, 
    1.151043e-08, 1.143336e-08, 1.159052e-08, 1.154135e-08, 1.166487e-08, 
    1.158287e-08, 1.168141e-08, 1.166251e-08, 1.171941e-08, 1.170311e-08, 
    1.177589e-08, 1.172693e-08, 1.181362e-08, 1.17642e-08, 1.177193e-08, 
    1.172532e-08, 1.144888e-08, 1.150084e-08, 1.14458e-08, 1.145321e-08, 
    1.144988e-08, 1.140947e-08, 1.13891e-08, 1.134646e-08, 1.13542e-08, 
    1.138552e-08, 1.145654e-08, 1.143243e-08, 1.149319e-08, 1.149182e-08, 
    1.155947e-08, 1.152897e-08, 1.164269e-08, 1.161037e-08, 1.170379e-08, 
    1.168029e-08, 1.170269e-08, 1.16959e-08, 1.170277e-08, 1.166831e-08, 
    1.168308e-08, 1.165276e-08, 1.153468e-08, 1.156938e-08, 1.14659e-08, 
    1.140369e-08, 1.136238e-08, 1.133306e-08, 1.133721e-08, 1.134511e-08, 
    1.138571e-08, 1.142388e-08, 1.145298e-08, 1.147244e-08, 1.149162e-08, 
    1.154967e-08, 1.158041e-08, 1.164923e-08, 1.163681e-08, 1.165785e-08, 
    1.167796e-08, 1.171171e-08, 1.170615e-08, 1.172102e-08, 1.16573e-08, 
    1.169965e-08, 1.162974e-08, 1.164886e-08, 1.149683e-08, 1.143894e-08, 
    1.141432e-08, 1.139279e-08, 1.134039e-08, 1.137657e-08, 1.136231e-08, 
    1.139625e-08, 1.141781e-08, 1.140715e-08, 1.147298e-08, 1.144738e-08, 
    1.158223e-08, 1.152414e-08, 1.167561e-08, 1.163936e-08, 1.16843e-08, 
    1.166137e-08, 1.170066e-08, 1.16653e-08, 1.172656e-08, 1.17399e-08, 
    1.173078e-08, 1.17658e-08, 1.166334e-08, 1.170268e-08, 1.140685e-08, 
    1.140859e-08, 1.141669e-08, 1.138107e-08, 1.137889e-08, 1.134625e-08, 
    1.137529e-08, 1.138766e-08, 1.141906e-08, 1.143764e-08, 1.145529e-08, 
    1.149412e-08, 1.153748e-08, 1.159813e-08, 1.164171e-08, 1.167092e-08, 
    1.165301e-08, 1.166883e-08, 1.165115e-08, 1.164286e-08, 1.17349e-08, 
    1.168322e-08, 1.176077e-08, 1.175647e-08, 1.172138e-08, 1.175696e-08, 
    1.140981e-08, 1.13998e-08, 1.136505e-08, 1.139224e-08, 1.134269e-08, 
    1.137043e-08, 1.138637e-08, 1.144791e-08, 1.146144e-08, 1.147398e-08, 
    1.149874e-08, 1.153053e-08, 1.158629e-08, 1.163482e-08, 1.167913e-08, 
    1.167588e-08, 1.167702e-08, 1.168692e-08, 1.16624e-08, 1.169094e-08, 
    1.169573e-08, 1.168321e-08, 1.17559e-08, 1.173513e-08, 1.175638e-08, 
    1.174286e-08, 1.140305e-08, 1.14199e-08, 1.141079e-08, 1.142791e-08, 
    1.141585e-08, 1.146947e-08, 1.148554e-08, 1.156078e-08, 1.15299e-08, 
    1.157905e-08, 1.15349e-08, 1.154272e-08, 1.158065e-08, 1.153728e-08, 
    1.163214e-08, 1.156782e-08, 1.16873e-08, 1.162306e-08, 1.169133e-08, 
    1.167893e-08, 1.169946e-08, 1.171784e-08, 1.174097e-08, 1.178364e-08, 
    1.177376e-08, 1.180945e-08, 1.144501e-08, 1.146685e-08, 1.146493e-08, 
    1.14878e-08, 1.150471e-08, 1.154137e-08, 1.160016e-08, 1.157805e-08, 
    1.161865e-08, 1.16268e-08, 1.156512e-08, 1.160299e-08, 1.148148e-08, 
    1.15011e-08, 1.148942e-08, 1.144673e-08, 1.158315e-08, 1.151313e-08, 
    1.164243e-08, 1.160449e-08, 1.171522e-08, 1.166015e-08, 1.176832e-08, 
    1.181457e-08, 1.185811e-08, 1.190898e-08, 1.147878e-08, 1.146393e-08, 
    1.149052e-08, 1.15273e-08, 1.156143e-08, 1.160681e-08, 1.161145e-08, 
    1.161995e-08, 1.164198e-08, 1.166049e-08, 1.162264e-08, 1.166514e-08, 
    1.150565e-08, 1.158922e-08, 1.145832e-08, 1.149773e-08, 1.152513e-08, 
    1.151311e-08, 1.157553e-08, 1.159024e-08, 1.165002e-08, 1.161912e-08, 
    1.180315e-08, 1.172172e-08, 1.194773e-08, 1.188456e-08, 1.145875e-08, 
    1.147873e-08, 1.154828e-08, 1.151519e-08, 1.160984e-08, 1.163314e-08, 
    1.165208e-08, 1.16763e-08, 1.167891e-08, 1.169326e-08, 1.166975e-08, 
    1.169233e-08, 1.16069e-08, 1.164508e-08, 1.154033e-08, 1.156582e-08, 
    1.15541e-08, 1.154123e-08, 1.158094e-08, 1.162323e-08, 1.162414e-08, 
    1.163771e-08, 1.167593e-08, 1.161022e-08, 1.181366e-08, 1.168801e-08, 
    1.150052e-08, 1.153901e-08, 1.154451e-08, 1.15296e-08, 1.16308e-08, 
    1.159413e-08, 1.169291e-08, 1.166621e-08, 1.170996e-08, 1.168822e-08, 
    1.168502e-08, 1.16571e-08, 1.163972e-08, 1.159581e-08, 1.156009e-08, 
    1.153176e-08, 1.153835e-08, 1.156946e-08, 1.162582e-08, 1.167915e-08, 
    1.166747e-08, 1.170663e-08, 1.160297e-08, 1.164644e-08, 1.162964e-08, 
    1.167344e-08, 1.157747e-08, 1.165919e-08, 1.155658e-08, 1.156557e-08, 
    1.15934e-08, 1.164938e-08, 1.166177e-08, 1.1675e-08, 1.166684e-08, 
    1.162725e-08, 1.162077e-08, 1.159273e-08, 1.158498e-08, 1.156362e-08, 
    1.154593e-08, 1.156209e-08, 1.157906e-08, 1.162727e-08, 1.167072e-08, 
    1.17181e-08, 1.17297e-08, 1.178505e-08, 1.173999e-08, 1.181436e-08, 
    1.175112e-08, 1.186059e-08, 1.166393e-08, 1.174927e-08, 1.159467e-08, 
    1.161132e-08, 1.164144e-08, 1.171054e-08, 1.167324e-08, 1.171686e-08, 
    1.162052e-08, 1.157054e-08, 1.155761e-08, 1.153348e-08, 1.155816e-08, 
    1.155615e-08, 1.157977e-08, 1.157218e-08, 1.162887e-08, 1.159842e-08, 
    1.168494e-08, 1.171652e-08, 1.180571e-08, 1.18604e-08, 1.191607e-08, 
    1.194066e-08, 1.194814e-08, 1.195127e-08 ;

 SOIL1N_TO_SOIL3N =
  1.34673e-10, 1.352711e-10, 1.351548e-10, 1.356372e-10, 1.353696e-10, 
    1.356855e-10, 1.347942e-10, 1.352948e-10, 1.349753e-10, 1.347268e-10, 
    1.365736e-10, 1.356588e-10, 1.375242e-10, 1.369406e-10, 1.384068e-10, 
    1.374334e-10, 1.386031e-10, 1.383788e-10, 1.390542e-10, 1.388607e-10, 
    1.397246e-10, 1.391435e-10, 1.401725e-10, 1.395858e-10, 1.396776e-10, 
    1.391243e-10, 1.358429e-10, 1.364597e-10, 1.358063e-10, 1.358943e-10, 
    1.358548e-10, 1.353751e-10, 1.351334e-10, 1.346273e-10, 1.347192e-10, 
    1.350909e-10, 1.359338e-10, 1.356477e-10, 1.363689e-10, 1.363526e-10, 
    1.371557e-10, 1.367936e-10, 1.381435e-10, 1.377598e-10, 1.388687e-10, 
    1.385898e-10, 1.388556e-10, 1.38775e-10, 1.388567e-10, 1.384476e-10, 
    1.386229e-10, 1.38263e-10, 1.368614e-10, 1.372732e-10, 1.36045e-10, 
    1.353065e-10, 1.348162e-10, 1.344682e-10, 1.345174e-10, 1.346112e-10, 
    1.350931e-10, 1.355463e-10, 1.358916e-10, 1.361226e-10, 1.363503e-10, 
    1.370394e-10, 1.374042e-10, 1.382211e-10, 1.380737e-10, 1.383234e-10, 
    1.385621e-10, 1.389627e-10, 1.388968e-10, 1.390733e-10, 1.383169e-10, 
    1.388196e-10, 1.379897e-10, 1.382167e-10, 1.364121e-10, 1.357249e-10, 
    1.354328e-10, 1.351771e-10, 1.345552e-10, 1.349847e-10, 1.348154e-10, 
    1.352182e-10, 1.354742e-10, 1.353476e-10, 1.36129e-10, 1.358252e-10, 
    1.374258e-10, 1.367363e-10, 1.385342e-10, 1.38104e-10, 1.386374e-10, 
    1.383652e-10, 1.388316e-10, 1.384118e-10, 1.39139e-10, 1.392974e-10, 
    1.391891e-10, 1.396049e-10, 1.383886e-10, 1.388556e-10, 1.35344e-10, 
    1.353647e-10, 1.354609e-10, 1.35038e-10, 1.350122e-10, 1.346248e-10, 
    1.349695e-10, 1.351163e-10, 1.35489e-10, 1.357095e-10, 1.359191e-10, 
    1.363799e-10, 1.368947e-10, 1.376146e-10, 1.381318e-10, 1.384786e-10, 
    1.38266e-10, 1.384537e-10, 1.382438e-10, 1.381455e-10, 1.39238e-10, 
    1.386245e-10, 1.395451e-10, 1.394941e-10, 1.390775e-10, 1.394999e-10, 
    1.353792e-10, 1.352604e-10, 1.348479e-10, 1.351707e-10, 1.345826e-10, 
    1.349117e-10, 1.35101e-10, 1.358315e-10, 1.35992e-10, 1.361408e-10, 
    1.364348e-10, 1.368121e-10, 1.37474e-10, 1.3805e-10, 1.38576e-10, 
    1.385374e-10, 1.38551e-10, 1.386685e-10, 1.383775e-10, 1.387163e-10, 
    1.387731e-10, 1.386245e-10, 1.394873e-10, 1.392408e-10, 1.394931e-10, 
    1.393325e-10, 1.35299e-10, 1.354989e-10, 1.353909e-10, 1.35594e-10, 
    1.354509e-10, 1.360873e-10, 1.362781e-10, 1.371712e-10, 1.368047e-10, 
    1.37388e-10, 1.368639e-10, 1.369568e-10, 1.37407e-10, 1.368923e-10, 
    1.380183e-10, 1.372548e-10, 1.38673e-10, 1.379105e-10, 1.387208e-10, 
    1.385737e-10, 1.388173e-10, 1.390355e-10, 1.393101e-10, 1.398166e-10, 
    1.396993e-10, 1.40123e-10, 1.35797e-10, 1.360563e-10, 1.360335e-10, 
    1.363049e-10, 1.365056e-10, 1.369407e-10, 1.376387e-10, 1.373762e-10, 
    1.378581e-10, 1.379548e-10, 1.372228e-10, 1.376722e-10, 1.362299e-10, 
    1.364629e-10, 1.363241e-10, 1.358174e-10, 1.374367e-10, 1.366056e-10, 
    1.381404e-10, 1.376901e-10, 1.390044e-10, 1.383507e-10, 1.396348e-10, 
    1.401837e-10, 1.407006e-10, 1.413045e-10, 1.361978e-10, 1.360216e-10, 
    1.363372e-10, 1.367737e-10, 1.371789e-10, 1.377175e-10, 1.377727e-10, 
    1.378736e-10, 1.38135e-10, 1.383548e-10, 1.379055e-10, 1.384099e-10, 
    1.365169e-10, 1.375088e-10, 1.35955e-10, 1.364228e-10, 1.36748e-10, 
    1.366054e-10, 1.373462e-10, 1.375209e-10, 1.382305e-10, 1.378637e-10, 
    1.400482e-10, 1.390816e-10, 1.417645e-10, 1.410146e-10, 1.359601e-10, 
    1.361972e-10, 1.370228e-10, 1.3663e-10, 1.377535e-10, 1.380301e-10, 
    1.38255e-10, 1.385424e-10, 1.385735e-10, 1.387438e-10, 1.384647e-10, 
    1.387327e-10, 1.377187e-10, 1.381718e-10, 1.369285e-10, 1.37231e-10, 
    1.370919e-10, 1.369392e-10, 1.374104e-10, 1.379125e-10, 1.379233e-10, 
    1.380843e-10, 1.38538e-10, 1.377581e-10, 1.401729e-10, 1.386814e-10, 
    1.364559e-10, 1.369128e-10, 1.369781e-10, 1.368011e-10, 1.380024e-10, 
    1.375671e-10, 1.387396e-10, 1.384227e-10, 1.38942e-10, 1.386839e-10, 
    1.38646e-10, 1.383146e-10, 1.381082e-10, 1.37587e-10, 1.37163e-10, 
    1.368268e-10, 1.369049e-10, 1.372743e-10, 1.379433e-10, 1.385762e-10, 
    1.384376e-10, 1.389025e-10, 1.37672e-10, 1.381879e-10, 1.379885e-10, 
    1.385085e-10, 1.373693e-10, 1.383393e-10, 1.371213e-10, 1.372281e-10, 
    1.375584e-10, 1.382229e-10, 1.3837e-10, 1.38527e-10, 1.384301e-10, 
    1.379603e-10, 1.378833e-10, 1.375504e-10, 1.374585e-10, 1.372048e-10, 
    1.369949e-10, 1.371867e-10, 1.373882e-10, 1.379605e-10, 1.384762e-10, 
    1.390386e-10, 1.391763e-10, 1.398334e-10, 1.392984e-10, 1.401812e-10, 
    1.394306e-10, 1.407301e-10, 1.383956e-10, 1.394086e-10, 1.375735e-10, 
    1.377711e-10, 1.381287e-10, 1.389489e-10, 1.385061e-10, 1.390239e-10, 
    1.378803e-10, 1.37287e-10, 1.371335e-10, 1.368472e-10, 1.371401e-10, 
    1.371163e-10, 1.373966e-10, 1.373065e-10, 1.379795e-10, 1.37618e-10, 
    1.38645e-10, 1.390199e-10, 1.400786e-10, 1.407278e-10, 1.413887e-10, 
    1.416805e-10, 1.417693e-10, 1.418065e-10 ;

 SOIL1N_vr =
  2.497618, 2.497612, 2.497613, 2.497607, 2.49761, 2.497607, 2.497617, 
    2.497611, 2.497615, 2.497617, 2.497597, 2.497607, 2.497587, 2.497593, 
    2.497577, 2.497588, 2.497575, 2.497578, 2.49757, 2.497572, 2.497563, 
    2.497569, 2.497558, 2.497565, 2.497564, 2.49757, 2.497605, 2.497598, 
    2.497606, 2.497605, 2.497605, 2.49761, 2.497613, 2.497618, 2.497617, 
    2.497613, 2.497604, 2.497607, 2.4976, 2.4976, 2.497591, 2.497595, 
    2.49758, 2.497584, 2.497572, 2.497576, 2.497572, 2.497573, 2.497572, 
    2.497577, 2.497575, 2.497579, 2.497594, 2.49759, 2.497603, 2.497611, 
    2.497616, 2.49762, 2.49762, 2.497619, 2.497613, 2.497608, 2.497605, 
    2.497602, 2.4976, 2.497592, 2.497588, 2.497579, 2.497581, 2.497578, 
    2.497576, 2.497571, 2.497572, 2.49757, 2.497578, 2.497573, 2.497582, 
    2.497579, 2.497599, 2.497607, 2.49761, 2.497612, 2.497619, 2.497615, 
    2.497616, 2.497612, 2.497609, 2.497611, 2.497602, 2.497605, 2.497588, 
    2.497596, 2.497576, 2.497581, 2.497575, 2.497578, 2.497573, 2.497577, 
    2.49757, 2.497568, 2.497569, 2.497565, 2.497578, 2.497572, 2.497611, 
    2.49761, 2.497609, 2.497614, 2.497614, 2.497618, 2.497615, 2.497613, 
    2.497609, 2.497607, 2.497604, 2.497599, 2.497594, 2.497586, 2.49758, 
    2.497577, 2.497579, 2.497577, 2.497579, 2.49758, 2.497568, 2.497575, 
    2.497565, 2.497566, 2.49757, 2.497566, 2.49761, 2.497612, 2.497616, 
    2.497612, 2.497619, 2.497615, 2.497613, 2.497605, 2.497604, 2.497602, 
    2.497599, 2.497595, 2.497587, 2.497581, 2.497576, 2.497576, 2.497576, 
    2.497575, 2.497578, 2.497574, 2.497573, 2.497575, 2.497566, 2.497568, 
    2.497566, 2.497567, 2.497611, 2.497609, 2.49761, 2.497608, 2.497609, 
    2.497602, 2.497601, 2.497591, 2.497595, 2.497588, 2.497594, 2.497593, 
    2.497588, 2.497594, 2.497582, 2.49759, 2.497575, 2.497583, 2.497574, 
    2.497576, 2.497573, 2.497571, 2.497568, 2.497562, 2.497563, 2.497559, 
    2.497606, 2.497603, 2.497603, 2.4976, 2.497598, 2.497593, 2.497586, 
    2.497589, 2.497583, 2.497582, 2.49759, 2.497585, 2.497601, 2.497598, 
    2.4976, 2.497606, 2.497588, 2.497597, 2.49758, 2.497585, 2.497571, 
    2.497578, 2.497564, 2.497558, 2.497553, 2.497546, 2.497601, 2.497603, 
    2.4976, 2.497595, 2.497591, 2.497585, 2.497584, 2.497583, 2.49758, 
    2.497578, 2.497583, 2.497577, 2.497598, 2.497587, 2.497604, 2.497599, 
    2.497595, 2.497597, 2.497589, 2.497587, 2.497579, 2.497583, 2.49756, 
    2.49757, 2.497541, 2.497549, 2.497604, 2.497601, 2.497592, 2.497597, 
    2.497585, 2.497581, 2.497579, 2.497576, 2.497576, 2.497574, 2.497577, 
    2.497574, 2.497585, 2.49758, 2.497593, 2.49759, 2.497592, 2.497593, 
    2.497588, 2.497583, 2.497583, 2.497581, 2.497576, 2.497584, 2.497558, 
    2.497574, 2.497599, 2.497594, 2.497593, 2.497595, 2.497582, 2.497586, 
    2.497574, 2.497577, 2.497572, 2.497574, 2.497575, 2.497578, 2.497581, 
    2.497586, 2.497591, 2.497595, 2.497594, 2.49759, 2.497582, 2.497576, 
    2.497577, 2.497572, 2.497585, 2.49758, 2.497582, 2.497576, 2.497589, 
    2.497578, 2.497591, 2.49759, 2.497586, 2.497579, 2.497578, 2.497576, 
    2.497577, 2.497582, 2.497583, 2.497587, 2.497588, 2.49759, 2.497593, 
    2.497591, 2.497588, 2.497582, 2.497577, 2.497571, 2.497569, 2.497562, 
    2.497568, 2.497558, 2.497566, 2.497552, 2.497577, 2.497566, 2.497586, 
    2.497584, 2.49758, 2.497571, 2.497576, 2.497571, 2.497583, 2.49759, 
    2.497591, 2.497594, 2.497591, 2.497591, 2.497588, 2.497589, 2.497582, 
    2.497586, 2.497575, 2.497571, 2.497559, 2.497552, 2.497545, 2.497542, 
    2.497541, 2.497541,
  2.497897, 2.49789, 2.497891, 2.497885, 2.497888, 2.497884, 2.497896, 
    2.497889, 2.497893, 2.497897, 2.497872, 2.497884, 2.497859, 2.497867, 
    2.497847, 2.49786, 2.497845, 2.497848, 2.497839, 2.497841, 2.49783, 
    2.497838, 2.497824, 2.497832, 2.49783, 2.497838, 2.497882, 2.497874, 
    2.497882, 2.497881, 2.497882, 2.497888, 2.497891, 2.497898, 2.497897, 
    2.497892, 2.49788, 2.497884, 2.497875, 2.497875, 2.497864, 2.497869, 
    2.497851, 2.497856, 2.497841, 2.497845, 2.497841, 2.497843, 2.497841, 
    2.497847, 2.497844, 2.497849, 2.497868, 2.497863, 2.497879, 2.497889, 
    2.497895, 2.4979, 2.4979, 2.497898, 2.497892, 2.497886, 2.497881, 
    2.497878, 2.497875, 2.497866, 2.497861, 2.49785, 2.497852, 2.497849, 
    2.497845, 2.49784, 2.497841, 2.497838, 2.497849, 2.497842, 2.497853, 
    2.49785, 2.497874, 2.497883, 2.497887, 2.497891, 2.497899, 2.497893, 
    2.497895, 2.49789, 2.497887, 2.497888, 2.497878, 2.497882, 2.49786, 
    2.49787, 2.497846, 2.497851, 2.497844, 2.497848, 2.497842, 2.497847, 
    2.497838, 2.497835, 2.497837, 2.497831, 2.497848, 2.497841, 2.497889, 
    2.497888, 2.497887, 2.497893, 2.497893, 2.497898, 2.497894, 2.497891, 
    2.497886, 2.497884, 2.497881, 2.497874, 2.497868, 2.497858, 2.497851, 
    2.497846, 2.497849, 2.497847, 2.497849, 2.497851, 2.497836, 2.497844, 
    2.497832, 2.497833, 2.497838, 2.497833, 2.497888, 2.49789, 2.497895, 
    2.497891, 2.497899, 2.497894, 2.497892, 2.497882, 2.49788, 2.497878, 
    2.497874, 2.497869, 2.49786, 2.497852, 2.497845, 2.497846, 2.497845, 
    2.497844, 2.497848, 2.497843, 2.497843, 2.497844, 2.497833, 2.497836, 
    2.497833, 2.497835, 2.497889, 2.497886, 2.497888, 2.497885, 2.497887, 
    2.497879, 2.497876, 2.497864, 2.497869, 2.497861, 2.497868, 2.497867, 
    2.497861, 2.497868, 2.497853, 2.497863, 2.497844, 2.497854, 2.497843, 
    2.497845, 2.497842, 2.497839, 2.497835, 2.497828, 2.49783, 2.497824, 
    2.497882, 2.497879, 2.497879, 2.497875, 2.497873, 2.497867, 2.497858, 
    2.497861, 2.497855, 2.497854, 2.497863, 2.497857, 2.497877, 2.497874, 
    2.497875, 2.497882, 2.49786, 2.497872, 2.497851, 2.497857, 2.497839, 
    2.497848, 2.497831, 2.497824, 2.497817, 2.497809, 2.497877, 2.497879, 
    2.497875, 2.497869, 2.497864, 2.497857, 2.497856, 2.497854, 2.497851, 
    2.497848, 2.497854, 2.497847, 2.497873, 2.497859, 2.49788, 2.497874, 
    2.49787, 2.497872, 2.497862, 2.497859, 2.49785, 2.497855, 2.497825, 
    2.497838, 2.497802, 2.497813, 2.49788, 2.497877, 2.497866, 2.497871, 
    2.497856, 2.497852, 2.497849, 2.497846, 2.497845, 2.497843, 2.497847, 
    2.497843, 2.497857, 2.497851, 2.497867, 2.497863, 2.497865, 2.497867, 
    2.497861, 2.497854, 2.497854, 2.497852, 2.497846, 2.497856, 2.497824, 
    2.497844, 2.497874, 2.497867, 2.497867, 2.497869, 2.497853, 2.497859, 
    2.497843, 2.497847, 2.49784, 2.497844, 2.497844, 2.497849, 2.497851, 
    2.497858, 2.497864, 2.497869, 2.497868, 2.497863, 2.497854, 2.497845, 
    2.497847, 2.497841, 2.497857, 2.49785, 2.497853, 2.497846, 2.497861, 
    2.497848, 2.497865, 2.497863, 2.497859, 2.49785, 2.497848, 2.497846, 
    2.497847, 2.497853, 2.497854, 2.497859, 2.49786, 2.497864, 2.497866, 
    2.497864, 2.497861, 2.497853, 2.497846, 2.497839, 2.497837, 2.497828, 
    2.497835, 2.497824, 2.497834, 2.497816, 2.497848, 2.497834, 2.497859, 
    2.497856, 2.497851, 2.49784, 2.497846, 2.497839, 2.497854, 2.497862, 
    2.497864, 2.497868, 2.497864, 2.497865, 2.497861, 2.497862, 2.497853, 
    2.497858, 2.497844, 2.497839, 2.497825, 2.497816, 2.497808, 2.497804, 
    2.497802, 2.497802,
  2.498027, 2.498018, 2.498019, 2.498012, 2.498016, 2.498012, 2.498025, 
    2.498018, 2.498022, 2.498026, 2.497999, 2.498012, 2.497985, 2.497993, 
    2.497972, 2.497986, 2.497969, 2.497972, 2.497962, 2.497965, 2.497952, 
    2.497961, 2.497946, 2.497955, 2.497953, 2.497961, 2.498009, 2.498, 
    2.49801, 2.498009, 2.498009, 2.498016, 2.49802, 2.498027, 2.498026, 
    2.49802, 2.498008, 2.498012, 2.498002, 2.498002, 2.49799, 2.497995, 
    2.497976, 2.497981, 2.497965, 2.497969, 2.497965, 2.497966, 2.497965, 
    2.497971, 2.497969, 2.497974, 2.497994, 2.497988, 2.498006, 2.498017, 
    2.498024, 2.49803, 2.498029, 2.498028, 2.49802, 2.498014, 2.498009, 
    2.498005, 2.498002, 2.497992, 2.497987, 2.497974, 2.497977, 2.497973, 
    2.49797, 2.497964, 2.497965, 2.497962, 2.497973, 2.497966, 2.497978, 
    2.497975, 2.498001, 2.498011, 2.498015, 2.498019, 2.498028, 2.498022, 
    2.498024, 2.498019, 2.498015, 2.498017, 2.498005, 2.49801, 2.497986, 
    2.497996, 2.49797, 2.497976, 2.497968, 2.497972, 2.497966, 2.497972, 
    2.497961, 2.497959, 2.49796, 2.497954, 2.497972, 2.497965, 2.498017, 
    2.498016, 2.498015, 2.498021, 2.498022, 2.498027, 2.498022, 2.49802, 
    2.498015, 2.498011, 2.498008, 2.498002, 2.497994, 2.497983, 2.497976, 
    2.497971, 2.497974, 2.497971, 2.497974, 2.497976, 2.49796, 2.497969, 
    2.497955, 2.497956, 2.497962, 2.497956, 2.498016, 2.498018, 2.498024, 
    2.498019, 2.498028, 2.498023, 2.49802, 2.498009, 2.498007, 2.498005, 
    2.498001, 2.497995, 2.497985, 2.497977, 2.497969, 2.49797, 2.49797, 
    2.497968, 2.497972, 2.497967, 2.497967, 2.497969, 2.497956, 2.49796, 
    2.497956, 2.497958, 2.498017, 2.498014, 2.498016, 2.498013, 2.498015, 
    2.498006, 2.498003, 2.49799, 2.497995, 2.497987, 2.497994, 2.497993, 
    2.497987, 2.497994, 2.497977, 2.497989, 2.497968, 2.497979, 2.497967, 
    2.497969, 2.497966, 2.497962, 2.497959, 2.497951, 2.497953, 2.497947, 
    2.49801, 2.498006, 2.498007, 2.498003, 2.498, 2.497993, 2.497983, 
    2.497987, 2.49798, 2.497978, 2.497989, 2.497983, 2.498004, 2.498, 
    2.498002, 2.49801, 2.497986, 2.497998, 2.497976, 2.497982, 2.497963, 
    2.497973, 2.497954, 2.497946, 2.497938, 2.497929, 2.498004, 2.498007, 
    2.498002, 2.497996, 2.49799, 2.497982, 2.497981, 2.49798, 2.497976, 
    2.497972, 2.497979, 2.497972, 2.497999, 2.497985, 2.498008, 2.498001, 
    2.497996, 2.497998, 2.497987, 2.497985, 2.497974, 2.49798, 2.497948, 
    2.497962, 2.497923, 2.497934, 2.498008, 2.498004, 2.497992, 2.497998, 
    2.497981, 2.497977, 2.497974, 2.49797, 2.497969, 2.497967, 2.497971, 
    2.497967, 2.497982, 2.497975, 2.497993, 2.497989, 2.497991, 2.497993, 
    2.497986, 2.497979, 2.497979, 2.497977, 2.49797, 2.497981, 2.497946, 
    2.497968, 2.498, 2.497994, 2.497993, 2.497995, 2.497978, 2.497984, 
    2.497967, 2.497972, 2.497964, 2.497968, 2.497968, 2.497973, 2.497976, 
    2.497984, 2.49799, 2.497995, 2.497994, 2.497988, 2.497979, 2.497969, 
    2.497971, 2.497965, 2.497983, 2.497975, 2.497978, 2.49797, 2.497987, 
    2.497973, 2.497991, 2.497989, 2.497984, 2.497974, 2.497972, 2.49797, 
    2.497972, 2.497978, 2.497979, 2.497984, 2.497986, 2.497989, 2.497993, 
    2.49799, 2.497987, 2.497978, 2.497971, 2.497962, 2.497961, 2.497951, 
    2.497959, 2.497946, 2.497957, 2.497938, 2.497972, 2.497957, 2.497984, 
    2.497981, 2.497976, 2.497964, 2.49797, 2.497963, 2.497979, 2.497988, 
    2.49799, 2.497995, 2.49799, 2.497991, 2.497987, 2.497988, 2.497978, 
    2.497983, 2.497968, 2.497963, 2.497947, 2.497938, 2.497928, 2.497924, 
    2.497923, 2.497922,
  2.498126, 2.498117, 2.498119, 2.498111, 2.498116, 2.498111, 2.498124, 
    2.498117, 2.498122, 2.498125, 2.498097, 2.498111, 2.498083, 2.498092, 
    2.49807, 2.498085, 2.498067, 2.49807, 2.49806, 2.498063, 2.49805, 
    2.498059, 2.498044, 2.498052, 2.498051, 2.498059, 2.498108, 2.498099, 
    2.498109, 2.498108, 2.498108, 2.498115, 2.498119, 2.498127, 2.498125, 
    2.49812, 2.498107, 2.498111, 2.498101, 2.498101, 2.498089, 2.498094, 
    2.498074, 2.49808, 2.498063, 2.498067, 2.498063, 2.498065, 2.498063, 
    2.49807, 2.498067, 2.498072, 2.498093, 2.498087, 2.498105, 2.498116, 
    2.498124, 2.498129, 2.498128, 2.498127, 2.49812, 2.498113, 2.498108, 
    2.498104, 2.498101, 2.498091, 2.498085, 2.498073, 2.498075, 2.498071, 
    2.498068, 2.498062, 2.498063, 2.49806, 2.498071, 2.498064, 2.498076, 
    2.498073, 2.4981, 2.49811, 2.498115, 2.498118, 2.498128, 2.498121, 
    2.498124, 2.498118, 2.498114, 2.498116, 2.498104, 2.498109, 2.498085, 
    2.498095, 2.498068, 2.498075, 2.498067, 2.498071, 2.498064, 2.49807, 
    2.498059, 2.498057, 2.498058, 2.498052, 2.49807, 2.498063, 2.498116, 
    2.498116, 2.498114, 2.498121, 2.498121, 2.498127, 2.498122, 2.498119, 
    2.498114, 2.498111, 2.498107, 2.4981, 2.498093, 2.498082, 2.498074, 
    2.498069, 2.498072, 2.498069, 2.498073, 2.498074, 2.498058, 2.498067, 
    2.498053, 2.498054, 2.49806, 2.498054, 2.498115, 2.498117, 2.498123, 
    2.498118, 2.498127, 2.498122, 2.49812, 2.498109, 2.498106, 2.498104, 
    2.4981, 2.498094, 2.498084, 2.498075, 2.498068, 2.498068, 2.498068, 
    2.498066, 2.49807, 2.498065, 2.498065, 2.498067, 2.498054, 2.498058, 
    2.498054, 2.498056, 2.498116, 2.498114, 2.498115, 2.498112, 2.498114, 
    2.498105, 2.498102, 2.498089, 2.498094, 2.498085, 2.498093, 2.498092, 
    2.498085, 2.498093, 2.498076, 2.498087, 2.498066, 2.498077, 2.498065, 
    2.498068, 2.498064, 2.498061, 2.498057, 2.498049, 2.498051, 2.498044, 
    2.498109, 2.498105, 2.498106, 2.498101, 2.498099, 2.498092, 2.498081, 
    2.498085, 2.498078, 2.498077, 2.498088, 2.498081, 2.498103, 2.498099, 
    2.498101, 2.498109, 2.498085, 2.498097, 2.498074, 2.498081, 2.498061, 
    2.498071, 2.498052, 2.498044, 2.498036, 2.498027, 2.498103, 2.498106, 
    2.498101, 2.498095, 2.498088, 2.49808, 2.49808, 2.498078, 2.498074, 
    2.498071, 2.498078, 2.49807, 2.498098, 2.498084, 2.498107, 2.4981, 
    2.498095, 2.498097, 2.498086, 2.498083, 2.498073, 2.498078, 2.498045, 
    2.49806, 2.49802, 2.498031, 2.498107, 2.498103, 2.498091, 2.498097, 
    2.49808, 2.498076, 2.498072, 2.498068, 2.498068, 2.498065, 2.498069, 
    2.498065, 2.49808, 2.498074, 2.498092, 2.498088, 2.49809, 2.498092, 
    2.498085, 2.498077, 2.498077, 2.498075, 2.498068, 2.49808, 2.498044, 
    2.498066, 2.498099, 2.498092, 2.498091, 2.498094, 2.498076, 2.498083, 
    2.498065, 2.49807, 2.498062, 2.498066, 2.498066, 2.498071, 2.498075, 
    2.498082, 2.498089, 2.498094, 2.498092, 2.498087, 2.498077, 2.498068, 
    2.49807, 2.498063, 2.498081, 2.498073, 2.498076, 2.498069, 2.498085, 
    2.498071, 2.498089, 2.498088, 2.498083, 2.498073, 2.498071, 2.498068, 
    2.49807, 2.498077, 2.498078, 2.498083, 2.498084, 2.498088, 2.498091, 
    2.498088, 2.498085, 2.498077, 2.498069, 2.498061, 2.498059, 2.498049, 
    2.498057, 2.498044, 2.498055, 2.498035, 2.49807, 2.498055, 2.498083, 
    2.49808, 2.498074, 2.498062, 2.498069, 2.498061, 2.498078, 2.498087, 
    2.498089, 2.498093, 2.498089, 2.498089, 2.498085, 2.498086, 2.498076, 
    2.498082, 2.498066, 2.498061, 2.498045, 2.498035, 2.498025, 2.498021, 
    2.49802, 2.498019,
  2.498263, 2.498255, 2.498256, 2.49825, 2.498253, 2.498249, 2.498261, 
    2.498254, 2.498259, 2.498262, 2.498237, 2.498249, 2.498224, 2.498232, 
    2.498212, 2.498225, 2.498209, 2.498212, 2.498203, 2.498206, 2.498194, 
    2.498202, 2.498188, 2.498196, 2.498194, 2.498202, 2.498247, 2.498238, 
    2.498247, 2.498246, 2.498247, 2.498253, 2.498256, 2.498263, 2.498262, 
    2.498257, 2.498245, 2.49825, 2.49824, 2.49824, 2.498229, 2.498234, 
    2.498215, 2.498221, 2.498205, 2.498209, 2.498206, 2.498207, 2.498206, 
    2.498211, 2.498209, 2.498214, 2.498233, 2.498227, 2.498244, 2.498254, 
    2.498261, 2.498266, 2.498265, 2.498264, 2.498257, 2.498251, 2.498246, 
    2.498243, 2.49824, 2.49823, 2.498225, 2.498214, 2.498216, 2.498213, 
    2.49821, 2.498204, 2.498205, 2.498203, 2.498213, 2.498206, 2.498218, 
    2.498214, 2.498239, 2.498248, 2.498252, 2.498256, 2.498264, 2.498259, 
    2.498261, 2.498255, 2.498252, 2.498254, 2.498243, 2.498247, 2.498225, 
    2.498235, 2.49821, 2.498216, 2.498209, 2.498212, 2.498206, 2.498212, 
    2.498202, 2.4982, 2.498201, 2.498195, 2.498212, 2.498206, 2.498254, 
    2.498253, 2.498252, 2.498258, 2.498258, 2.498263, 2.498259, 2.498257, 
    2.498252, 2.498249, 2.498246, 2.49824, 2.498232, 2.498223, 2.498216, 
    2.498211, 2.498214, 2.498211, 2.498214, 2.498215, 2.4982, 2.498209, 
    2.498196, 2.498197, 2.498203, 2.498197, 2.498253, 2.498255, 2.49826, 
    2.498256, 2.498264, 2.49826, 2.498257, 2.498247, 2.498245, 2.498243, 
    2.498239, 2.498234, 2.498224, 2.498217, 2.498209, 2.49821, 2.49821, 
    2.498208, 2.498212, 2.498208, 2.498207, 2.498209, 2.498197, 2.4982, 
    2.498197, 2.498199, 2.498254, 2.498251, 2.498253, 2.49825, 2.498252, 
    2.498244, 2.498241, 2.498229, 2.498234, 2.498226, 2.498233, 2.498232, 
    2.498225, 2.498233, 2.498217, 2.498228, 2.498208, 2.498219, 2.498208, 
    2.498209, 2.498206, 2.498203, 2.498199, 2.498193, 2.498194, 2.498188, 
    2.498247, 2.498244, 2.498244, 2.49824, 2.498238, 2.498232, 2.498222, 
    2.498226, 2.498219, 2.498218, 2.498228, 2.498222, 2.498241, 2.498238, 
    2.49824, 2.498247, 2.498225, 2.498236, 2.498215, 2.498222, 2.498204, 
    2.498213, 2.498195, 2.498188, 2.49818, 2.498172, 2.498242, 2.498244, 
    2.49824, 2.498234, 2.498229, 2.498221, 2.49822, 2.498219, 2.498215, 
    2.498213, 2.498219, 2.498212, 2.498238, 2.498224, 2.498245, 2.498239, 
    2.498235, 2.498236, 2.498226, 2.498224, 2.498214, 2.498219, 2.498189, 
    2.498203, 2.498166, 2.498176, 2.498245, 2.498242, 2.498231, 2.498236, 
    2.498221, 2.498217, 2.498214, 2.49821, 2.498209, 2.498207, 2.498211, 
    2.498207, 2.498221, 2.498215, 2.498232, 2.498228, 2.49823, 2.498232, 
    2.498225, 2.498219, 2.498219, 2.498216, 2.49821, 2.498221, 2.498188, 
    2.498208, 2.498239, 2.498232, 2.498231, 2.498234, 2.498217, 2.498223, 
    2.498207, 2.498212, 2.498204, 2.498208, 2.498209, 2.498213, 2.498216, 
    2.498223, 2.498229, 2.498233, 2.498232, 2.498227, 2.498218, 2.498209, 
    2.498211, 2.498205, 2.498222, 2.498215, 2.498218, 2.49821, 2.498226, 
    2.498213, 2.498229, 2.498228, 2.498223, 2.498214, 2.498212, 2.49821, 
    2.498212, 2.498218, 2.498219, 2.498224, 2.498225, 2.498228, 2.498231, 
    2.498229, 2.498226, 2.498218, 2.498211, 2.498203, 2.498201, 2.498192, 
    2.4982, 2.498188, 2.498198, 2.49818, 2.498212, 2.498198, 2.498223, 
    2.49822, 2.498216, 2.498204, 2.49821, 2.498204, 2.498219, 2.498227, 
    2.498229, 2.498233, 2.498229, 2.49823, 2.498226, 2.498227, 2.498218, 
    2.498223, 2.498209, 2.498204, 2.498189, 2.49818, 2.498171, 2.498167, 
    2.498166, 2.498165,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  5.981638e-08, 6.008199e-08, 6.003036e-08, 6.02446e-08, 6.012576e-08, 
    6.026604e-08, 5.987024e-08, 6.009252e-08, 5.995062e-08, 5.98403e-08, 
    6.06604e-08, 6.025416e-08, 6.108253e-08, 6.082337e-08, 6.147447e-08, 
    6.104219e-08, 6.156164e-08, 6.146202e-08, 6.176194e-08, 6.167601e-08, 
    6.205964e-08, 6.18016e-08, 6.225856e-08, 6.199802e-08, 6.203877e-08, 
    6.179308e-08, 6.033592e-08, 6.060981e-08, 6.031969e-08, 6.035874e-08, 
    6.034122e-08, 6.01282e-08, 6.002085e-08, 5.979609e-08, 5.98369e-08, 
    6.000199e-08, 6.037631e-08, 6.024924e-08, 6.056951e-08, 6.056229e-08, 
    6.091889e-08, 6.07581e-08, 6.135755e-08, 6.118717e-08, 6.167959e-08, 
    6.155575e-08, 6.167377e-08, 6.163799e-08, 6.167424e-08, 6.149261e-08, 
    6.157043e-08, 6.14106e-08, 6.07882e-08, 6.09711e-08, 6.042565e-08, 
    6.009773e-08, 5.987998e-08, 5.972547e-08, 5.974731e-08, 5.978895e-08, 
    6.000295e-08, 6.020419e-08, 6.035756e-08, 6.046015e-08, 6.056124e-08, 
    6.086724e-08, 6.102924e-08, 6.1392e-08, 6.132655e-08, 6.143745e-08, 
    6.154342e-08, 6.172134e-08, 6.169206e-08, 6.177044e-08, 6.143453e-08, 
    6.165777e-08, 6.128926e-08, 6.139004e-08, 6.058868e-08, 6.028353e-08, 
    6.015379e-08, 6.004028e-08, 5.97641e-08, 5.995481e-08, 5.987963e-08, 
    6.005851e-08, 6.017218e-08, 6.011597e-08, 6.046295e-08, 6.032805e-08, 
    6.103884e-08, 6.073265e-08, 6.153106e-08, 6.133998e-08, 6.157686e-08, 
    6.145599e-08, 6.16631e-08, 6.14767e-08, 6.179962e-08, 6.186993e-08, 
    6.182188e-08, 6.200649e-08, 6.146637e-08, 6.167377e-08, 6.011439e-08, 
    6.012355e-08, 6.016627e-08, 5.99785e-08, 5.996701e-08, 5.979497e-08, 
    5.994806e-08, 6.001325e-08, 6.017877e-08, 6.027668e-08, 6.036975e-08, 
    6.05744e-08, 6.080298e-08, 6.112266e-08, 6.135237e-08, 6.150636e-08, 
    6.141194e-08, 6.149529e-08, 6.14021e-08, 6.135843e-08, 6.184358e-08, 
    6.157115e-08, 6.197993e-08, 6.195732e-08, 6.17723e-08, 6.195986e-08, 
    6.012999e-08, 6.007723e-08, 5.989406e-08, 6.003741e-08, 5.977623e-08, 
    5.992241e-08, 6.000648e-08, 6.033085e-08, 6.040214e-08, 6.046823e-08, 
    6.059878e-08, 6.076632e-08, 6.106026e-08, 6.131605e-08, 6.154959e-08, 
    6.153248e-08, 6.15385e-08, 6.159067e-08, 6.146144e-08, 6.161189e-08, 
    6.163714e-08, 6.157112e-08, 6.195428e-08, 6.184481e-08, 6.195683e-08, 
    6.188556e-08, 6.009439e-08, 6.018316e-08, 6.013519e-08, 6.02254e-08, 
    6.016185e-08, 6.044446e-08, 6.05292e-08, 6.092577e-08, 6.076302e-08, 
    6.102206e-08, 6.078934e-08, 6.083057e-08, 6.103049e-08, 6.080192e-08, 
    6.130193e-08, 6.096291e-08, 6.159269e-08, 6.125408e-08, 6.161392e-08, 
    6.154858e-08, 6.165677e-08, 6.175366e-08, 6.187557e-08, 6.210053e-08, 
    6.204844e-08, 6.223657e-08, 6.031553e-08, 6.043068e-08, 6.042055e-08, 
    6.054108e-08, 6.063021e-08, 6.082344e-08, 6.113338e-08, 6.101683e-08, 
    6.123081e-08, 6.127377e-08, 6.094868e-08, 6.114826e-08, 6.050777e-08, 
    6.061122e-08, 6.054963e-08, 6.032461e-08, 6.104366e-08, 6.067461e-08, 
    6.135616e-08, 6.11562e-08, 6.173984e-08, 6.144956e-08, 6.201976e-08, 
    6.226353e-08, 6.249304e-08, 6.276121e-08, 6.049354e-08, 6.04153e-08, 
    6.055541e-08, 6.074928e-08, 6.09292e-08, 6.116839e-08, 6.119287e-08, 
    6.123769e-08, 6.135377e-08, 6.145138e-08, 6.125185e-08, 6.147585e-08, 
    6.063521e-08, 6.107571e-08, 6.03857e-08, 6.059344e-08, 6.073785e-08, 
    6.067452e-08, 6.10035e-08, 6.108105e-08, 6.139619e-08, 6.123328e-08, 
    6.220336e-08, 6.177412e-08, 6.296546e-08, 6.263246e-08, 6.038795e-08, 
    6.049328e-08, 6.085988e-08, 6.068545e-08, 6.118437e-08, 6.130718e-08, 
    6.140704e-08, 6.153468e-08, 6.154847e-08, 6.16241e-08, 6.150017e-08, 
    6.161921e-08, 6.11689e-08, 6.137012e-08, 6.081799e-08, 6.095235e-08, 
    6.089054e-08, 6.082274e-08, 6.103202e-08, 6.125498e-08, 6.125976e-08, 
    6.133126e-08, 6.153272e-08, 6.118639e-08, 6.225874e-08, 6.15964e-08, 
    6.060814e-08, 6.081102e-08, 6.084002e-08, 6.076142e-08, 6.129487e-08, 
    6.110157e-08, 6.162226e-08, 6.148153e-08, 6.171212e-08, 6.159753e-08, 
    6.158067e-08, 6.143351e-08, 6.134189e-08, 6.111043e-08, 6.092213e-08, 
    6.077283e-08, 6.080754e-08, 6.097154e-08, 6.126863e-08, 6.154971e-08, 
    6.148814e-08, 6.16946e-08, 6.114819e-08, 6.137729e-08, 6.128873e-08, 
    6.151964e-08, 6.101373e-08, 6.144449e-08, 6.090362e-08, 6.095105e-08, 
    6.109773e-08, 6.139281e-08, 6.145812e-08, 6.152784e-08, 6.148482e-08, 
    6.127618e-08, 6.124199e-08, 6.109417e-08, 6.105335e-08, 6.094072e-08, 
    6.084748e-08, 6.093267e-08, 6.102213e-08, 6.127626e-08, 6.15053e-08, 
    6.175504e-08, 6.181617e-08, 6.210796e-08, 6.187041e-08, 6.226242e-08, 
    6.192911e-08, 6.250615e-08, 6.146948e-08, 6.191932e-08, 6.110441e-08, 
    6.119219e-08, 6.135096e-08, 6.171517e-08, 6.151856e-08, 6.174851e-08, 
    6.124066e-08, 6.09772e-08, 6.090905e-08, 6.07819e-08, 6.091197e-08, 
    6.090139e-08, 6.102585e-08, 6.098585e-08, 6.12847e-08, 6.112417e-08, 
    6.158024e-08, 6.17467e-08, 6.221686e-08, 6.250511e-08, 6.279861e-08, 
    6.292818e-08, 6.296762e-08, 6.298411e-08 ;

 SOIL1_HR_S3 =
  7.098643e-10, 7.130175e-10, 7.124045e-10, 7.149479e-10, 7.135371e-10, 
    7.152025e-10, 7.105036e-10, 7.131426e-10, 7.114579e-10, 7.101482e-10, 
    7.198844e-10, 7.150615e-10, 7.248961e-10, 7.218193e-10, 7.295494e-10, 
    7.244172e-10, 7.305844e-10, 7.294016e-10, 7.329624e-10, 7.319423e-10, 
    7.364971e-10, 7.334333e-10, 7.388588e-10, 7.357655e-10, 7.362492e-10, 
    7.333322e-10, 7.160322e-10, 7.192839e-10, 7.158394e-10, 7.163031e-10, 
    7.160951e-10, 7.135662e-10, 7.122917e-10, 7.096234e-10, 7.101078e-10, 
    7.120677e-10, 7.165116e-10, 7.150032e-10, 7.188055e-10, 7.187196e-10, 
    7.229533e-10, 7.210443e-10, 7.281614e-10, 7.261384e-10, 7.319848e-10, 
    7.305144e-10, 7.319158e-10, 7.314908e-10, 7.319212e-10, 7.297647e-10, 
    7.306886e-10, 7.287911e-10, 7.214017e-10, 7.235731e-10, 7.170975e-10, 
    7.132044e-10, 7.106193e-10, 7.087849e-10, 7.090442e-10, 7.095385e-10, 
    7.120792e-10, 7.144683e-10, 7.16289e-10, 7.17507e-10, 7.187073e-10, 
    7.223401e-10, 7.242635e-10, 7.285704e-10, 7.277932e-10, 7.291099e-10, 
    7.303681e-10, 7.324804e-10, 7.321327e-10, 7.330634e-10, 7.290753e-10, 
    7.317257e-10, 7.273505e-10, 7.285471e-10, 7.19033e-10, 7.154101e-10, 
    7.1387e-10, 7.125223e-10, 7.092436e-10, 7.115077e-10, 7.106152e-10, 
    7.127388e-10, 7.140882e-10, 7.134209e-10, 7.175404e-10, 7.159387e-10, 
    7.243774e-10, 7.207422e-10, 7.302213e-10, 7.279528e-10, 7.307651e-10, 
    7.2933e-10, 7.31789e-10, 7.29576e-10, 7.334098e-10, 7.342447e-10, 
    7.336741e-10, 7.358659e-10, 7.294533e-10, 7.319157e-10, 7.134022e-10, 
    7.13511e-10, 7.140181e-10, 7.117889e-10, 7.116526e-10, 7.096101e-10, 
    7.114275e-10, 7.122015e-10, 7.141665e-10, 7.153288e-10, 7.164338e-10, 
    7.188635e-10, 7.215772e-10, 7.253726e-10, 7.280998e-10, 7.29928e-10, 
    7.28807e-10, 7.297967e-10, 7.286903e-10, 7.281718e-10, 7.339317e-10, 
    7.306973e-10, 7.355507e-10, 7.352821e-10, 7.330855e-10, 7.353124e-10, 
    7.135874e-10, 7.129611e-10, 7.107864e-10, 7.124882e-10, 7.093877e-10, 
    7.111231e-10, 7.12121e-10, 7.15972e-10, 7.168184e-10, 7.17603e-10, 
    7.191528e-10, 7.21142e-10, 7.246317e-10, 7.276685e-10, 7.304413e-10, 
    7.302381e-10, 7.303097e-10, 7.30929e-10, 7.293948e-10, 7.311809e-10, 
    7.314807e-10, 7.306969e-10, 7.352461e-10, 7.339464e-10, 7.352764e-10, 
    7.344301e-10, 7.131647e-10, 7.142186e-10, 7.136491e-10, 7.147201e-10, 
    7.139656e-10, 7.173207e-10, 7.183268e-10, 7.23035e-10, 7.211028e-10, 
    7.241782e-10, 7.214152e-10, 7.219048e-10, 7.242783e-10, 7.215646e-10, 
    7.27501e-10, 7.234759e-10, 7.309531e-10, 7.269329e-10, 7.312051e-10, 
    7.304293e-10, 7.317138e-10, 7.328642e-10, 7.343117e-10, 7.369824e-10, 
    7.36364e-10, 7.385978e-10, 7.1579e-10, 7.171572e-10, 7.170369e-10, 
    7.184678e-10, 7.195261e-10, 7.218201e-10, 7.254998e-10, 7.24116e-10, 
    7.266565e-10, 7.271665e-10, 7.23307e-10, 7.256765e-10, 7.180723e-10, 
    7.193006e-10, 7.185694e-10, 7.158978e-10, 7.244347e-10, 7.200532e-10, 
    7.281448e-10, 7.257707e-10, 7.327001e-10, 7.292537e-10, 7.360235e-10, 
    7.389179e-10, 7.416427e-10, 7.448269e-10, 7.179035e-10, 7.169745e-10, 
    7.18638e-10, 7.209396e-10, 7.230757e-10, 7.259155e-10, 7.262062e-10, 
    7.267382e-10, 7.281165e-10, 7.292753e-10, 7.269063e-10, 7.295659e-10, 
    7.195853e-10, 7.248152e-10, 7.166232e-10, 7.190895e-10, 7.20804e-10, 
    7.20052e-10, 7.239579e-10, 7.248785e-10, 7.2862e-10, 7.266859e-10, 
    7.382034e-10, 7.331071e-10, 7.47252e-10, 7.432982e-10, 7.166499e-10, 
    7.179004e-10, 7.222528e-10, 7.201818e-10, 7.261052e-10, 7.275633e-10, 
    7.287489e-10, 7.302643e-10, 7.304281e-10, 7.31326e-10, 7.298546e-10, 
    7.312679e-10, 7.259215e-10, 7.283106e-10, 7.217554e-10, 7.233506e-10, 
    7.226167e-10, 7.218118e-10, 7.242964e-10, 7.269436e-10, 7.270003e-10, 
    7.278492e-10, 7.30241e-10, 7.261292e-10, 7.388609e-10, 7.309971e-10, 
    7.19264e-10, 7.216727e-10, 7.220169e-10, 7.210838e-10, 7.274171e-10, 
    7.251221e-10, 7.313041e-10, 7.296332e-10, 7.323711e-10, 7.310105e-10, 
    7.308104e-10, 7.290631e-10, 7.279753e-10, 7.252273e-10, 7.229917e-10, 
    7.212192e-10, 7.216314e-10, 7.235785e-10, 7.271055e-10, 7.304428e-10, 
    7.297117e-10, 7.321629e-10, 7.256756e-10, 7.283956e-10, 7.273442e-10, 
    7.300857e-10, 7.240793e-10, 7.291935e-10, 7.227721e-10, 7.233351e-10, 
    7.250766e-10, 7.2858e-10, 7.293554e-10, 7.30183e-10, 7.296723e-10, 
    7.271951e-10, 7.267894e-10, 7.250343e-10, 7.245496e-10, 7.232125e-10, 
    7.221055e-10, 7.231169e-10, 7.241791e-10, 7.271962e-10, 7.299155e-10, 
    7.328805e-10, 7.336063e-10, 7.370708e-10, 7.342503e-10, 7.389047e-10, 
    7.349473e-10, 7.417985e-10, 7.294902e-10, 7.348311e-10, 7.251559e-10, 
    7.261981e-10, 7.280831e-10, 7.324072e-10, 7.300729e-10, 7.32803e-10, 
    7.267735e-10, 7.236456e-10, 7.228366e-10, 7.213269e-10, 7.228711e-10, 
    7.227455e-10, 7.242232e-10, 7.237483e-10, 7.272964e-10, 7.253905e-10, 
    7.308053e-10, 7.327816e-10, 7.383636e-10, 7.417861e-10, 7.452708e-10, 
    7.468094e-10, 7.472777e-10, 7.474735e-10 ;

 SOIL2C =
  5.783958, 5.783965, 5.783963, 5.783968, 5.783966, 5.783968, 5.783959, 
    5.783965, 5.783961, 5.783959, 5.783978, 5.783968, 5.783987, 5.783981, 
    5.783996, 5.783986, 5.783998, 5.783996, 5.784003, 5.784001, 5.784009, 
    5.784004, 5.784014, 5.784008, 5.784009, 5.784003, 5.78397, 5.783977, 
    5.78397, 5.783971, 5.78397, 5.783966, 5.783963, 5.783958, 5.783959, 
    5.783963, 5.783971, 5.783968, 5.783976, 5.783976, 5.783984, 5.78398, 
    5.783993, 5.783989, 5.784001, 5.783998, 5.784001, 5.784, 5.784001, 
    5.783997, 5.783998, 5.783995, 5.78398, 5.783985, 5.783972, 5.783965, 
    5.78396, 5.783957, 5.783957, 5.783958, 5.783963, 5.783967, 5.783971, 
    5.783973, 5.783975, 5.783982, 5.783986, 5.783994, 5.783993, 5.783995, 
    5.783998, 5.784002, 5.784001, 5.784003, 5.783995, 5.784, 5.783992, 
    5.783994, 5.783976, 5.783969, 5.783966, 5.783964, 5.783957, 5.783961, 
    5.78396, 5.783964, 5.783967, 5.783965, 5.783973, 5.78397, 5.783986, 
    5.783979, 5.783998, 5.783993, 5.783998, 5.783996, 5.784, 5.783996, 
    5.784004, 5.784005, 5.784004, 5.784008, 5.783996, 5.784001, 5.783965, 
    5.783966, 5.783967, 5.783962, 5.783962, 5.783958, 5.783961, 5.783963, 
    5.783967, 5.783969, 5.783971, 5.783976, 5.783981, 5.783988, 5.783993, 
    5.783997, 5.783995, 5.783997, 5.783995, 5.783994, 5.784005, 5.783998, 
    5.784008, 5.784007, 5.784003, 5.784007, 5.783966, 5.783964, 5.78396, 
    5.783963, 5.783957, 5.783961, 5.783963, 5.78397, 5.783972, 5.783973, 
    5.783976, 5.78398, 5.783987, 5.783993, 5.783998, 5.783998, 5.783998, 
    5.783999, 5.783996, 5.783999, 5.784, 5.783998, 5.784007, 5.784005, 
    5.784007, 5.784006, 5.783965, 5.783967, 5.783966, 5.783967, 5.783966, 
    5.783973, 5.783975, 5.783984, 5.78398, 5.783986, 5.78398, 5.783981, 
    5.783986, 5.783981, 5.783992, 5.783985, 5.783999, 5.783991, 5.783999, 
    5.783998, 5.784, 5.784002, 5.784005, 5.78401, 5.784009, 5.784013, 
    5.78397, 5.783972, 5.783972, 5.783975, 5.783977, 5.783981, 5.783988, 
    5.783986, 5.78399, 5.783991, 5.783984, 5.783989, 5.783974, 5.783977, 
    5.783975, 5.78397, 5.783987, 5.783978, 5.783993, 5.783989, 5.784002, 
    5.783996, 5.784009, 5.784014, 5.784019, 5.784026, 5.783974, 5.783972, 
    5.783975, 5.783979, 5.783984, 5.783989, 5.78399, 5.783991, 5.783993, 
    5.783996, 5.783991, 5.783996, 5.783977, 5.783987, 5.783971, 5.783976, 
    5.783979, 5.783978, 5.783986, 5.783987, 5.783994, 5.783991, 5.784013, 
    5.784003, 5.78403, 5.784022, 5.783971, 5.783974, 5.783982, 5.783978, 
    5.783989, 5.783992, 5.783995, 5.783998, 5.783998, 5.783999, 5.783997, 
    5.783999, 5.783989, 5.783994, 5.783981, 5.783984, 5.783983, 5.783981, 
    5.783986, 5.783991, 5.783991, 5.783993, 5.783998, 5.783989, 5.784014, 
    5.783999, 5.783977, 5.783981, 5.783982, 5.78398, 5.783992, 5.783988, 
    5.783999, 5.783996, 5.784001, 5.783999, 5.783998, 5.783995, 5.783993, 
    5.783988, 5.783984, 5.78398, 5.783981, 5.783985, 5.783991, 5.783998, 
    5.783997, 5.784001, 5.783988, 5.783994, 5.783992, 5.783997, 5.783986, 
    5.783996, 5.783983, 5.783984, 5.783988, 5.783994, 5.783996, 5.783998, 
    5.783997, 5.783992, 5.783991, 5.783988, 5.783987, 5.783984, 5.783982, 
    5.783984, 5.783986, 5.783992, 5.783997, 5.784002, 5.784004, 5.78401, 
    5.784005, 5.784014, 5.784007, 5.784019, 5.783996, 5.784006, 5.783988, 
    5.78399, 5.783993, 5.784002, 5.783997, 5.784002, 5.783991, 5.783985, 
    5.783983, 5.78398, 5.783983, 5.783983, 5.783986, 5.783985, 5.783992, 
    5.783988, 5.783998, 5.784002, 5.784013, 5.784019, 5.784026, 5.784029, 
    5.78403, 5.78403 ;

 SOIL2C_TO_SOIL1C =
  1.058223e-09, 1.062926e-09, 1.062012e-09, 1.065804e-09, 1.0637e-09, 
    1.066184e-09, 1.059177e-09, 1.063112e-09, 1.0606e-09, 1.058647e-09, 
    1.073166e-09, 1.065974e-09, 1.080639e-09, 1.076051e-09, 1.087578e-09, 
    1.079925e-09, 1.089122e-09, 1.087358e-09, 1.092668e-09, 1.091147e-09, 
    1.097939e-09, 1.09337e-09, 1.10146e-09, 1.096848e-09, 1.097569e-09, 
    1.093219e-09, 1.067421e-09, 1.07227e-09, 1.067134e-09, 1.067825e-09, 
    1.067515e-09, 1.063744e-09, 1.061843e-09, 1.057864e-09, 1.058587e-09, 
    1.061509e-09, 1.068136e-09, 1.065887e-09, 1.071557e-09, 1.071429e-09, 
    1.077742e-09, 1.074896e-09, 1.085509e-09, 1.082492e-09, 1.09121e-09, 
    1.089017e-09, 1.091107e-09, 1.090473e-09, 1.091115e-09, 1.087899e-09, 
    1.089277e-09, 1.086448e-09, 1.075429e-09, 1.078666e-09, 1.06901e-09, 
    1.063204e-09, 1.059349e-09, 1.056614e-09, 1.057e-09, 1.057738e-09, 
    1.061526e-09, 1.065089e-09, 1.067804e-09, 1.069621e-09, 1.07141e-09, 
    1.076828e-09, 1.079696e-09, 1.086118e-09, 1.08496e-09, 1.086923e-09, 
    1.088799e-09, 1.091949e-09, 1.091431e-09, 1.092818e-09, 1.086871e-09, 
    1.090824e-09, 1.084299e-09, 1.086084e-09, 1.071896e-09, 1.066494e-09, 
    1.064197e-09, 1.062187e-09, 1.057298e-09, 1.060674e-09, 1.059343e-09, 
    1.06251e-09, 1.064522e-09, 1.063527e-09, 1.06967e-09, 1.067282e-09, 
    1.079866e-09, 1.074445e-09, 1.08858e-09, 1.085197e-09, 1.089391e-09, 
    1.087251e-09, 1.090918e-09, 1.087618e-09, 1.093335e-09, 1.09458e-09, 
    1.093729e-09, 1.096997e-09, 1.087435e-09, 1.091107e-09, 1.063499e-09, 
    1.063661e-09, 1.064418e-09, 1.061094e-09, 1.06089e-09, 1.057844e-09, 
    1.060555e-09, 1.061709e-09, 1.064639e-09, 1.066372e-09, 1.06802e-09, 
    1.071643e-09, 1.07569e-09, 1.08135e-09, 1.085417e-09, 1.088143e-09, 
    1.086471e-09, 1.087947e-09, 1.086297e-09, 1.085524e-09, 1.094113e-09, 
    1.08929e-09, 1.096527e-09, 1.096127e-09, 1.092851e-09, 1.096172e-09, 
    1.063776e-09, 1.062841e-09, 1.059598e-09, 1.062136e-09, 1.057513e-09, 
    1.060101e-09, 1.061589e-09, 1.067332e-09, 1.068594e-09, 1.069764e-09, 
    1.072075e-09, 1.075041e-09, 1.080245e-09, 1.084774e-09, 1.088908e-09, 
    1.088605e-09, 1.088712e-09, 1.089636e-09, 1.087348e-09, 1.090011e-09, 
    1.090458e-09, 1.08929e-09, 1.096073e-09, 1.094135e-09, 1.096118e-09, 
    1.094856e-09, 1.063145e-09, 1.064717e-09, 1.063868e-09, 1.065465e-09, 
    1.064339e-09, 1.069343e-09, 1.070843e-09, 1.077864e-09, 1.074983e-09, 
    1.079569e-09, 1.075449e-09, 1.076179e-09, 1.079718e-09, 1.075671e-09, 
    1.084524e-09, 1.078522e-09, 1.089672e-09, 1.083677e-09, 1.090047e-09, 
    1.088891e-09, 1.090806e-09, 1.092521e-09, 1.09468e-09, 1.098662e-09, 
    1.09774e-09, 1.101071e-09, 1.06706e-09, 1.069099e-09, 1.06892e-09, 
    1.071053e-09, 1.072632e-09, 1.076052e-09, 1.08154e-09, 1.079476e-09, 
    1.083264e-09, 1.084025e-09, 1.07827e-09, 1.081803e-09, 1.070464e-09, 
    1.072295e-09, 1.071205e-09, 1.067221e-09, 1.079951e-09, 1.073417e-09, 
    1.085484e-09, 1.081944e-09, 1.092277e-09, 1.087137e-09, 1.097232e-09, 
    1.101548e-09, 1.105611e-09, 1.110359e-09, 1.070212e-09, 1.068826e-09, 
    1.071307e-09, 1.074739e-09, 1.077925e-09, 1.082159e-09, 1.082593e-09, 
    1.083386e-09, 1.085442e-09, 1.08717e-09, 1.083637e-09, 1.087603e-09, 
    1.07272e-09, 1.080519e-09, 1.068303e-09, 1.071981e-09, 1.074537e-09, 
    1.073416e-09, 1.07924e-09, 1.080613e-09, 1.086192e-09, 1.083308e-09, 
    1.100483e-09, 1.092883e-09, 1.113975e-09, 1.10808e-09, 1.068342e-09, 
    1.070207e-09, 1.076698e-09, 1.073609e-09, 1.082442e-09, 1.084617e-09, 
    1.086385e-09, 1.088645e-09, 1.088889e-09, 1.090228e-09, 1.088033e-09, 
    1.090141e-09, 1.082169e-09, 1.085731e-09, 1.075956e-09, 1.078335e-09, 
    1.07724e-09, 1.07604e-09, 1.079745e-09, 1.083692e-09, 1.083777e-09, 
    1.085043e-09, 1.08861e-09, 1.082478e-09, 1.101463e-09, 1.089737e-09, 
    1.072241e-09, 1.075833e-09, 1.076346e-09, 1.074954e-09, 1.084399e-09, 
    1.080976e-09, 1.090195e-09, 1.087703e-09, 1.091786e-09, 1.089757e-09, 
    1.089459e-09, 1.086853e-09, 1.085231e-09, 1.081133e-09, 1.0778e-09, 
    1.075156e-09, 1.075771e-09, 1.078674e-09, 1.083934e-09, 1.088911e-09, 
    1.08782e-09, 1.091476e-09, 1.081802e-09, 1.085858e-09, 1.08429e-09, 
    1.088378e-09, 1.079421e-09, 1.087048e-09, 1.077472e-09, 1.078312e-09, 
    1.080909e-09, 1.086133e-09, 1.087289e-09, 1.088523e-09, 1.087762e-09, 
    1.084068e-09, 1.083463e-09, 1.080845e-09, 1.080123e-09, 1.078129e-09, 
    1.076478e-09, 1.077986e-09, 1.07957e-09, 1.084069e-09, 1.088124e-09, 
    1.092546e-09, 1.093628e-09, 1.098794e-09, 1.094588e-09, 1.101529e-09, 
    1.095627e-09, 1.105844e-09, 1.08749e-09, 1.095454e-09, 1.081027e-09, 
    1.082581e-09, 1.085392e-09, 1.09184e-09, 1.088359e-09, 1.09243e-09, 
    1.083439e-09, 1.078775e-09, 1.077568e-09, 1.075317e-09, 1.07762e-09, 
    1.077432e-09, 1.079636e-09, 1.078928e-09, 1.084219e-09, 1.081377e-09, 
    1.089451e-09, 1.092398e-09, 1.100722e-09, 1.105825e-09, 1.111021e-09, 
    1.113316e-09, 1.114014e-09, 1.114306e-09 ;

 SOIL2C_TO_SOIL3C =
  7.558738e-11, 7.592325e-11, 7.585797e-11, 7.612889e-11, 7.597861e-11, 
    7.615601e-11, 7.565548e-11, 7.593658e-11, 7.575714e-11, 7.561762e-11, 
    7.66547e-11, 7.614098e-11, 7.718853e-11, 7.68608e-11, 7.768417e-11, 
    7.713752e-11, 7.779442e-11, 7.766842e-11, 7.80477e-11, 7.793904e-11, 
    7.842418e-11, 7.809785e-11, 7.867573e-11, 7.834626e-11, 7.839778e-11, 
    7.808709e-11, 7.624437e-11, 7.659074e-11, 7.622385e-11, 7.627324e-11, 
    7.625107e-11, 7.59817e-11, 7.584595e-11, 7.556172e-11, 7.561332e-11, 
    7.582209e-11, 7.629545e-11, 7.613477e-11, 7.653977e-11, 7.653063e-11, 
    7.698158e-11, 7.677825e-11, 7.753632e-11, 7.732085e-11, 7.794358e-11, 
    7.778695e-11, 7.793621e-11, 7.789096e-11, 7.79368e-11, 7.77071e-11, 
    7.780551e-11, 7.76034e-11, 7.681632e-11, 7.70476e-11, 7.635785e-11, 
    7.594317e-11, 7.566781e-11, 7.547241e-11, 7.550003e-11, 7.555269e-11, 
    7.582331e-11, 7.607779e-11, 7.627173e-11, 7.640148e-11, 7.652932e-11, 
    7.691627e-11, 7.712114e-11, 7.757989e-11, 7.749711e-11, 7.763735e-11, 
    7.777137e-11, 7.799635e-11, 7.795933e-11, 7.805845e-11, 7.763367e-11, 
    7.791597e-11, 7.744996e-11, 7.75774e-11, 7.656401e-11, 7.617812e-11, 
    7.601406e-11, 7.587051e-11, 7.552127e-11, 7.576244e-11, 7.566737e-11, 
    7.589357e-11, 7.603732e-11, 7.596623e-11, 7.640502e-11, 7.623442e-11, 
    7.713328e-11, 7.674607e-11, 7.775573e-11, 7.75141e-11, 7.781366e-11, 
    7.76608e-11, 7.792272e-11, 7.7687e-11, 7.809535e-11, 7.818427e-11, 
    7.812351e-11, 7.835695e-11, 7.767393e-11, 7.793621e-11, 7.596423e-11, 
    7.597582e-11, 7.602984e-11, 7.579239e-11, 7.577786e-11, 7.556031e-11, 
    7.57539e-11, 7.583634e-11, 7.604565e-11, 7.616945e-11, 7.628716e-11, 
    7.654596e-11, 7.683502e-11, 7.723928e-11, 7.752977e-11, 7.772449e-11, 
    7.760509e-11, 7.77105e-11, 7.759266e-11, 7.753743e-11, 7.815094e-11, 
    7.780643e-11, 7.832338e-11, 7.829477e-11, 7.806081e-11, 7.829799e-11, 
    7.598396e-11, 7.591724e-11, 7.56856e-11, 7.586688e-11, 7.553661e-11, 
    7.572147e-11, 7.582777e-11, 7.623797e-11, 7.632812e-11, 7.64117e-11, 
    7.657678e-11, 7.678865e-11, 7.716037e-11, 7.748383e-11, 7.777917e-11, 
    7.775753e-11, 7.776515e-11, 7.783112e-11, 7.76677e-11, 7.785795e-11, 
    7.788988e-11, 7.780639e-11, 7.829094e-11, 7.815251e-11, 7.829416e-11, 
    7.820403e-11, 7.593894e-11, 7.60512e-11, 7.599054e-11, 7.610462e-11, 
    7.602424e-11, 7.638163e-11, 7.648879e-11, 7.699029e-11, 7.678448e-11, 
    7.711206e-11, 7.681776e-11, 7.68699e-11, 7.712272e-11, 7.683366e-11, 
    7.746599e-11, 7.703726e-11, 7.783368e-11, 7.740547e-11, 7.786052e-11, 
    7.777789e-11, 7.79147e-11, 7.803724e-11, 7.819141e-11, 7.847588e-11, 
    7.841001e-11, 7.864793e-11, 7.621859e-11, 7.636421e-11, 7.63514e-11, 
    7.650382e-11, 7.661654e-11, 7.686089e-11, 7.725282e-11, 7.710544e-11, 
    7.737604e-11, 7.743036e-11, 7.701926e-11, 7.727165e-11, 7.646168e-11, 
    7.659252e-11, 7.651463e-11, 7.623007e-11, 7.713939e-11, 7.667268e-11, 
    7.753456e-11, 7.728169e-11, 7.801976e-11, 7.765267e-11, 7.837374e-11, 
    7.868202e-11, 7.897225e-11, 7.931138e-11, 7.644371e-11, 7.634475e-11, 
    7.652195e-11, 7.67671e-11, 7.699462e-11, 7.729711e-11, 7.732807e-11, 
    7.738473e-11, 7.753154e-11, 7.765497e-11, 7.740264e-11, 7.768592e-11, 
    7.662285e-11, 7.71799e-11, 7.630733e-11, 7.657004e-11, 7.675265e-11, 
    7.667256e-11, 7.708859e-11, 7.718666e-11, 7.758517e-11, 7.737917e-11, 
    7.860592e-11, 7.80631e-11, 7.956968e-11, 7.914857e-11, 7.631017e-11, 
    7.644337e-11, 7.690697e-11, 7.668638e-11, 7.731731e-11, 7.747263e-11, 
    7.759891e-11, 7.776032e-11, 7.777776e-11, 7.78734e-11, 7.771667e-11, 
    7.786721e-11, 7.729775e-11, 7.755221e-11, 7.685399e-11, 7.702391e-11, 
    7.694574e-11, 7.686e-11, 7.712465e-11, 7.740661e-11, 7.741265e-11, 
    7.750307e-11, 7.775783e-11, 7.731987e-11, 7.867595e-11, 7.783837e-11, 
    7.658862e-11, 7.684518e-11, 7.688185e-11, 7.678246e-11, 7.745705e-11, 
    7.72126e-11, 7.787106e-11, 7.76931e-11, 7.798471e-11, 7.78398e-11, 
    7.781847e-11, 7.763237e-11, 7.751651e-11, 7.722381e-11, 7.698568e-11, 
    7.679688e-11, 7.684078e-11, 7.704818e-11, 7.742387e-11, 7.777932e-11, 
    7.770146e-11, 7.796255e-11, 7.727156e-11, 7.756127e-11, 7.744929e-11, 
    7.774129e-11, 7.710152e-11, 7.764626e-11, 7.696229e-11, 7.702226e-11, 
    7.720775e-11, 7.758091e-11, 7.76635e-11, 7.775166e-11, 7.769727e-11, 
    7.743341e-11, 7.739018e-11, 7.720324e-11, 7.715163e-11, 7.70092e-11, 
    7.689129e-11, 7.699901e-11, 7.711216e-11, 7.743352e-11, 7.772316e-11, 
    7.803897e-11, 7.811628e-11, 7.848529e-11, 7.818488e-11, 7.868062e-11, 
    7.825911e-11, 7.898883e-11, 7.767786e-11, 7.824674e-11, 7.72162e-11, 
    7.732721e-11, 7.752798e-11, 7.798857e-11, 7.773993e-11, 7.803072e-11, 
    7.738849e-11, 7.705533e-11, 7.696915e-11, 7.680835e-11, 7.697283e-11, 
    7.695945e-11, 7.711685e-11, 7.706627e-11, 7.74442e-11, 7.724119e-11, 
    7.781794e-11, 7.802843e-11, 7.862299e-11, 7.898752e-11, 7.935867e-11, 
    7.952254e-11, 7.957242e-11, 7.959327e-11 ;

 SOIL2C_vr =
  20.00596, 20.00598, 20.00597, 20.00599, 20.00598, 20.00599, 20.00596, 
    20.00598, 20.00597, 20.00596, 20.00601, 20.00599, 20.00604, 20.00602, 
    20.00606, 20.00603, 20.00607, 20.00606, 20.00608, 20.00607, 20.0061, 
    20.00608, 20.00611, 20.00609, 20.00609, 20.00608, 20.00599, 20.00601, 
    20.00599, 20.00599, 20.00599, 20.00598, 20.00597, 20.00596, 20.00596, 
    20.00597, 20.00599, 20.00599, 20.006, 20.006, 20.00603, 20.00602, 
    20.00605, 20.00604, 20.00607, 20.00607, 20.00607, 20.00607, 20.00607, 
    20.00606, 20.00607, 20.00606, 20.00602, 20.00603, 20.006, 20.00598, 
    20.00596, 20.00595, 20.00595, 20.00596, 20.00597, 20.00598, 20.00599, 
    20.006, 20.006, 20.00602, 20.00603, 20.00606, 20.00605, 20.00606, 
    20.00607, 20.00607, 20.00607, 20.00608, 20.00606, 20.00607, 20.00605, 
    20.00606, 20.00601, 20.00599, 20.00598, 20.00597, 20.00595, 20.00597, 
    20.00596, 20.00597, 20.00598, 20.00598, 20.006, 20.00599, 20.00603, 
    20.00602, 20.00606, 20.00605, 20.00607, 20.00606, 20.00607, 20.00606, 
    20.00608, 20.00608, 20.00608, 20.00609, 20.00606, 20.00607, 20.00598, 
    20.00598, 20.00598, 20.00597, 20.00597, 20.00596, 20.00597, 20.00597, 
    20.00598, 20.00599, 20.00599, 20.00601, 20.00602, 20.00604, 20.00605, 
    20.00606, 20.00606, 20.00606, 20.00606, 20.00605, 20.00608, 20.00607, 
    20.00609, 20.00609, 20.00608, 20.00609, 20.00598, 20.00598, 20.00596, 
    20.00597, 20.00596, 20.00597, 20.00597, 20.00599, 20.00599, 20.006, 
    20.00601, 20.00602, 20.00603, 20.00605, 20.00607, 20.00606, 20.00606, 
    20.00607, 20.00606, 20.00607, 20.00607, 20.00607, 20.00609, 20.00608, 
    20.00609, 20.00608, 20.00598, 20.00598, 20.00598, 20.00598, 20.00598, 
    20.006, 20.006, 20.00603, 20.00602, 20.00603, 20.00602, 20.00602, 
    20.00603, 20.00602, 20.00605, 20.00603, 20.00607, 20.00605, 20.00607, 
    20.00607, 20.00607, 20.00608, 20.00608, 20.0061, 20.0061, 20.00611, 
    20.00599, 20.006, 20.006, 20.006, 20.00601, 20.00602, 20.00604, 20.00603, 
    20.00605, 20.00605, 20.00603, 20.00604, 20.006, 20.00601, 20.006, 
    20.00599, 20.00603, 20.00601, 20.00605, 20.00604, 20.00608, 20.00606, 
    20.00609, 20.00611, 20.00612, 20.00614, 20.006, 20.00599, 20.006, 
    20.00602, 20.00603, 20.00604, 20.00604, 20.00605, 20.00605, 20.00606, 
    20.00605, 20.00606, 20.00601, 20.00604, 20.00599, 20.00601, 20.00602, 
    20.00601, 20.00603, 20.00604, 20.00606, 20.00605, 20.00611, 20.00608, 
    20.00615, 20.00613, 20.00599, 20.006, 20.00602, 20.00601, 20.00604, 
    20.00605, 20.00606, 20.00606, 20.00607, 20.00607, 20.00606, 20.00607, 
    20.00604, 20.00605, 20.00602, 20.00603, 20.00603, 20.00602, 20.00603, 
    20.00605, 20.00605, 20.00605, 20.00606, 20.00604, 20.00611, 20.00607, 
    20.00601, 20.00602, 20.00602, 20.00602, 20.00605, 20.00604, 20.00607, 
    20.00606, 20.00607, 20.00607, 20.00607, 20.00606, 20.00605, 20.00604, 
    20.00603, 20.00602, 20.00602, 20.00603, 20.00605, 20.00607, 20.00606, 
    20.00607, 20.00604, 20.00605, 20.00605, 20.00606, 20.00603, 20.00606, 
    20.00603, 20.00603, 20.00604, 20.00606, 20.00606, 20.00606, 20.00606, 
    20.00605, 20.00605, 20.00604, 20.00603, 20.00603, 20.00602, 20.00603, 
    20.00603, 20.00605, 20.00606, 20.00608, 20.00608, 20.0061, 20.00608, 
    20.00611, 20.00609, 20.00612, 20.00606, 20.00609, 20.00604, 20.00604, 
    20.00605, 20.00607, 20.00606, 20.00608, 20.00605, 20.00603, 20.00603, 
    20.00602, 20.00603, 20.00603, 20.00603, 20.00603, 20.00605, 20.00604, 
    20.00607, 20.00608, 20.00611, 20.00612, 20.00614, 20.00615, 20.00615, 
    20.00615,
  20.00537, 20.0054, 20.00539, 20.00541, 20.0054, 20.00541, 20.00538, 
    20.0054, 20.00538, 20.00538, 20.00544, 20.00541, 20.00547, 20.00545, 
    20.0055, 20.00547, 20.00551, 20.0055, 20.00553, 20.00552, 20.00555, 
    20.00553, 20.00556, 20.00554, 20.00555, 20.00553, 20.00541, 20.00544, 
    20.00541, 20.00542, 20.00541, 20.0054, 20.00539, 20.00537, 20.00538, 
    20.00539, 20.00542, 20.00541, 20.00543, 20.00543, 20.00546, 20.00545, 
    20.00549, 20.00548, 20.00552, 20.00551, 20.00552, 20.00552, 20.00552, 
    20.0055, 20.00551, 20.0055, 20.00545, 20.00546, 20.00542, 20.0054, 
    20.00538, 20.00537, 20.00537, 20.00537, 20.00539, 20.00541, 20.00542, 
    20.00542, 20.00543, 20.00546, 20.00547, 20.0055, 20.00549, 20.0055, 
    20.00551, 20.00552, 20.00552, 20.00553, 20.0055, 20.00552, 20.00549, 
    20.0055, 20.00543, 20.00541, 20.0054, 20.00539, 20.00537, 20.00539, 
    20.00538, 20.00539, 20.0054, 20.0054, 20.00542, 20.00541, 20.00547, 
    20.00545, 20.00551, 20.00549, 20.00551, 20.0055, 20.00552, 20.0055, 
    20.00553, 20.00553, 20.00553, 20.00554, 20.0055, 20.00552, 20.0054, 
    20.0054, 20.0054, 20.00539, 20.00539, 20.00537, 20.00538, 20.00539, 
    20.0054, 20.00541, 20.00542, 20.00543, 20.00545, 20.00548, 20.00549, 
    20.0055, 20.0055, 20.0055, 20.0055, 20.00549, 20.00553, 20.00551, 
    20.00554, 20.00554, 20.00553, 20.00554, 20.0054, 20.0054, 20.00538, 
    20.00539, 20.00537, 20.00538, 20.00539, 20.00541, 20.00542, 20.00542, 
    20.00544, 20.00545, 20.00547, 20.00549, 20.00551, 20.00551, 20.00551, 
    20.00551, 20.0055, 20.00551, 20.00552, 20.00551, 20.00554, 20.00553, 
    20.00554, 20.00554, 20.0054, 20.0054, 20.0054, 20.00541, 20.0054, 
    20.00542, 20.00543, 20.00546, 20.00545, 20.00547, 20.00545, 20.00545, 
    20.00547, 20.00545, 20.00549, 20.00546, 20.00551, 20.00549, 20.00551, 
    20.00551, 20.00552, 20.00552, 20.00553, 20.00555, 20.00555, 20.00556, 
    20.00541, 20.00542, 20.00542, 20.00543, 20.00544, 20.00545, 20.00548, 
    20.00547, 20.00548, 20.00549, 20.00546, 20.00548, 20.00543, 20.00544, 
    20.00543, 20.00541, 20.00547, 20.00544, 20.00549, 20.00548, 20.00552, 
    20.0055, 20.00554, 20.00556, 20.00558, 20.0056, 20.00543, 20.00542, 
    20.00543, 20.00545, 20.00546, 20.00548, 20.00548, 20.00549, 20.00549, 
    20.0055, 20.00549, 20.0055, 20.00544, 20.00547, 20.00542, 20.00544, 
    20.00545, 20.00544, 20.00547, 20.00547, 20.0055, 20.00548, 20.00556, 
    20.00553, 20.00562, 20.00559, 20.00542, 20.00543, 20.00546, 20.00544, 
    20.00548, 20.00549, 20.0055, 20.00551, 20.00551, 20.00551, 20.0055, 
    20.00551, 20.00548, 20.0055, 20.00545, 20.00546, 20.00546, 20.00545, 
    20.00547, 20.00549, 20.00549, 20.00549, 20.00551, 20.00548, 20.00556, 
    20.00551, 20.00544, 20.00545, 20.00545, 20.00545, 20.00549, 20.00547, 
    20.00551, 20.0055, 20.00552, 20.00551, 20.00551, 20.0055, 20.00549, 
    20.00547, 20.00546, 20.00545, 20.00545, 20.00546, 20.00549, 20.00551, 
    20.0055, 20.00552, 20.00548, 20.0055, 20.00549, 20.00551, 20.00547, 
    20.0055, 20.00546, 20.00546, 20.00547, 20.0055, 20.0055, 20.00551, 
    20.0055, 20.00549, 20.00549, 20.00547, 20.00547, 20.00546, 20.00546, 
    20.00546, 20.00547, 20.00549, 20.0055, 20.00552, 20.00553, 20.00555, 
    20.00553, 20.00556, 20.00554, 20.00558, 20.0055, 20.00554, 20.00547, 
    20.00548, 20.00549, 20.00552, 20.00551, 20.00552, 20.00549, 20.00546, 
    20.00546, 20.00545, 20.00546, 20.00546, 20.00547, 20.00546, 20.00549, 
    20.00548, 20.00551, 20.00552, 20.00556, 20.00558, 20.0056, 20.00562, 
    20.00562, 20.00562,
  20.00504, 20.00507, 20.00506, 20.00508, 20.00507, 20.00508, 20.00505, 
    20.00507, 20.00506, 20.00505, 20.00512, 20.00508, 20.00515, 20.00513, 
    20.00518, 20.00515, 20.00519, 20.00518, 20.00521, 20.0052, 20.00523, 
    20.00521, 20.00525, 20.00523, 20.00523, 20.00521, 20.00509, 20.00511, 
    20.00509, 20.00509, 20.00509, 20.00507, 20.00506, 20.00504, 20.00505, 
    20.00506, 20.00509, 20.00508, 20.00511, 20.00511, 20.00514, 20.00513, 
    20.00517, 20.00516, 20.0052, 20.00519, 20.0052, 20.0052, 20.0052, 
    20.00519, 20.00519, 20.00518, 20.00513, 20.00514, 20.0051, 20.00507, 
    20.00505, 20.00504, 20.00504, 20.00504, 20.00506, 20.00508, 20.00509, 
    20.0051, 20.00511, 20.00513, 20.00515, 20.00518, 20.00517, 20.00518, 
    20.00519, 20.00521, 20.0052, 20.00521, 20.00518, 20.0052, 20.00517, 
    20.00518, 20.00511, 20.00508, 20.00507, 20.00506, 20.00504, 20.00506, 
    20.00505, 20.00507, 20.00508, 20.00507, 20.0051, 20.00509, 20.00515, 
    20.00512, 20.00519, 20.00517, 20.00519, 20.00518, 20.0052, 20.00519, 
    20.00521, 20.00522, 20.00521, 20.00523, 20.00518, 20.0052, 20.00507, 
    20.00507, 20.00507, 20.00506, 20.00506, 20.00504, 20.00506, 20.00506, 
    20.00508, 20.00508, 20.00509, 20.00511, 20.00513, 20.00516, 20.00517, 
    20.00519, 20.00518, 20.00519, 20.00518, 20.00517, 20.00522, 20.00519, 
    20.00523, 20.00523, 20.00521, 20.00523, 20.00507, 20.00507, 20.00505, 
    20.00506, 20.00504, 20.00505, 20.00506, 20.00509, 20.00509, 20.0051, 
    20.00511, 20.00513, 20.00515, 20.00517, 20.00519, 20.00519, 20.00519, 
    20.0052, 20.00518, 20.0052, 20.0052, 20.00519, 20.00523, 20.00522, 
    20.00523, 20.00522, 20.00507, 20.00508, 20.00507, 20.00508, 20.00507, 
    20.0051, 20.00511, 20.00514, 20.00513, 20.00515, 20.00513, 20.00513, 
    20.00515, 20.00513, 20.00517, 20.00514, 20.0052, 20.00517, 20.0052, 
    20.00519, 20.0052, 20.00521, 20.00522, 20.00524, 20.00523, 20.00525, 
    20.00509, 20.0051, 20.0051, 20.00511, 20.00511, 20.00513, 20.00516, 
    20.00515, 20.00517, 20.00517, 20.00514, 20.00516, 20.0051, 20.00511, 
    20.00511, 20.00509, 20.00515, 20.00512, 20.00517, 20.00516, 20.00521, 
    20.00518, 20.00523, 20.00525, 20.00527, 20.00529, 20.0051, 20.0051, 
    20.00511, 20.00512, 20.00514, 20.00516, 20.00516, 20.00517, 20.00517, 
    20.00518, 20.00517, 20.00518, 20.00511, 20.00515, 20.00509, 20.00511, 
    20.00512, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 20.00525, 
    20.00521, 20.00531, 20.00528, 20.00509, 20.0051, 20.00513, 20.00512, 
    20.00516, 20.00517, 20.00518, 20.00519, 20.00519, 20.0052, 20.00519, 
    20.0052, 20.00516, 20.00518, 20.00513, 20.00514, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00517, 20.00517, 20.00519, 20.00516, 20.00525, 
    20.0052, 20.00511, 20.00513, 20.00513, 20.00513, 20.00517, 20.00515, 
    20.0052, 20.00519, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00515, 20.00514, 20.00513, 20.00513, 20.00514, 20.00517, 20.00519, 
    20.00519, 20.0052, 20.00516, 20.00518, 20.00517, 20.00519, 20.00515, 
    20.00518, 20.00514, 20.00514, 20.00515, 20.00518, 20.00518, 20.00519, 
    20.00519, 20.00517, 20.00517, 20.00515, 20.00515, 20.00514, 20.00513, 
    20.00514, 20.00515, 20.00517, 20.00519, 20.00521, 20.00521, 20.00524, 
    20.00522, 20.00525, 20.00522, 20.00527, 20.00518, 20.00522, 20.00515, 
    20.00516, 20.00517, 20.00521, 20.00519, 20.00521, 20.00517, 20.00514, 
    20.00514, 20.00513, 20.00514, 20.00514, 20.00515, 20.00514, 20.00517, 
    20.00516, 20.00519, 20.00521, 20.00525, 20.00527, 20.0053, 20.00531, 
    20.00531, 20.00531,
  20.00479, 20.00481, 20.00481, 20.00483, 20.00482, 20.00483, 20.0048, 
    20.00481, 20.0048, 20.00479, 20.00486, 20.00483, 20.0049, 20.00488, 
    20.00493, 20.0049, 20.00494, 20.00493, 20.00496, 20.00495, 20.00498, 
    20.00496, 20.005, 20.00498, 20.00498, 20.00496, 20.00484, 20.00486, 
    20.00484, 20.00484, 20.00484, 20.00482, 20.00481, 20.00479, 20.00479, 
    20.00481, 20.00484, 20.00483, 20.00486, 20.00486, 20.00489, 20.00487, 
    20.00492, 20.00491, 20.00495, 20.00494, 20.00495, 20.00495, 20.00495, 
    20.00494, 20.00494, 20.00493, 20.00488, 20.00489, 20.00484, 20.00482, 
    20.0048, 20.00478, 20.00479, 20.00479, 20.00481, 20.00482, 20.00484, 
    20.00485, 20.00485, 20.00488, 20.0049, 20.00493, 20.00492, 20.00493, 
    20.00494, 20.00496, 20.00495, 20.00496, 20.00493, 20.00495, 20.00492, 
    20.00493, 20.00486, 20.00483, 20.00482, 20.00481, 20.00479, 20.0048, 
    20.0048, 20.00481, 20.00482, 20.00482, 20.00485, 20.00484, 20.0049, 
    20.00487, 20.00494, 20.00492, 20.00494, 20.00493, 20.00495, 20.00493, 
    20.00496, 20.00497, 20.00496, 20.00498, 20.00493, 20.00495, 20.00482, 
    20.00482, 20.00482, 20.0048, 20.0048, 20.00479, 20.0048, 20.00481, 
    20.00482, 20.00483, 20.00484, 20.00486, 20.00488, 20.0049, 20.00492, 
    20.00494, 20.00493, 20.00494, 20.00493, 20.00492, 20.00496, 20.00494, 
    20.00498, 20.00497, 20.00496, 20.00498, 20.00482, 20.00481, 20.0048, 
    20.00481, 20.00479, 20.0048, 20.00481, 20.00484, 20.00484, 20.00485, 
    20.00486, 20.00487, 20.0049, 20.00492, 20.00494, 20.00494, 20.00494, 
    20.00494, 20.00493, 20.00495, 20.00495, 20.00494, 20.00497, 20.00496, 
    20.00497, 20.00497, 20.00481, 20.00482, 20.00482, 20.00483, 20.00482, 
    20.00484, 20.00485, 20.00489, 20.00487, 20.00489, 20.00488, 20.00488, 
    20.0049, 20.00488, 20.00492, 20.00489, 20.00494, 20.00492, 20.00495, 
    20.00494, 20.00495, 20.00496, 20.00497, 20.00499, 20.00498, 20.005, 
    20.00483, 20.00484, 20.00484, 20.00485, 20.00486, 20.00488, 20.0049, 
    20.00489, 20.00491, 20.00492, 20.00489, 20.00491, 20.00485, 20.00486, 
    20.00485, 20.00484, 20.0049, 20.00487, 20.00492, 20.00491, 20.00496, 
    20.00493, 20.00498, 20.005, 20.00502, 20.00504, 20.00485, 20.00484, 
    20.00485, 20.00487, 20.00489, 20.00491, 20.00491, 20.00491, 20.00492, 
    20.00493, 20.00492, 20.00493, 20.00486, 20.0049, 20.00484, 20.00486, 
    20.00487, 20.00487, 20.00489, 20.0049, 20.00493, 20.00491, 20.005, 
    20.00496, 20.00506, 20.00503, 20.00484, 20.00485, 20.00488, 20.00487, 
    20.00491, 20.00492, 20.00493, 20.00494, 20.00494, 20.00495, 20.00494, 
    20.00495, 20.00491, 20.00492, 20.00488, 20.00489, 20.00488, 20.00488, 
    20.0049, 20.00492, 20.00492, 20.00492, 20.00494, 20.00491, 20.005, 
    20.00494, 20.00486, 20.00488, 20.00488, 20.00487, 20.00492, 20.0049, 
    20.00495, 20.00493, 20.00495, 20.00494, 20.00494, 20.00493, 20.00492, 
    20.0049, 20.00489, 20.00487, 20.00488, 20.00489, 20.00492, 20.00494, 
    20.00493, 20.00495, 20.00491, 20.00492, 20.00492, 20.00494, 20.00489, 
    20.00493, 20.00488, 20.00489, 20.0049, 20.00493, 20.00493, 20.00494, 
    20.00493, 20.00492, 20.00491, 20.0049, 20.0049, 20.00489, 20.00488, 
    20.00489, 20.00489, 20.00492, 20.00494, 20.00496, 20.00496, 20.00499, 
    20.00497, 20.005, 20.00497, 20.00502, 20.00493, 20.00497, 20.0049, 
    20.00491, 20.00492, 20.00496, 20.00494, 20.00496, 20.00491, 20.00489, 
    20.00488, 20.00487, 20.00488, 20.00488, 20.00489, 20.00489, 20.00492, 
    20.0049, 20.00494, 20.00496, 20.005, 20.00502, 20.00505, 20.00506, 
    20.00506, 20.00506,
  20.00425, 20.00427, 20.00427, 20.00428, 20.00427, 20.00428, 20.00425, 
    20.00427, 20.00426, 20.00425, 20.00431, 20.00428, 20.00434, 20.00433, 
    20.00437, 20.00434, 20.00438, 20.00437, 20.0044, 20.00439, 20.00442, 
    20.0044, 20.00443, 20.00441, 20.00442, 20.0044, 20.00429, 20.00431, 
    20.00429, 20.00429, 20.00429, 20.00427, 20.00426, 20.00425, 20.00425, 
    20.00426, 20.00429, 20.00428, 20.00431, 20.00431, 20.00433, 20.00432, 
    20.00437, 20.00435, 20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 
    20.00438, 20.00438, 20.00437, 20.00432, 20.00434, 20.0043, 20.00427, 
    20.00426, 20.00424, 20.00424, 20.00425, 20.00426, 20.00428, 20.00429, 
    20.0043, 20.00431, 20.00433, 20.00434, 20.00437, 20.00436, 20.00437, 
    20.00438, 20.00439, 20.00439, 20.0044, 20.00437, 20.00439, 20.00436, 
    20.00437, 20.00431, 20.00429, 20.00427, 20.00427, 20.00425, 20.00426, 
    20.00426, 20.00427, 20.00428, 20.00427, 20.0043, 20.00429, 20.00434, 
    20.00432, 20.00438, 20.00436, 20.00438, 20.00437, 20.00439, 20.00438, 
    20.0044, 20.0044, 20.0044, 20.00441, 20.00437, 20.00439, 20.00427, 
    20.00427, 20.00428, 20.00426, 20.00426, 20.00425, 20.00426, 20.00426, 
    20.00428, 20.00428, 20.00429, 20.00431, 20.00432, 20.00435, 20.00437, 
    20.00438, 20.00437, 20.00438, 20.00437, 20.00437, 20.0044, 20.00438, 
    20.00441, 20.00441, 20.0044, 20.00441, 20.00427, 20.00427, 20.00426, 
    20.00427, 20.00425, 20.00426, 20.00426, 20.00429, 20.00429, 20.0043, 
    20.00431, 20.00432, 20.00434, 20.00436, 20.00438, 20.00438, 20.00438, 
    20.00438, 20.00437, 20.00438, 20.00439, 20.00438, 20.00441, 20.0044, 
    20.00441, 20.00441, 20.00427, 20.00428, 20.00427, 20.00428, 20.00428, 
    20.0043, 20.0043, 20.00433, 20.00432, 20.00434, 20.00432, 20.00433, 
    20.00434, 20.00432, 20.00436, 20.00434, 20.00438, 20.00436, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.0044, 20.00442, 20.00442, 20.00443, 
    20.00429, 20.0043, 20.0043, 20.0043, 20.00431, 20.00433, 20.00435, 
    20.00434, 20.00436, 20.00436, 20.00434, 20.00435, 20.0043, 20.00431, 
    20.0043, 20.00429, 20.00434, 20.00431, 20.00437, 20.00435, 20.00439, 
    20.00437, 20.00442, 20.00443, 20.00445, 20.00447, 20.0043, 20.0043, 
    20.0043, 20.00432, 20.00433, 20.00435, 20.00435, 20.00436, 20.00437, 
    20.00437, 20.00436, 20.00438, 20.00431, 20.00434, 20.00429, 20.00431, 
    20.00432, 20.00431, 20.00434, 20.00434, 20.00437, 20.00436, 20.00443, 
    20.0044, 20.00449, 20.00446, 20.00429, 20.0043, 20.00433, 20.00431, 
    20.00435, 20.00436, 20.00437, 20.00438, 20.00438, 20.00438, 20.00438, 
    20.00438, 20.00435, 20.00437, 20.00433, 20.00434, 20.00433, 20.00433, 
    20.00434, 20.00436, 20.00436, 20.00436, 20.00438, 20.00435, 20.00443, 
    20.00438, 20.00431, 20.00432, 20.00433, 20.00432, 20.00436, 20.00435, 
    20.00438, 20.00438, 20.00439, 20.00438, 20.00438, 20.00437, 20.00436, 
    20.00435, 20.00433, 20.00432, 20.00432, 20.00434, 20.00436, 20.00438, 
    20.00438, 20.00439, 20.00435, 20.00437, 20.00436, 20.00438, 20.00434, 
    20.00437, 20.00433, 20.00434, 20.00435, 20.00437, 20.00437, 20.00438, 
    20.00438, 20.00436, 20.00436, 20.00434, 20.00434, 20.00433, 20.00433, 
    20.00433, 20.00434, 20.00436, 20.00438, 20.0044, 20.0044, 20.00442, 
    20.0044, 20.00443, 20.00441, 20.00445, 20.00437, 20.00441, 20.00435, 
    20.00435, 20.00437, 20.00439, 20.00438, 20.00439, 20.00436, 20.00434, 
    20.00433, 20.00432, 20.00433, 20.00433, 20.00434, 20.00434, 20.00436, 
    20.00435, 20.00438, 20.00439, 20.00443, 20.00445, 20.00447, 20.00448, 
    20.00449, 20.00449,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258144, 0.525815, 0.5258148, 0.5258153, 0.525815, 0.5258153, 0.5258145, 
    0.525815, 0.5258147, 0.5258145, 0.5258161, 0.5258153, 0.525817, 
    0.5258165, 0.5258178, 0.5258169, 0.525818, 0.5258178, 0.5258184, 
    0.5258182, 0.5258191, 0.5258185, 0.5258195, 0.5258189, 0.525819, 
    0.5258185, 0.5258155, 0.525816, 0.5258154, 0.5258155, 0.5258155, 
    0.5258151, 0.5258148, 0.5258144, 0.5258144, 0.5258148, 0.5258155, 
    0.5258153, 0.525816, 0.525816, 0.5258167, 0.5258163, 0.5258176, 
    0.5258172, 0.5258182, 0.525818, 0.5258182, 0.5258182, 0.5258182, 
    0.5258179, 0.525818, 0.5258177, 0.5258164, 0.5258168, 0.5258157, 
    0.525815, 0.5258145, 0.5258142, 0.5258142, 0.5258144, 0.5258148, 
    0.5258152, 0.5258155, 0.5258157, 0.525816, 0.5258166, 0.5258169, 
    0.5258176, 0.5258175, 0.5258178, 0.525818, 0.5258183, 0.5258183, 
    0.5258185, 0.5258178, 0.5258182, 0.5258175, 0.5258176, 0.525816, 
    0.5258154, 0.5258151, 0.5258149, 0.5258143, 0.5258147, 0.5258145, 
    0.5258149, 0.5258151, 0.525815, 0.5258157, 0.5258155, 0.5258169, 
    0.5258163, 0.5258179, 0.5258176, 0.525818, 0.5258178, 0.5258182, 
    0.5258178, 0.5258185, 0.5258186, 0.5258185, 0.5258189, 0.5258178, 
    0.5258182, 0.525815, 0.525815, 0.5258151, 0.5258147, 0.5258147, 
    0.5258144, 0.5258147, 0.5258148, 0.5258151, 0.5258154, 0.5258155, 
    0.525816, 0.5258164, 0.5258171, 0.5258176, 0.5258179, 0.5258177, 
    0.5258179, 0.5258177, 0.5258176, 0.5258186, 0.525818, 0.5258189, 
    0.5258188, 0.5258185, 0.5258188, 0.5258151, 0.525815, 0.5258145, 
    0.5258148, 0.5258143, 0.5258146, 0.5258148, 0.5258155, 0.5258156, 
    0.5258157, 0.525816, 0.5258164, 0.525817, 0.5258175, 0.525818, 0.5258179, 
    0.525818, 0.525818, 0.5258178, 0.5258181, 0.5258182, 0.525818, 0.5258188, 
    0.5258186, 0.5258188, 0.5258187, 0.525815, 0.5258151, 0.5258151, 
    0.5258152, 0.5258151, 0.5258157, 0.5258158, 0.5258167, 0.5258164, 
    0.5258169, 0.5258164, 0.5258165, 0.5258169, 0.5258164, 0.5258175, 
    0.5258168, 0.525818, 0.5258174, 0.5258181, 0.525818, 0.5258182, 
    0.5258184, 0.5258186, 0.5258191, 0.525819, 0.5258194, 0.5258154, 
    0.5258157, 0.5258157, 0.5258159, 0.5258161, 0.5258165, 0.5258171, 
    0.5258169, 0.5258173, 0.5258174, 0.5258167, 0.5258172, 0.5258158, 
    0.525816, 0.5258159, 0.5258154, 0.5258169, 0.5258162, 0.5258176, 
    0.5258172, 0.5258184, 0.5258178, 0.5258189, 0.5258195, 0.52582, 
    0.5258205, 0.5258158, 0.5258157, 0.5258159, 0.5258163, 0.5258167, 
    0.5258172, 0.5258173, 0.5258173, 0.5258176, 0.5258178, 0.5258174, 
    0.5258178, 0.5258161, 0.525817, 0.5258156, 0.525816, 0.5258163, 
    0.5258162, 0.5258169, 0.525817, 0.5258177, 0.5258173, 0.5258194, 
    0.5258185, 0.5258209, 0.5258203, 0.5258156, 0.5258158, 0.5258166, 
    0.5258162, 0.5258172, 0.5258175, 0.5258177, 0.5258179, 0.525818, 
    0.5258182, 0.5258179, 0.5258181, 0.5258172, 0.5258176, 0.5258165, 
    0.5258167, 0.5258166, 0.5258165, 0.5258169, 0.5258174, 0.5258174, 
    0.5258175, 0.5258179, 0.5258172, 0.5258195, 0.5258181, 0.525816, 
    0.5258164, 0.5258165, 0.5258164, 0.5258175, 0.525817, 0.5258181, 
    0.5258179, 0.5258183, 0.5258181, 0.525818, 0.5258178, 0.5258176, 
    0.5258171, 0.5258167, 0.5258164, 0.5258164, 0.5258168, 0.5258174, 
    0.525818, 0.5258179, 0.5258183, 0.5258172, 0.5258176, 0.5258175, 
    0.5258179, 0.5258169, 0.5258178, 0.5258167, 0.5258167, 0.525817, 
    0.5258176, 0.5258178, 0.5258179, 0.5258179, 0.5258174, 0.5258173, 
    0.525817, 0.525817, 0.5258167, 0.5258166, 0.5258167, 0.5258169, 
    0.5258174, 0.5258179, 0.5258184, 0.5258185, 0.5258191, 0.5258186, 
    0.5258195, 0.5258188, 0.52582, 0.5258178, 0.5258188, 0.525817, 0.5258173, 
    0.5258176, 0.5258183, 0.5258179, 0.5258184, 0.5258173, 0.5258168, 
    0.5258167, 0.5258164, 0.5258167, 0.5258166, 0.5258169, 0.5258168, 
    0.5258175, 0.5258171, 0.525818, 0.5258184, 0.5258194, 0.52582, 0.5258206, 
    0.5258209, 0.5258209, 0.525821 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -7.709882e-21, 7.709882e-21, 1.541976e-20, 1.003089e-36, 2.569961e-21, 
    -1.003089e-36, 2.312965e-20, -5.139921e-21, 1.28498e-20, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    1.027984e-20, -7.709882e-21, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, -2.569961e-21, 0, -1.28498e-20, 
    1.003089e-36, 1.027984e-20, 1.027984e-20, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 5.139921e-21, 1.003089e-36, 2.569961e-21, 
    -7.709882e-21, 1.003089e-36, 5.139921e-21, -2.569961e-21, -1.003089e-36, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, -1.027984e-20, 2.826957e-20, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 1.027984e-20, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, 1.798972e-20, 1.541976e-20, -2.569961e-21, 
    5.139921e-21, -2.055969e-20, -1.28498e-20, 1.28498e-20, -1.28498e-20, 
    -2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -3.083953e-20, -1.027984e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    -1.027984e-20, -1.798972e-20, 7.709882e-21, -2.569961e-21, -7.709882e-21, 
    1.541976e-20, 5.139921e-21, 1.28498e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -1.027984e-20, 0, -2.569961e-21, -1.003089e-36, 
    1.28498e-20, 5.139921e-21, 1.003089e-36, -1.027984e-20, -2.569961e-21, 
    -1.28498e-20, -2.312965e-20, -1.798972e-20, 5.139921e-21, 1.003089e-36, 
    2.569961e-21, 1.003089e-36, -1.027984e-20, -7.709882e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, -2.055969e-20, 
    1.541976e-20, -7.709882e-21, 5.139921e-21, 1.28498e-20, 1.541976e-20, 
    -7.709882e-21, -1.28498e-20, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -1.027984e-20, -3.083953e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -1.798972e-20, 0, 2.569961e-21, -2.569961e-21, -1.28498e-20, 
    1.003089e-36, -1.541976e-20, -1.798972e-20, -1.28498e-20, -1.027984e-20, 
    5.139921e-21, 1.541976e-20, 7.709882e-21, 2.569961e-21, -1.027984e-20, 0, 
    1.027984e-20, -7.709882e-21, -5.139921e-21, -1.541976e-20, -1.798972e-20, 
    7.709882e-21, 1.28498e-20, 1.798972e-20, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, -2.055969e-20, 1.28498e-20, 
    -5.139921e-21, -2.312965e-20, -1.28498e-20, -2.569961e-21, -1.798972e-20, 
    -7.709882e-21, 1.541976e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, -1.003089e-36, 1.541976e-20, 2.569961e-21, -1.541976e-20, 
    1.003089e-36, 5.139921e-21, -7.709882e-21, 1.541976e-20, 1.541976e-20, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 2.569961e-20, 
    5.139921e-21, 1.798972e-20, 2.569961e-21, 1.798972e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, -2.312965e-20, -2.055969e-20, 1.28498e-20, 
    1.003089e-36, -2.569961e-21, -2.312965e-20, 2.569961e-21, 1.003089e-36, 
    1.28498e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -2.312965e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 2.055969e-20, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -2.055969e-20, 2.569961e-20, 2.569961e-21, 
    0, 2.826957e-20, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 2.312965e-20, 2.569961e-21, -7.709882e-21, 
    -1.28498e-20, -7.709882e-21, 2.569961e-21, -7.709882e-21, 1.28498e-20, 
    -2.569961e-21, -1.541976e-20, -2.569961e-21, 1.28498e-20, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, -2.569961e-21, 1.003089e-36, -5.139921e-21, 
    1.003089e-36, -1.28498e-20, -1.027984e-20, 2.055969e-20, -1.28498e-20, 
    -2.055969e-20, 1.28498e-20, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    1.003089e-36, 1.28498e-20, -1.541976e-20, 0, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.541976e-20, -7.709882e-21, 7.709882e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 1.027984e-20, 1.28498e-20, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, -5.139921e-21, 2.055969e-20, -2.312965e-20, 
    7.709882e-21, 1.541976e-20, 7.709882e-21, -5.139921e-21, -1.003089e-36, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    1.541976e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, -2.569961e-21, 
    0, 1.003089e-36, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, -5.139921e-21,
  -5.139921e-21, 7.709882e-21, 1.28498e-20, -2.569961e-21, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, 7.709882e-21, 1.28498e-20, -1.541976e-20, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, 0, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, -1.003089e-36, -7.709882e-21, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, 7.709882e-21, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, 2.569961e-21, -7.709882e-21, 
    1.003089e-36, 2.569961e-21, -5.139921e-21, -1.027984e-20, -1.003089e-36, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    7.709882e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -1.28498e-20, 0, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, -1.003089e-36, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 2.055969e-20, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 0, 2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, 1.003089e-36, 1.28498e-20, 
    -2.569961e-21, 1.027984e-20, -7.709882e-21, -1.027984e-20, 0, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    0, 2.569961e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -1.28498e-20, -7.709882e-21, -2.569961e-21, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 
    1.28498e-20, -1.027984e-20, -7.709882e-21, -7.709882e-21, 0, 0, 
    5.139921e-21, 2.569961e-21, -2.569961e-20, -2.569961e-21, 0, 
    1.003089e-36, -2.569961e-21, -7.709882e-21, 1.027984e-20, 0, 
    7.709882e-21, 0, 0, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 1.003089e-36, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    1.003089e-36, 1.798972e-20, 0, 1.027984e-20, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -1.798972e-20, -1.027984e-20, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, -7.709882e-21, 0, 0, 1.28498e-20, 
    5.139921e-21, 7.709882e-21, 0, 2.569961e-21, 7.709882e-21, 0, 
    -1.027984e-20, 0, 5.139921e-21, 0, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 0, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, 0, -7.709882e-21, 
    -1.027984e-20, 1.027984e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, 0, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, 1.027984e-20, -1.003089e-36, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 1.003089e-36, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 1.541976e-20, 2.569961e-21, -1.28498e-20, -2.569961e-21, 
    7.709882e-21, 0, -7.709882e-21, -1.027984e-20, -2.569961e-21, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, -1.28498e-20, 0, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 5.139921e-21, 0, 0, 0, 
    5.139921e-21, 1.003089e-36, -1.003089e-36, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 0, -7.709882e-21, 7.709882e-21, -1.003089e-36, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, 1.798972e-20, 5.139921e-21, 2.569961e-21, 
    1.003089e-36, -1.003089e-36, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    1.003089e-36, 7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, 1.003089e-36, 0, 
    2.055969e-20, 0, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -1.003089e-36, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 0, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 1.003089e-36, -2.569961e-21, 
    1.798972e-20, 2.569961e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 0, 5.139921e-21, 0, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, 1.798972e-20, 7.709882e-21, 1.28498e-20, 
    2.569961e-21, -1.003089e-36, 0, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21,
  -2.569961e-21, 2.569961e-21, 1.003089e-36, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.003089e-36, 1.28498e-20, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, -1.798972e-20, -2.569961e-21, 
    0, -1.003089e-36, 5.139921e-21, -1.28498e-20, -1.541976e-20, 1.28498e-20, 
    1.003089e-36, -1.027984e-20, 5.139921e-21, 1.28498e-20, -1.541976e-20, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    1.798972e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, -7.709882e-21, 
    1.28498e-20, 2.569961e-21, -1.541976e-20, 1.003089e-36, -7.709882e-21, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -1.027984e-20, 5.139921e-21, 
    1.28498e-20, 7.709882e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -2.312965e-20, 2.569961e-21, 
    -1.027984e-20, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 0, 0, 1.798972e-20, 1.003089e-36, 
    7.709882e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.28498e-20, -2.569961e-21, 0, 
    -2.569961e-21, -5.139921e-21, -2.055969e-20, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, 7.709882e-21, 1.28498e-20, -2.569961e-21, 5.139921e-21, 0, 
    -1.798972e-20, -1.003089e-36, 5.139921e-21, 0, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 1.027984e-20, 
    5.139921e-21, -1.003089e-36, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, 2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 0, -2.569961e-21, 
    1.28498e-20, -2.569961e-21, 0, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, -1.798972e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 0, 
    7.709882e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 1.003089e-36, 
    -2.055969e-20, 1.027984e-20, -1.28498e-20, -5.139921e-21, 0, 
    -1.28498e-20, 7.709882e-21, -7.709882e-21, -1.027984e-20, -1.28498e-20, 
    -5.139921e-21, 1.541976e-20, 1.003089e-36, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 1.541976e-20, 
    0, 2.569961e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, -2.055969e-20, -1.28498e-20, 5.139921e-21, 7.709882e-21, 
    -1.28498e-20, 7.709882e-21, 0, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    1.28498e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.28498e-20, 0, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 1.541976e-20, 0, 
    1.003089e-36, 7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -1.28498e-20, -7.709882e-21, -7.709882e-21, -1.003089e-36, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, 1.28498e-20, 0, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 1.027984e-20, -1.003089e-36, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 0, -5.139921e-21, -1.541976e-20, 
    1.541976e-20, 2.569961e-21, 7.709882e-21, 1.003089e-36, -7.709882e-21, 
    -1.28498e-20, 7.709882e-21, -2.569961e-21, 0, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 1.027984e-20, 1.541976e-20, 0, 1.003089e-36, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, 
    0, -1.027984e-20, -7.709882e-21, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, 1.28498e-20, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 1.798972e-20, 
    1.027984e-20, 7.709882e-21, -5.139921e-21, -7.709882e-21, -7.709882e-21, 
    -1.28498e-20, 7.709882e-21, 7.709882e-21, -1.027984e-20, 7.709882e-21, 
    -5.139921e-21, -1.027984e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, 0, 2.569961e-21, 
    -1.541976e-20, -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21,
  1.027984e-20, 5.139921e-21, -1.003089e-36, 1.027984e-20, 2.569961e-21, 
    1.027984e-20, -1.541976e-20, 0, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 0, 1.541976e-20, 1.798972e-20, 7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -2.569961e-21, -1.003089e-36, 
    5.139921e-21, -7.709882e-21, -7.709882e-21, -1.28498e-20, 1.003089e-36, 
    -7.709882e-21, -7.709882e-21, 1.027984e-20, -7.709882e-21, -1.798972e-20, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -1.28498e-20, 1.28498e-20, -2.569961e-21, -1.027984e-20, 
    0, -5.139921e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -5.139921e-21, -7.709882e-21, 1.003089e-36, 7.709882e-21, 
    -1.28498e-20, 2.569961e-21, -5.139921e-21, -2.569961e-21, 1.541976e-20, 
    -1.798972e-20, -1.027984e-20, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -7.709882e-21, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, -7.709882e-21, -2.569961e-20, 5.139921e-21, 
    -2.569961e-21, 1.28498e-20, 1.541976e-20, -1.28498e-20, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -1.003089e-36, 5.139921e-21, 1.28498e-20, 
    0, -2.569961e-21, 1.027984e-20, -1.027984e-20, -1.541976e-20, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.055969e-20, 
    7.709882e-21, 1.027984e-20, -7.709882e-21, 5.139921e-21, -1.28498e-20, 
    1.027984e-20, -1.541976e-20, -2.569961e-21, 0, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.541976e-20, -2.569961e-21, -1.28498e-20, 1.027984e-20, 0, 
    7.709882e-21, 2.569961e-21, -1.798972e-20, -1.003089e-36, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, -1.28498e-20, 
    1.28498e-20, 1.28498e-20, 2.569961e-21, 1.027984e-20, 0, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -2.055969e-20, 
    -7.709882e-21, -3.083953e-20, -5.139921e-21, 1.541976e-20, 1.003089e-36, 
    -1.28498e-20, 0, -1.541976e-20, -5.139921e-21, 2.569961e-20, 0, 
    -5.139921e-21, -1.798972e-20, -1.28498e-20, 0, 5.139921e-21, 
    -1.28498e-20, 0, 2.569961e-21, -1.28498e-20, 1.541976e-20, 7.709882e-21, 
    1.003089e-36, 0, 2.569961e-21, 2.569961e-21, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, -1.003089e-36, -1.541976e-20, 5.139921e-21, 5.139921e-21, 
    1.003089e-36, 1.027984e-20, 7.709882e-21, 1.003089e-36, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, 0, -1.541976e-20, -2.569961e-21, 
    -2.055969e-20, -1.003089e-36, -5.139921e-21, -2.569961e-21, 
    -2.055969e-20, 2.312965e-20, -2.569961e-21, 1.541976e-20, 1.28498e-20, 
    1.003089e-36, -2.569961e-21, 0, 5.139921e-21, -5.139921e-21, 
    -1.28498e-20, -1.027984e-20, 1.027984e-20, 1.28498e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, 0, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 1.003089e-36, -2.826957e-20, -1.28498e-20, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -1.28498e-20, -2.569961e-21, 5.139921e-21, 1.28498e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 1.003089e-36, 1.798972e-20, -5.139921e-21, 
    1.003089e-36, -1.003089e-36, -2.569961e-21, -5.139921e-21, 1.003089e-36, 
    -7.709882e-21, 1.003089e-36, 1.541976e-20, 5.139921e-21, 2.312965e-20, 
    1.027984e-20, 2.569961e-21, 7.709882e-21, -7.709882e-21, 1.541976e-20, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, -1.28498e-20, 7.709882e-21, 
    1.541976e-20, -1.027984e-20, -1.003089e-36, 5.139921e-21, 0, 
    -7.709882e-21, 1.027984e-20, -1.003089e-36, 2.569961e-21, -1.027984e-20, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    0, -5.139921e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    2.569961e-21, 1.798972e-20, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    2.055969e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, -7.709882e-21, 
    -1.541976e-20, 1.003089e-36, -2.569961e-21, -1.28498e-20, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, -7.709882e-21, -2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -1.541976e-20, -1.28498e-20, 2.569961e-21, -2.569961e-20, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, -1.798972e-20, 0, 5.139921e-21, 
    -7.709882e-21, 5.139921e-21, -1.003089e-36, -7.709882e-21, 5.139921e-21, 
    5.139921e-21,
  2.055969e-20, -1.541976e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, 5.139921e-21, -7.709882e-21, 
    -1.027984e-20, 5.139921e-21, 0, -1.28498e-20, -1.798972e-20, 
    -5.139921e-21, 0, -1.003089e-36, 1.027984e-20, 7.709882e-21, 
    -1.541976e-20, -2.312965e-20, 1.28498e-20, -1.027984e-20, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, 1.003089e-36, -1.541976e-20, -1.28498e-20, 0, 
    -7.709882e-21, 1.541976e-20, 7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -1.28498e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, 2.569961e-21, 
    7.709882e-21, 7.709882e-21, 2.055969e-20, -2.569961e-21, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -2.055969e-20, 1.798972e-20, 1.027984e-20, -2.569961e-21, 
    1.798972e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, 1.798972e-20, 1.28498e-20, 
    2.569961e-21, 2.569961e-21, 1.003089e-36, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -2.055969e-20, 2.569961e-21, 5.139921e-21, -2.055969e-20, 
    -2.826957e-20, -1.003089e-36, -1.027984e-20, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, 2.569961e-21, -7.709882e-21, 2.312965e-20, 5.139921e-21, 
    2.569961e-21, -2.826957e-20, -3.009266e-36, 1.541976e-20, 7.709882e-21, 
    1.003089e-36, -1.027984e-20, -1.027984e-20, -1.798972e-20, 1.798972e-20, 
    -5.139921e-21, 1.798972e-20, 2.312965e-20, 2.055969e-20, -1.027984e-20, 
    -2.569961e-21, -1.027984e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 1.28498e-20, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, 0, 2.055969e-20, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -1.003089e-36, 5.139921e-21, 2.569961e-21, -1.798972e-20, -1.003089e-36, 
    -7.709882e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    0, 1.003089e-36, 2.569961e-21, 1.027984e-20, 7.709882e-21, 1.027984e-20, 
    1.003089e-36, -2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -1.798972e-20, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, -5.139921e-21, 1.003089e-36, 1.541976e-20, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, 0, 2.312965e-20, 
    7.709882e-21, 1.798972e-20, 1.003089e-36, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 2.312965e-20, -1.027984e-20, 1.798972e-20, 
    0, -2.569961e-21, 2.312965e-20, 1.28498e-20, 2.569961e-21, 1.541976e-20, 
    2.055969e-20, -1.798972e-20, 1.28498e-20, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, 1.798972e-20, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 1.28498e-20, 
    -7.709882e-21, -2.569961e-21, 1.798972e-20, 5.139921e-21, 5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    1.28498e-20, 0, 5.139921e-21, -2.569961e-21, -7.709882e-21, 0, 
    2.569961e-21, -2.055969e-20, -1.027984e-20, -5.139921e-21, -1.28498e-20, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 1.541976e-20, -2.569961e-21, -1.003089e-36, 
    2.569961e-20, -2.569961e-21, -1.027984e-20, 0, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 1.28498e-20, -2.569961e-20, 2.569961e-21, 5.139921e-21, 
    -1.541976e-20, 7.709882e-21, -1.28498e-20, 2.569961e-21, -5.139921e-21, 
    -1.003089e-36, 1.541976e-20, -5.139921e-21, 7.709882e-21, 1.003089e-36, 
    7.709882e-21, 2.569961e-21, -1.798972e-20, -5.139921e-21, -2.569961e-21, 
    1.798972e-20, 2.569961e-21, -7.709882e-21, -2.569961e-21, -1.003089e-36, 
    5.139921e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -1.003089e-36, 1.027984e-20, -1.027984e-20, 2.312965e-20, 
    -5.139921e-21, 1.798972e-20, 7.709882e-21, 7.709882e-21, 2.055969e-20, 
    -7.709882e-21, 5.139921e-21, 1.003089e-36, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -7.709882e-21, 1.003089e-36, 1.798972e-20, 
    -2.312965e-20, 0, -1.798972e-20, 1.027984e-20, 7.709882e-21, 
    -7.709882e-21, 1.28498e-20, 2.569961e-21, -1.28498e-20, 1.027984e-20, 
    -1.28498e-20, -7.709882e-21, -7.709882e-21, -1.28498e-20, 5.139921e-21, 
    2.569961e-21, -1.541976e-20, 1.003089e-36, -1.027984e-20, -1.027984e-20, 
    2.569961e-20, -2.569961e-21, -7.709882e-21, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 1.003089e-36, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, 1.027984e-20, -7.709882e-21, 1.798972e-20, 1.798972e-20, 
    -1.541976e-20,
  6.259376e-29, 6.259382e-29, 6.259381e-29, 6.259386e-29, 6.259384e-29, 
    6.259387e-29, 6.259378e-29, 6.259382e-29, 6.259379e-29, 6.259376e-29, 
    6.259396e-29, 6.259387e-29, 6.259406e-29, 6.2594e-29, 6.259415e-29, 
    6.259405e-29, 6.259417e-29, 6.259415e-29, 6.259422e-29, 6.25942e-29, 
    6.259429e-29, 6.259423e-29, 6.259434e-29, 6.259428e-29, 6.259428e-29, 
    6.259423e-29, 6.259388e-29, 6.259394e-29, 6.259388e-29, 6.259389e-29, 
    6.259388e-29, 6.259384e-29, 6.259381e-29, 6.259376e-29, 6.259376e-29, 
    6.259381e-29, 6.259389e-29, 6.259386e-29, 6.259394e-29, 6.259394e-29, 
    6.259402e-29, 6.259398e-29, 6.259413e-29, 6.259408e-29, 6.25942e-29, 
    6.259417e-29, 6.25942e-29, 6.259419e-29, 6.25942e-29, 6.259416e-29, 
    6.259417e-29, 6.259414e-29, 6.259399e-29, 6.259404e-29, 6.25939e-29, 
    6.259382e-29, 6.259378e-29, 6.259374e-29, 6.259375e-29, 6.259375e-29, 
    6.259381e-29, 6.259385e-29, 6.259389e-29, 6.259391e-29, 6.259394e-29, 
    6.259401e-29, 6.259405e-29, 6.259413e-29, 6.259411e-29, 6.259414e-29, 
    6.259417e-29, 6.259421e-29, 6.25942e-29, 6.259422e-29, 6.259414e-29, 
    6.259419e-29, 6.259411e-29, 6.259413e-29, 6.259394e-29, 6.259387e-29, 
    6.259384e-29, 6.259381e-29, 6.259375e-29, 6.259379e-29, 6.259378e-29, 
    6.259382e-29, 6.259384e-29, 6.259383e-29, 6.259391e-29, 6.259388e-29, 
    6.259405e-29, 6.259398e-29, 6.259416e-29, 6.259412e-29, 6.259417e-29, 
    6.259415e-29, 6.25942e-29, 6.259415e-29, 6.259423e-29, 6.259425e-29, 
    6.259423e-29, 6.259428e-29, 6.259415e-29, 6.25942e-29, 6.259383e-29, 
    6.259384e-29, 6.259384e-29, 6.25938e-29, 6.259379e-29, 6.259376e-29, 
    6.259379e-29, 6.259381e-29, 6.259385e-29, 6.259387e-29, 6.259389e-29, 
    6.259394e-29, 6.259399e-29, 6.259407e-29, 6.259412e-29, 6.259416e-29, 
    6.259414e-29, 6.259416e-29, 6.259413e-29, 6.259413e-29, 6.259424e-29, 
    6.259417e-29, 6.259427e-29, 6.259426e-29, 6.259422e-29, 6.259426e-29, 
    6.259384e-29, 6.259382e-29, 6.259378e-29, 6.259381e-29, 6.259375e-29, 
    6.259379e-29, 6.259381e-29, 6.259388e-29, 6.25939e-29, 6.259391e-29, 
    6.259394e-29, 6.259399e-29, 6.259405e-29, 6.259411e-29, 6.259417e-29, 
    6.259417e-29, 6.259417e-29, 6.259418e-29, 6.259415e-29, 6.259419e-29, 
    6.259419e-29, 6.259417e-29, 6.259426e-29, 6.259424e-29, 6.259426e-29, 
    6.259425e-29, 6.259382e-29, 6.259385e-29, 6.259384e-29, 6.259385e-29, 
    6.259384e-29, 6.259391e-29, 6.259393e-29, 6.259402e-29, 6.259398e-29, 
    6.259405e-29, 6.259399e-29, 6.2594e-29, 6.259405e-29, 6.259399e-29, 
    6.259411e-29, 6.259403e-29, 6.259418e-29, 6.25941e-29, 6.259419e-29, 
    6.259417e-29, 6.259419e-29, 6.259422e-29, 6.259425e-29, 6.25943e-29, 
    6.259429e-29, 6.259433e-29, 6.259388e-29, 6.25939e-29, 6.25939e-29, 
    6.259393e-29, 6.259395e-29, 6.2594e-29, 6.259407e-29, 6.259404e-29, 
    6.25941e-29, 6.25941e-29, 6.259403e-29, 6.259408e-29, 6.259392e-29, 
    6.259395e-29, 6.259393e-29, 6.259388e-29, 6.259405e-29, 6.259396e-29, 
    6.259413e-29, 6.259408e-29, 6.259422e-29, 6.259414e-29, 6.259428e-29, 
    6.259434e-29, 6.259439e-29, 6.259446e-29, 6.259392e-29, 6.25939e-29, 
    6.259393e-29, 6.259398e-29, 6.259402e-29, 6.259408e-29, 6.259408e-29, 
    6.25941e-29, 6.259413e-29, 6.259414e-29, 6.25941e-29, 6.259415e-29, 
    6.259395e-29, 6.259406e-29, 6.25939e-29, 6.259394e-29, 6.259398e-29, 
    6.259396e-29, 6.259404e-29, 6.259406e-29, 6.259413e-29, 6.25941e-29, 
    6.259432e-29, 6.259422e-29, 6.25945e-29, 6.259443e-29, 6.25939e-29, 
    6.259392e-29, 6.259401e-29, 6.259396e-29, 6.259408e-29, 6.259411e-29, 
    6.259414e-29, 6.259417e-29, 6.259417e-29, 6.259419e-29, 6.259416e-29, 
    6.259419e-29, 6.259408e-29, 6.259413e-29, 6.2594e-29, 6.259403e-29, 
    6.259401e-29, 6.2594e-29, 6.259405e-29, 6.25941e-29, 6.25941e-29, 
    6.259412e-29, 6.259417e-29, 6.259408e-29, 6.259434e-29, 6.259418e-29, 
    6.259394e-29, 6.259399e-29, 6.2594e-29, 6.259398e-29, 6.259411e-29, 
    6.259407e-29, 6.259419e-29, 6.259416e-29, 6.259421e-29, 6.259418e-29, 
    6.259417e-29, 6.259414e-29, 6.259412e-29, 6.259407e-29, 6.259402e-29, 
    6.259399e-29, 6.259399e-29, 6.259404e-29, 6.25941e-29, 6.259417e-29, 
    6.259416e-29, 6.25942e-29, 6.259407e-29, 6.259413e-29, 6.259411e-29, 
    6.259416e-29, 6.259404e-29, 6.259414e-29, 6.259402e-29, 6.259403e-29, 
    6.259407e-29, 6.259413e-29, 6.259415e-29, 6.259416e-29, 6.259416e-29, 
    6.259411e-29, 6.25941e-29, 6.259406e-29, 6.259405e-29, 6.259402e-29, 
    6.259401e-29, 6.259402e-29, 6.259405e-29, 6.259411e-29, 6.259416e-29, 
    6.259422e-29, 6.259423e-29, 6.25943e-29, 6.259425e-29, 6.259434e-29, 
    6.259426e-29, 6.25944e-29, 6.259415e-29, 6.259426e-29, 6.259407e-29, 
    6.259408e-29, 6.259412e-29, 6.259421e-29, 6.259416e-29, 6.259422e-29, 
    6.25941e-29, 6.259404e-29, 6.259402e-29, 6.259399e-29, 6.259402e-29, 
    6.259402e-29, 6.259405e-29, 6.259404e-29, 6.259411e-29, 6.259407e-29, 
    6.259417e-29, 6.259422e-29, 6.259432e-29, 6.25944e-29, 6.259446e-29, 
    6.259449e-29, 6.25945e-29, 6.25945e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.137825e-10, 2.147324e-10, 2.145478e-10, 2.15314e-10, 2.14889e-10, 
    2.153907e-10, 2.139751e-10, 2.147701e-10, 2.142626e-10, 2.13868e-10, 
    2.168012e-10, 2.153482e-10, 2.18311e-10, 2.173841e-10, 2.197128e-10, 
    2.181667e-10, 2.200246e-10, 2.196683e-10, 2.20741e-10, 2.204336e-10, 
    2.218058e-10, 2.208828e-10, 2.225172e-10, 2.215854e-10, 2.217311e-10, 
    2.208524e-10, 2.156407e-10, 2.166203e-10, 2.155826e-10, 2.157223e-10, 
    2.156596e-10, 2.148977e-10, 2.145138e-10, 2.137099e-10, 2.138559e-10, 
    2.144463e-10, 2.157851e-10, 2.153307e-10, 2.164761e-10, 2.164503e-10, 
    2.177257e-10, 2.171506e-10, 2.192947e-10, 2.186852e-10, 2.204465e-10, 
    2.200035e-10, 2.204256e-10, 2.202977e-10, 2.204273e-10, 2.197777e-10, 
    2.20056e-10, 2.194844e-10, 2.172583e-10, 2.179124e-10, 2.159616e-10, 
    2.147888e-10, 2.140099e-10, 2.134573e-10, 2.135354e-10, 2.136844e-10, 
    2.144498e-10, 2.151695e-10, 2.15718e-10, 2.16085e-10, 2.164466e-10, 
    2.17541e-10, 2.181204e-10, 2.194179e-10, 2.191838e-10, 2.195804e-10, 
    2.199594e-10, 2.205958e-10, 2.20491e-10, 2.207714e-10, 2.1957e-10, 
    2.203684e-10, 2.190504e-10, 2.194108e-10, 2.165447e-10, 2.154533e-10, 
    2.149893e-10, 2.145833e-10, 2.135955e-10, 2.142776e-10, 2.140087e-10, 
    2.146485e-10, 2.15055e-10, 2.14854e-10, 2.16095e-10, 2.156125e-10, 
    2.181547e-10, 2.170596e-10, 2.199152e-10, 2.192318e-10, 2.20079e-10, 
    2.196467e-10, 2.203875e-10, 2.197208e-10, 2.208757e-10, 2.211272e-10, 
    2.209554e-10, 2.216156e-10, 2.196838e-10, 2.204256e-10, 2.148483e-10, 
    2.148811e-10, 2.150339e-10, 2.143623e-10, 2.143212e-10, 2.137059e-10, 
    2.142534e-10, 2.144866e-10, 2.150786e-10, 2.154288e-10, 2.157617e-10, 
    2.164936e-10, 2.173112e-10, 2.184545e-10, 2.192761e-10, 2.198269e-10, 
    2.194891e-10, 2.197873e-10, 2.19454e-10, 2.192978e-10, 2.21033e-10, 
    2.200586e-10, 2.215207e-10, 2.214398e-10, 2.20778e-10, 2.214489e-10, 
    2.149041e-10, 2.147155e-10, 2.140603e-10, 2.14573e-10, 2.136389e-10, 
    2.141617e-10, 2.144624e-10, 2.156225e-10, 2.158775e-10, 2.161139e-10, 
    2.165808e-10, 2.1718e-10, 2.182313e-10, 2.191462e-10, 2.199815e-10, 
    2.199203e-10, 2.199418e-10, 2.201284e-10, 2.196662e-10, 2.202043e-10, 
    2.202946e-10, 2.200585e-10, 2.214289e-10, 2.210374e-10, 2.21438e-10, 
    2.211831e-10, 2.147768e-10, 2.150943e-10, 2.149227e-10, 2.152454e-10, 
    2.150181e-10, 2.160288e-10, 2.163319e-10, 2.177503e-10, 2.171682e-10, 
    2.180947e-10, 2.172623e-10, 2.174098e-10, 2.181249e-10, 2.173073e-10, 
    2.190957e-10, 2.178832e-10, 2.201357e-10, 2.189246e-10, 2.202116e-10, 
    2.199779e-10, 2.203648e-10, 2.207114e-10, 2.211474e-10, 2.21952e-10, 
    2.217657e-10, 2.224386e-10, 2.155677e-10, 2.159796e-10, 2.159433e-10, 
    2.163744e-10, 2.166932e-10, 2.173843e-10, 2.184928e-10, 2.18076e-10, 
    2.188413e-10, 2.18995e-10, 2.178323e-10, 2.185461e-10, 2.162553e-10, 
    2.166253e-10, 2.16405e-10, 2.156002e-10, 2.18172e-10, 2.16852e-10, 
    2.192897e-10, 2.185745e-10, 2.206619e-10, 2.196237e-10, 2.216631e-10, 
    2.22535e-10, 2.233558e-10, 2.24315e-10, 2.162044e-10, 2.159245e-10, 
    2.164257e-10, 2.171191e-10, 2.177626e-10, 2.186181e-10, 2.187056e-10, 
    2.188659e-10, 2.192811e-10, 2.196302e-10, 2.189166e-10, 2.197177e-10, 
    2.167111e-10, 2.182866e-10, 2.158187e-10, 2.165617e-10, 2.170782e-10, 
    2.168517e-10, 2.180283e-10, 2.183057e-10, 2.194328e-10, 2.188502e-10, 
    2.223198e-10, 2.207845e-10, 2.250456e-10, 2.238545e-10, 2.158268e-10, 
    2.162035e-10, 2.175147e-10, 2.168908e-10, 2.186752e-10, 2.191145e-10, 
    2.194716e-10, 2.199282e-10, 2.199775e-10, 2.20248e-10, 2.198047e-10, 
    2.202305e-10, 2.186199e-10, 2.193396e-10, 2.173648e-10, 2.178454e-10, 
    2.176243e-10, 2.173818e-10, 2.181303e-10, 2.189278e-10, 2.189449e-10, 
    2.192006e-10, 2.199212e-10, 2.186825e-10, 2.225178e-10, 2.201489e-10, 
    2.166143e-10, 2.173399e-10, 2.174436e-10, 2.171625e-10, 2.190705e-10, 
    2.183791e-10, 2.202414e-10, 2.197381e-10, 2.205628e-10, 2.20153e-10, 
    2.200927e-10, 2.195663e-10, 2.192386e-10, 2.184108e-10, 2.177373e-10, 
    2.172033e-10, 2.173275e-10, 2.17914e-10, 2.189766e-10, 2.199819e-10, 
    2.197617e-10, 2.205001e-10, 2.185458e-10, 2.193652e-10, 2.190485e-10, 
    2.198744e-10, 2.180649e-10, 2.196056e-10, 2.176711e-10, 2.178407e-10, 
    2.183654e-10, 2.194207e-10, 2.196544e-10, 2.199037e-10, 2.197498e-10, 
    2.190036e-10, 2.188813e-10, 2.183526e-10, 2.182066e-10, 2.178038e-10, 
    2.174703e-10, 2.17775e-10, 2.18095e-10, 2.190039e-10, 2.198231e-10, 
    2.207163e-10, 2.209349e-10, 2.219786e-10, 2.211289e-10, 2.22531e-10, 
    2.213389e-10, 2.234028e-10, 2.19695e-10, 2.213039e-10, 2.183893e-10, 
    2.187032e-10, 2.192711e-10, 2.205737e-10, 2.198705e-10, 2.20693e-10, 
    2.188765e-10, 2.179343e-10, 2.176905e-10, 2.172357e-10, 2.177009e-10, 
    2.176631e-10, 2.181083e-10, 2.179652e-10, 2.190341e-10, 2.184599e-10, 
    2.200911e-10, 2.206865e-10, 2.223681e-10, 2.23399e-10, 2.244488e-10, 
    2.249122e-10, 2.250533e-10, 2.251123e-10 ;

 SOIL2N_TO_SOIL3N =
  1.527018e-11, 1.533803e-11, 1.532484e-11, 1.537957e-11, 1.534921e-11, 
    1.538505e-11, 1.528394e-11, 1.534072e-11, 1.530447e-11, 1.527629e-11, 
    1.54858e-11, 1.538202e-11, 1.559364e-11, 1.552743e-11, 1.569377e-11, 
    1.558334e-11, 1.571604e-11, 1.569059e-11, 1.576721e-11, 1.574526e-11, 
    1.584327e-11, 1.577734e-11, 1.589409e-11, 1.582753e-11, 1.583794e-11, 
    1.577517e-11, 1.54029e-11, 1.547288e-11, 1.539876e-11, 1.540874e-11, 
    1.540426e-11, 1.534984e-11, 1.532241e-11, 1.526499e-11, 1.527542e-11, 
    1.531759e-11, 1.541322e-11, 1.538076e-11, 1.546258e-11, 1.546073e-11, 
    1.555183e-11, 1.551076e-11, 1.56639e-11, 1.562037e-11, 1.574618e-11, 
    1.571454e-11, 1.574469e-11, 1.573555e-11, 1.574481e-11, 1.56984e-11, 
    1.571829e-11, 1.567746e-11, 1.551845e-11, 1.556517e-11, 1.542583e-11, 
    1.534205e-11, 1.528642e-11, 1.524695e-11, 1.525253e-11, 1.526317e-11, 
    1.531784e-11, 1.536925e-11, 1.540843e-11, 1.543464e-11, 1.546047e-11, 
    1.553864e-11, 1.558003e-11, 1.56727e-11, 1.565598e-11, 1.568431e-11, 
    1.571139e-11, 1.575684e-11, 1.574936e-11, 1.576938e-11, 1.568357e-11, 
    1.57406e-11, 1.564646e-11, 1.56722e-11, 1.546748e-11, 1.538952e-11, 
    1.535638e-11, 1.532738e-11, 1.525682e-11, 1.530554e-11, 1.528634e-11, 
    1.533203e-11, 1.536107e-11, 1.534671e-11, 1.543536e-11, 1.540089e-11, 
    1.558248e-11, 1.550426e-11, 1.570823e-11, 1.565941e-11, 1.571993e-11, 
    1.568905e-11, 1.574196e-11, 1.569434e-11, 1.577684e-11, 1.57948e-11, 
    1.578253e-11, 1.582969e-11, 1.56917e-11, 1.574469e-11, 1.534631e-11, 
    1.534865e-11, 1.535956e-11, 1.531159e-11, 1.530866e-11, 1.526471e-11, 
    1.530382e-11, 1.532047e-11, 1.536276e-11, 1.538777e-11, 1.541155e-11, 
    1.546383e-11, 1.552223e-11, 1.560389e-11, 1.566258e-11, 1.570192e-11, 
    1.56778e-11, 1.569909e-11, 1.567529e-11, 1.566413e-11, 1.578807e-11, 
    1.571847e-11, 1.58229e-11, 1.581713e-11, 1.576986e-11, 1.581778e-11, 
    1.53503e-11, 1.533682e-11, 1.529002e-11, 1.532664e-11, 1.525992e-11, 
    1.529727e-11, 1.531874e-11, 1.540161e-11, 1.541982e-11, 1.543671e-11, 
    1.547006e-11, 1.551286e-11, 1.558795e-11, 1.56533e-11, 1.571296e-11, 
    1.570859e-11, 1.571013e-11, 1.572346e-11, 1.569044e-11, 1.572888e-11, 
    1.573533e-11, 1.571846e-11, 1.581635e-11, 1.578838e-11, 1.5817e-11, 
    1.579879e-11, 1.53412e-11, 1.536388e-11, 1.535162e-11, 1.537467e-11, 
    1.535843e-11, 1.543063e-11, 1.545228e-11, 1.555359e-11, 1.551202e-11, 
    1.557819e-11, 1.551874e-11, 1.552927e-11, 1.558035e-11, 1.552195e-11, 
    1.564969e-11, 1.556308e-11, 1.572398e-11, 1.563747e-11, 1.57294e-11, 
    1.571271e-11, 1.574034e-11, 1.57651e-11, 1.579624e-11, 1.585371e-11, 
    1.584041e-11, 1.588847e-11, 1.539769e-11, 1.542711e-11, 1.542452e-11, 
    1.545532e-11, 1.547809e-11, 1.552745e-11, 1.560663e-11, 1.557686e-11, 
    1.563152e-11, 1.56425e-11, 1.555945e-11, 1.561043e-11, 1.544681e-11, 
    1.547324e-11, 1.54575e-11, 1.540001e-11, 1.558371e-11, 1.548943e-11, 
    1.566355e-11, 1.561246e-11, 1.576157e-11, 1.568741e-11, 1.583308e-11, 
    1.589536e-11, 1.595399e-11, 1.60225e-11, 1.544317e-11, 1.542318e-11, 
    1.545898e-11, 1.55085e-11, 1.555447e-11, 1.561558e-11, 1.562183e-11, 
    1.563328e-11, 1.566294e-11, 1.568787e-11, 1.56369e-11, 1.569412e-11, 
    1.547936e-11, 1.55919e-11, 1.541562e-11, 1.546869e-11, 1.550559e-11, 
    1.54894e-11, 1.557345e-11, 1.559326e-11, 1.567377e-11, 1.563216e-11, 
    1.587998e-11, 1.577032e-11, 1.607468e-11, 1.598961e-11, 1.54162e-11, 
    1.544311e-11, 1.553676e-11, 1.54922e-11, 1.561966e-11, 1.565104e-11, 
    1.567655e-11, 1.570915e-11, 1.571268e-11, 1.5732e-11, 1.570034e-11, 
    1.573075e-11, 1.561571e-11, 1.566712e-11, 1.552606e-11, 1.556039e-11, 
    1.554459e-11, 1.552727e-11, 1.558074e-11, 1.56377e-11, 1.563892e-11, 
    1.565719e-11, 1.570865e-11, 1.562018e-11, 1.589413e-11, 1.572492e-11, 
    1.547245e-11, 1.552428e-11, 1.553169e-11, 1.551161e-11, 1.564789e-11, 
    1.559851e-11, 1.573153e-11, 1.569558e-11, 1.575449e-11, 1.572521e-11, 
    1.57209e-11, 1.568331e-11, 1.56599e-11, 1.560077e-11, 1.555266e-11, 
    1.551452e-11, 1.552339e-11, 1.556529e-11, 1.564118e-11, 1.5713e-11, 
    1.569726e-11, 1.575001e-11, 1.561042e-11, 1.566894e-11, 1.564632e-11, 
    1.570531e-11, 1.557606e-11, 1.568611e-11, 1.554794e-11, 1.556005e-11, 
    1.559753e-11, 1.567291e-11, 1.56896e-11, 1.570741e-11, 1.569642e-11, 
    1.564311e-11, 1.563438e-11, 1.559662e-11, 1.558619e-11, 1.555741e-11, 
    1.553359e-11, 1.555536e-11, 1.557821e-11, 1.564314e-11, 1.570165e-11, 
    1.576545e-11, 1.578107e-11, 1.585561e-11, 1.579492e-11, 1.589507e-11, 
    1.580992e-11, 1.595734e-11, 1.56925e-11, 1.580742e-11, 1.559923e-11, 
    1.562166e-11, 1.566222e-11, 1.575527e-11, 1.570503e-11, 1.576378e-11, 
    1.563404e-11, 1.556673e-11, 1.554932e-11, 1.551684e-11, 1.555007e-11, 
    1.554736e-11, 1.557916e-11, 1.556894e-11, 1.564529e-11, 1.560428e-11, 
    1.57208e-11, 1.576332e-11, 1.588343e-11, 1.595708e-11, 1.603206e-11, 
    1.606516e-11, 1.607523e-11, 1.607945e-11 ;

 SOIL2N_vr =
  1.818724, 1.818725, 1.818725, 1.818726, 1.818725, 1.818726, 1.818724, 
    1.818725, 1.818724, 1.818724, 1.818728, 1.818726, 1.818731, 1.818729, 
    1.818733, 1.81873, 1.818733, 1.818733, 1.818734, 1.818734, 1.818736, 
    1.818735, 1.818737, 1.818736, 1.818736, 1.818735, 1.818726, 1.818728, 
    1.818726, 1.818727, 1.818726, 1.818725, 1.818725, 1.818723, 1.818724, 
    1.818725, 1.818727, 1.818726, 1.818728, 1.818728, 1.81873, 1.818729, 
    1.818732, 1.818731, 1.818734, 1.818733, 1.818734, 1.818734, 1.818734, 
    1.818733, 1.818733, 1.818732, 1.818729, 1.81873, 1.818727, 1.818725, 
    1.818724, 1.818723, 1.818723, 1.818723, 1.818725, 1.818726, 1.818727, 
    1.818727, 1.818728, 1.818729, 1.81873, 1.818732, 1.818732, 1.818733, 
    1.818733, 1.818734, 1.818734, 1.818734, 1.818733, 1.818734, 1.818732, 
    1.818732, 1.818728, 1.818726, 1.818725, 1.818725, 1.818723, 1.818724, 
    1.818724, 1.818725, 1.818725, 1.818725, 1.818727, 1.818726, 1.81873, 
    1.818729, 1.818733, 1.818732, 1.818733, 1.818733, 1.818734, 1.818733, 
    1.818735, 1.818735, 1.818735, 1.818736, 1.818733, 1.818734, 1.818725, 
    1.818725, 1.818725, 1.818724, 1.818724, 1.818723, 1.818724, 1.818725, 
    1.818726, 1.818726, 1.818727, 1.818728, 1.818729, 1.818731, 1.818732, 
    1.818733, 1.818732, 1.818733, 1.818732, 1.818732, 1.818735, 1.818733, 
    1.818736, 1.818735, 1.818734, 1.818735, 1.818725, 1.818725, 1.818724, 
    1.818725, 1.818723, 1.818724, 1.818725, 1.818726, 1.818727, 1.818727, 
    1.818728, 1.818729, 1.81873, 1.818732, 1.818733, 1.818733, 1.818733, 
    1.818733, 1.818733, 1.818734, 1.818734, 1.818733, 1.818735, 1.818735, 
    1.818735, 1.818735, 1.818725, 1.818726, 1.818725, 1.818726, 1.818725, 
    1.818727, 1.818727, 1.81873, 1.818729, 1.81873, 1.818729, 1.818729, 
    1.81873, 1.818729, 1.818732, 1.81873, 1.818733, 1.818732, 1.818734, 
    1.818733, 1.818734, 1.818734, 1.818735, 1.818736, 1.818736, 1.818737, 
    1.818726, 1.818727, 1.818727, 1.818728, 1.818728, 1.818729, 1.818731, 
    1.81873, 1.818731, 1.818732, 1.81873, 1.818731, 1.818727, 1.818728, 
    1.818728, 1.818726, 1.81873, 1.818728, 1.818732, 1.818731, 1.818734, 
    1.818733, 1.818736, 1.818737, 1.818738, 1.81874, 1.818727, 1.818727, 
    1.818728, 1.818729, 1.81873, 1.818731, 1.818731, 1.818731, 1.818732, 
    1.818733, 1.818732, 1.818733, 1.818728, 1.818731, 1.818727, 1.818728, 
    1.818729, 1.818728, 1.81873, 1.818731, 1.818732, 1.818731, 1.818737, 
    1.818734, 1.818741, 1.818739, 1.818727, 1.818727, 1.818729, 1.818728, 
    1.818731, 1.818732, 1.818732, 1.818733, 1.818733, 1.818734, 1.818733, 
    1.818734, 1.818731, 1.818732, 1.818729, 1.81873, 1.81873, 1.818729, 
    1.81873, 1.818732, 1.818732, 1.818732, 1.818733, 1.818731, 1.818737, 
    1.818733, 1.818728, 1.818729, 1.818729, 1.818729, 1.818732, 1.818731, 
    1.818734, 1.818733, 1.818734, 1.818733, 1.818733, 1.818733, 1.818732, 
    1.818731, 1.81873, 1.818729, 1.818729, 1.81873, 1.818732, 1.818733, 
    1.818733, 1.818734, 1.818731, 1.818732, 1.818732, 1.818733, 1.81873, 
    1.818733, 1.81873, 1.81873, 1.818731, 1.818732, 1.818733, 1.818733, 
    1.818733, 1.818732, 1.818731, 1.818731, 1.81873, 1.81873, 1.818729, 
    1.81873, 1.81873, 1.818732, 1.818733, 1.818734, 1.818735, 1.818736, 
    1.818735, 1.818737, 1.818735, 1.818738, 1.818733, 1.818735, 1.818731, 
    1.818731, 1.818732, 1.818734, 1.818733, 1.818734, 1.818731, 1.81873, 
    1.81873, 1.818729, 1.81873, 1.81873, 1.81873, 1.81873, 1.818732, 
    1.818731, 1.818733, 1.818734, 1.818737, 1.818738, 1.81874, 1.818741, 
    1.818741, 1.818741,
  1.81867, 1.818672, 1.818672, 1.818673, 1.818673, 1.818674, 1.818671, 
    1.818672, 1.818671, 1.818671, 1.818676, 1.818673, 1.818679, 1.818678, 
    1.818682, 1.818679, 1.818683, 1.818682, 1.818684, 1.818684, 1.818686, 
    1.818684, 1.818688, 1.818686, 1.818686, 1.818684, 1.818674, 1.818676, 
    1.818674, 1.818674, 1.818674, 1.818673, 1.818672, 1.81867, 1.818671, 
    1.818672, 1.818674, 1.818673, 1.818676, 1.818676, 1.818678, 1.818677, 
    1.818681, 1.81868, 1.818684, 1.818683, 1.818684, 1.818683, 1.818684, 
    1.818682, 1.818683, 1.818682, 1.818677, 1.818679, 1.818675, 1.818672, 
    1.818671, 1.81867, 1.81867, 1.81867, 1.818672, 1.818673, 1.818674, 
    1.818675, 1.818676, 1.818678, 1.818679, 1.818681, 1.818681, 1.818682, 
    1.818683, 1.818684, 1.818684, 1.818684, 1.818682, 1.818683, 1.818681, 
    1.818681, 1.818676, 1.818674, 1.818673, 1.818672, 1.81867, 1.818671, 
    1.818671, 1.818672, 1.818673, 1.818673, 1.818675, 1.818674, 1.818679, 
    1.818677, 1.818682, 1.818681, 1.818683, 1.818682, 1.818683, 1.818682, 
    1.818684, 1.818685, 1.818684, 1.818686, 1.818682, 1.818684, 1.818673, 
    1.818673, 1.818673, 1.818672, 1.818671, 1.81867, 1.818671, 1.818672, 
    1.818673, 1.818674, 1.818674, 1.818676, 1.818677, 1.81868, 1.818681, 
    1.818682, 1.818682, 1.818682, 1.818682, 1.818681, 1.818685, 1.818683, 
    1.818686, 1.818685, 1.818684, 1.818686, 1.818673, 1.818672, 1.818671, 
    1.818672, 1.81867, 1.818671, 1.818672, 1.818674, 1.818675, 1.818675, 
    1.818676, 1.818677, 1.818679, 1.818681, 1.818683, 1.818683, 1.818683, 
    1.818683, 1.818682, 1.818683, 1.818683, 1.818683, 1.818685, 1.818685, 
    1.818685, 1.818685, 1.818672, 1.818673, 1.818673, 1.818673, 1.818673, 
    1.818675, 1.818675, 1.818678, 1.818677, 1.818679, 1.818677, 1.818678, 
    1.818679, 1.818677, 1.818681, 1.818678, 1.818683, 1.818681, 1.818683, 
    1.818683, 1.818683, 1.818684, 1.818685, 1.818686, 1.818686, 1.818687, 
    1.818674, 1.818675, 1.818675, 1.818676, 1.818676, 1.818678, 1.81868, 
    1.818679, 1.81868, 1.818681, 1.818678, 1.81868, 1.818675, 1.818676, 
    1.818676, 1.818674, 1.818679, 1.818676, 1.818681, 1.81868, 1.818684, 
    1.818682, 1.818686, 1.818688, 1.818689, 1.818691, 1.818675, 1.818675, 
    1.818676, 1.818677, 1.818678, 1.81868, 1.81868, 1.81868, 1.818681, 
    1.818682, 1.818681, 1.818682, 1.818676, 1.818679, 1.818674, 1.818676, 
    1.818677, 1.818676, 1.818679, 1.818679, 1.818682, 1.81868, 1.818687, 
    1.818684, 1.818692, 1.81869, 1.818674, 1.818675, 1.818678, 1.818677, 
    1.81868, 1.818681, 1.818682, 1.818683, 1.818683, 1.818683, 1.818682, 
    1.818683, 1.81868, 1.818681, 1.818678, 1.818678, 1.818678, 1.818678, 
    1.818679, 1.818681, 1.818681, 1.818681, 1.818683, 1.81868, 1.818688, 
    1.818683, 1.818676, 1.818677, 1.818678, 1.818677, 1.818681, 1.818679, 
    1.818683, 1.818682, 1.818684, 1.818683, 1.818683, 1.818682, 1.818681, 
    1.81868, 1.818678, 1.818677, 1.818677, 1.818679, 1.818681, 1.818683, 
    1.818682, 1.818684, 1.81868, 1.818681, 1.818681, 1.818682, 1.818679, 
    1.818682, 1.818678, 1.818678, 1.818679, 1.818681, 1.818682, 1.818682, 
    1.818682, 1.818681, 1.81868, 1.818679, 1.818679, 1.818678, 1.818678, 
    1.818678, 1.818679, 1.818681, 1.818682, 1.818684, 1.818684, 1.818686, 
    1.818685, 1.818688, 1.818685, 1.818689, 1.818682, 1.818685, 1.818679, 
    1.81868, 1.818681, 1.818684, 1.818682, 1.818684, 1.81868, 1.818679, 
    1.818678, 1.818677, 1.818678, 1.818678, 1.818679, 1.818679, 1.818681, 
    1.81868, 1.818683, 1.818684, 1.818687, 1.818689, 1.818691, 1.818692, 
    1.818693, 1.818693,
  1.81864, 1.818642, 1.818642, 1.818644, 1.818643, 1.818644, 1.818641, 
    1.818643, 1.818641, 1.818641, 1.818647, 1.818644, 1.81865, 1.818648, 
    1.818653, 1.81865, 1.818654, 1.818653, 1.818655, 1.818655, 1.818658, 
    1.818656, 1.818659, 1.818657, 1.818658, 1.818656, 1.818644, 1.818647, 
    1.818644, 1.818645, 1.818645, 1.818643, 1.818642, 1.81864, 1.818641, 
    1.818642, 1.818645, 1.818644, 1.818646, 1.818646, 1.818649, 1.818648, 
    1.818652, 1.818651, 1.818655, 1.818654, 1.818655, 1.818654, 1.818655, 
    1.818653, 1.818654, 1.818653, 1.818648, 1.818649, 1.818645, 1.818643, 
    1.818641, 1.81864, 1.81864, 1.81864, 1.818642, 1.818643, 1.818645, 
    1.818645, 1.818646, 1.818649, 1.81865, 1.818653, 1.818652, 1.818653, 
    1.818654, 1.818655, 1.818655, 1.818655, 1.818653, 1.818655, 1.818652, 
    1.818653, 1.818646, 1.818644, 1.818643, 1.818642, 1.81864, 1.818642, 
    1.818641, 1.818642, 1.818643, 1.818643, 1.818645, 1.818644, 1.81865, 
    1.818648, 1.818654, 1.818652, 1.818654, 1.818653, 1.818655, 1.818653, 
    1.818656, 1.818656, 1.818656, 1.818657, 1.818653, 1.818655, 1.818643, 
    1.818643, 1.818643, 1.818642, 1.818642, 1.81864, 1.818641, 1.818642, 
    1.818643, 1.818644, 1.818645, 1.818646, 1.818648, 1.81865, 1.818652, 
    1.818653, 1.818653, 1.818653, 1.818653, 1.818652, 1.818656, 1.818654, 
    1.818657, 1.818657, 1.818655, 1.818657, 1.818643, 1.818642, 1.818641, 
    1.818642, 1.81864, 1.818641, 1.818642, 1.818644, 1.818645, 1.818645, 
    1.818646, 1.818648, 1.81865, 1.818652, 1.818654, 1.818654, 1.818654, 
    1.818654, 1.818653, 1.818654, 1.818654, 1.818654, 1.818657, 1.818656, 
    1.818657, 1.818656, 1.818643, 1.818643, 1.818643, 1.818644, 1.818643, 
    1.818645, 1.818646, 1.818649, 1.818648, 1.81865, 1.818648, 1.818648, 
    1.81865, 1.818648, 1.818652, 1.818649, 1.818654, 1.818651, 1.818654, 
    1.818654, 1.818655, 1.818655, 1.818656, 1.818658, 1.818658, 1.818659, 
    1.818644, 1.818645, 1.818645, 1.818646, 1.818647, 1.818648, 1.818651, 
    1.81865, 1.818651, 1.818652, 1.818649, 1.818651, 1.818646, 1.818647, 
    1.818646, 1.818644, 1.81865, 1.818647, 1.818652, 1.818651, 1.818655, 
    1.818653, 1.818657, 1.818659, 1.818661, 1.818663, 1.818646, 1.818645, 
    1.818646, 1.818648, 1.818649, 1.818651, 1.818651, 1.818651, 1.818652, 
    1.818653, 1.818651, 1.818653, 1.818647, 1.81865, 1.818645, 1.818646, 
    1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 1.818659, 
    1.818655, 1.818665, 1.818662, 1.818645, 1.818646, 1.818648, 1.818647, 
    1.818651, 1.818652, 1.818653, 1.818654, 1.818654, 1.818654, 1.818653, 
    1.818654, 1.818651, 1.818652, 1.818648, 1.818649, 1.818649, 1.818648, 
    1.81865, 1.818651, 1.818652, 1.818652, 1.818654, 1.818651, 1.818659, 
    1.818654, 1.818647, 1.818648, 1.818648, 1.818648, 1.818652, 1.81865, 
    1.818654, 1.818653, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.81865, 1.818649, 1.818648, 1.818648, 1.818649, 1.818652, 1.818654, 
    1.818653, 1.818655, 1.818651, 1.818652, 1.818652, 1.818654, 1.81865, 
    1.818653, 1.818649, 1.818649, 1.81865, 1.818653, 1.818653, 1.818654, 
    1.818653, 1.818652, 1.818651, 1.81865, 1.81865, 1.818649, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818653, 1.818655, 1.818656, 1.818658, 
    1.818656, 1.818659, 1.818657, 1.818661, 1.818653, 1.818657, 1.81865, 
    1.818651, 1.818652, 1.818655, 1.818653, 1.818655, 1.818651, 1.818649, 
    1.818649, 1.818648, 1.818649, 1.818649, 1.81865, 1.818649, 1.818652, 
    1.81865, 1.818654, 1.818655, 1.818659, 1.818661, 1.818663, 1.818664, 
    1.818665, 1.818665,
  1.818617, 1.818619, 1.818619, 1.818621, 1.81862, 1.818621, 1.818618, 
    1.818619, 1.818618, 1.818618, 1.818624, 1.818621, 1.818627, 1.818625, 
    1.81863, 1.818627, 1.818631, 1.81863, 1.818633, 1.818632, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818635, 1.818633, 1.818621, 1.818624, 
    1.818621, 1.818622, 1.818622, 1.81862, 1.818619, 1.818617, 1.818617, 
    1.818619, 1.818622, 1.818621, 1.818623, 1.818623, 1.818626, 1.818625, 
    1.818629, 1.818628, 1.818632, 1.818631, 1.818632, 1.818632, 1.818632, 
    1.81863, 1.818631, 1.81863, 1.818625, 1.818626, 1.818622, 1.81862, 
    1.818618, 1.818617, 1.818617, 1.818617, 1.818619, 1.81862, 1.818622, 
    1.818622, 1.818623, 1.818626, 1.818627, 1.81863, 1.818629, 1.81863, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.81863, 1.818632, 1.818629, 
    1.81863, 1.818623, 1.818621, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818618, 1.818619, 1.81862, 1.81862, 1.818622, 1.818621, 1.818627, 
    1.818624, 1.818631, 1.818629, 1.818631, 1.81863, 1.818632, 1.81863, 
    1.818633, 1.818633, 1.818633, 1.818635, 1.81863, 1.818632, 1.81862, 
    1.81862, 1.81862, 1.818619, 1.818619, 1.818617, 1.818618, 1.818619, 
    1.81862, 1.818621, 1.818622, 1.818623, 1.818625, 1.818628, 1.818629, 
    1.818631, 1.81863, 1.81863, 1.81863, 1.818629, 1.818633, 1.818631, 
    1.818634, 1.818634, 1.818633, 1.818634, 1.81862, 1.818619, 1.818618, 
    1.818619, 1.818617, 1.818618, 1.818619, 1.818621, 1.818622, 1.818622, 
    1.818624, 1.818625, 1.818627, 1.818629, 1.818631, 1.818631, 1.818631, 
    1.818631, 1.81863, 1.818631, 1.818632, 1.818631, 1.818634, 1.818633, 
    1.818634, 1.818634, 1.818619, 1.81862, 1.81862, 1.818621, 1.81862, 
    1.818622, 1.818623, 1.818626, 1.818625, 1.818627, 1.818625, 1.818625, 
    1.818627, 1.818625, 1.818629, 1.818626, 1.818631, 1.818629, 1.818631, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.818635, 1.818635, 1.818636, 
    1.818621, 1.818622, 1.818622, 1.818623, 1.818624, 1.818625, 1.818628, 
    1.818627, 1.818628, 1.818629, 1.818626, 1.818628, 1.818623, 1.818624, 
    1.818623, 1.818621, 1.818627, 1.818624, 1.818629, 1.818628, 1.818632, 
    1.81863, 1.818635, 1.818637, 1.818638, 1.81864, 1.818623, 1.818622, 
    1.818623, 1.818625, 1.818626, 1.818628, 1.818628, 1.818628, 1.818629, 
    1.81863, 1.818629, 1.81863, 1.818624, 1.818627, 1.818622, 1.818623, 
    1.818625, 1.818624, 1.818627, 1.818627, 1.81863, 1.818628, 1.818636, 
    1.818633, 1.818642, 1.818639, 1.818622, 1.818623, 1.818626, 1.818624, 
    1.818628, 1.818629, 1.81863, 1.818631, 1.818631, 1.818632, 1.818631, 
    1.818631, 1.818628, 1.81863, 1.818625, 1.818626, 1.818626, 1.818625, 
    1.818627, 1.818629, 1.818629, 1.818629, 1.818631, 1.818628, 1.818636, 
    1.818631, 1.818624, 1.818625, 1.818625, 1.818625, 1.818629, 1.818627, 
    1.818632, 1.81863, 1.818632, 1.818631, 1.818631, 1.81863, 1.818629, 
    1.818627, 1.818626, 1.818625, 1.818625, 1.818626, 1.818629, 1.818631, 
    1.81863, 1.818632, 1.818628, 1.81863, 1.818629, 1.818631, 1.818627, 
    1.81863, 1.818626, 1.818626, 1.818627, 1.81863, 1.81863, 1.818631, 
    1.81863, 1.818629, 1.818629, 1.818627, 1.818627, 1.818626, 1.818625, 
    1.818626, 1.818627, 1.818629, 1.818631, 1.818632, 1.818633, 1.818635, 
    1.818633, 1.818637, 1.818634, 1.818638, 1.81863, 1.818634, 1.818627, 
    1.818628, 1.818629, 1.818632, 1.818631, 1.818632, 1.818629, 1.818626, 
    1.818626, 1.818625, 1.818626, 1.818626, 1.818627, 1.818627, 1.818629, 
    1.818628, 1.818631, 1.818632, 1.818636, 1.818638, 1.818641, 1.818642, 
    1.818642, 1.818642,
  1.818568, 1.81857, 1.81857, 1.818571, 1.81857, 1.818571, 1.818569, 1.81857, 
    1.818569, 1.818568, 1.818574, 1.818571, 1.818577, 1.818575, 1.81858, 
    1.818577, 1.81858, 1.818579, 1.818581, 1.818581, 1.818583, 1.818582, 
    1.818585, 1.818583, 1.818583, 1.818582, 1.818572, 1.818574, 1.818572, 
    1.818572, 1.818572, 1.81857, 1.81857, 1.818568, 1.818568, 1.818569, 
    1.818572, 1.818571, 1.818573, 1.818573, 1.818576, 1.818575, 1.818579, 
    1.818578, 1.818581, 1.81858, 1.818581, 1.818581, 1.818581, 1.81858, 
    1.81858, 1.818579, 1.818575, 1.818576, 1.818572, 1.81857, 1.818569, 
    1.818568, 1.818568, 1.818568, 1.818569, 1.818571, 1.818572, 1.818573, 
    1.818573, 1.818575, 1.818576, 1.818579, 1.818578, 1.818579, 1.81858, 
    1.818581, 1.818581, 1.818582, 1.818579, 1.818581, 1.818578, 1.818579, 
    1.818573, 1.818571, 1.81857, 1.81857, 1.818568, 1.818569, 1.818569, 
    1.81857, 1.818571, 1.81857, 1.818573, 1.818572, 1.818577, 1.818574, 
    1.81858, 1.818579, 1.81858, 1.818579, 1.818581, 1.81858, 1.818582, 
    1.818582, 1.818582, 1.818583, 1.818579, 1.818581, 1.81857, 1.81857, 
    1.818571, 1.818569, 1.818569, 1.818568, 1.818569, 1.81857, 1.818571, 
    1.818571, 1.818572, 1.818573, 1.818575, 1.818577, 1.818579, 1.81858, 
    1.818579, 1.81858, 1.818579, 1.818579, 1.818582, 1.81858, 1.818583, 
    1.818583, 1.818582, 1.818583, 1.81857, 1.81857, 1.818569, 1.81857, 
    1.818568, 1.818569, 1.818569, 1.818572, 1.818572, 1.818573, 1.818573, 
    1.818575, 1.818577, 1.818578, 1.81858, 1.81858, 1.81858, 1.81858, 
    1.818579, 1.81858, 1.818581, 1.81858, 1.818583, 1.818582, 1.818583, 
    1.818582, 1.81857, 1.818571, 1.81857, 1.818571, 1.81857, 1.818572, 
    1.818573, 1.818576, 1.818575, 1.818576, 1.818575, 1.818575, 1.818576, 
    1.818575, 1.818578, 1.818576, 1.81858, 1.818578, 1.818581, 1.81858, 
    1.818581, 1.818581, 1.818582, 1.818584, 1.818583, 1.818585, 1.818572, 
    1.818572, 1.818572, 1.818573, 1.818574, 1.818575, 1.818577, 1.818576, 
    1.818578, 1.818578, 1.818576, 1.818577, 1.818573, 1.818574, 1.818573, 
    1.818572, 1.818577, 1.818574, 1.818579, 1.818577, 1.818581, 1.818579, 
    1.818583, 1.818585, 1.818586, 1.818588, 1.818573, 1.818572, 1.818573, 
    1.818575, 1.818576, 1.818577, 1.818578, 1.818578, 1.818579, 1.818579, 
    1.818578, 1.81858, 1.818574, 1.818577, 1.818572, 1.818573, 1.818574, 
    1.818574, 1.818576, 1.818577, 1.818579, 1.818578, 1.818584, 1.818582, 
    1.81859, 1.818587, 1.818572, 1.818573, 1.818575, 1.818574, 1.818578, 
    1.818578, 1.818579, 1.81858, 1.81858, 1.818581, 1.81858, 1.818581, 
    1.818577, 1.818579, 1.818575, 1.818576, 1.818576, 1.818575, 1.818576, 
    1.818578, 1.818578, 1.818578, 1.81858, 1.818578, 1.818585, 1.81858, 
    1.818574, 1.818575, 1.818575, 1.818575, 1.818578, 1.818577, 1.818581, 
    1.81858, 1.818581, 1.81858, 1.81858, 1.818579, 1.818579, 1.818577, 
    1.818576, 1.818575, 1.818575, 1.818576, 1.818578, 1.81858, 1.81858, 
    1.818581, 1.818577, 1.818579, 1.818578, 1.81858, 1.818576, 1.818579, 
    1.818576, 1.818576, 1.818577, 1.818579, 1.818579, 1.81858, 1.81858, 
    1.818578, 1.818578, 1.818577, 1.818577, 1.818576, 1.818575, 1.818576, 
    1.818576, 1.818578, 1.81858, 1.818581, 1.818582, 1.818584, 1.818582, 
    1.818585, 1.818583, 1.818587, 1.818579, 1.818583, 1.818577, 1.818578, 
    1.818579, 1.818581, 1.81858, 1.818581, 1.818578, 1.818576, 1.818576, 
    1.818575, 1.818576, 1.818576, 1.818576, 1.818576, 1.818578, 1.818577, 
    1.81858, 1.818581, 1.818585, 1.818587, 1.818589, 1.818589, 1.81859, 
    1.81859,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.293384e-09, 1.299131e-09, 1.298014e-09, 1.30265e-09, 1.300078e-09, 
    1.303114e-09, 1.294549e-09, 1.299359e-09, 1.296289e-09, 1.293902e-09, 
    1.311647e-09, 1.302857e-09, 1.320781e-09, 1.315174e-09, 1.329262e-09, 
    1.319909e-09, 1.331149e-09, 1.328993e-09, 1.335483e-09, 1.333624e-09, 
    1.341925e-09, 1.336341e-09, 1.346229e-09, 1.340592e-09, 1.341473e-09, 
    1.336157e-09, 1.304626e-09, 1.310553e-09, 1.304275e-09, 1.30512e-09, 
    1.304741e-09, 1.300131e-09, 1.297808e-09, 1.292945e-09, 1.293828e-09, 
    1.2974e-09, 1.3055e-09, 1.30275e-09, 1.309681e-09, 1.309524e-09, 
    1.31724e-09, 1.313761e-09, 1.326733e-09, 1.323046e-09, 1.333701e-09, 
    1.331021e-09, 1.333575e-09, 1.332801e-09, 1.333585e-09, 1.329655e-09, 
    1.331339e-09, 1.32788e-09, 1.314413e-09, 1.31837e-09, 1.306568e-09, 
    1.299472e-09, 1.29476e-09, 1.291417e-09, 1.291889e-09, 1.29279e-09, 
    1.297421e-09, 1.301775e-09, 1.305094e-09, 1.307314e-09, 1.309502e-09, 
    1.316123e-09, 1.319628e-09, 1.327478e-09, 1.326062e-09, 1.328461e-09, 
    1.330755e-09, 1.334604e-09, 1.333971e-09, 1.335667e-09, 1.328398e-09, 
    1.333229e-09, 1.325255e-09, 1.327436e-09, 1.310095e-09, 1.303492e-09, 
    1.300685e-09, 1.298229e-09, 1.292253e-09, 1.29638e-09, 1.294753e-09, 
    1.298623e-09, 1.301083e-09, 1.299867e-09, 1.307375e-09, 1.304456e-09, 
    1.319836e-09, 1.313211e-09, 1.330487e-09, 1.326352e-09, 1.331478e-09, 
    1.328863e-09, 1.333344e-09, 1.329311e-09, 1.336298e-09, 1.33782e-09, 
    1.33678e-09, 1.340775e-09, 1.329087e-09, 1.333575e-09, 1.299832e-09, 
    1.300031e-09, 1.300955e-09, 1.296892e-09, 1.296643e-09, 1.292921e-09, 
    1.296233e-09, 1.297644e-09, 1.301226e-09, 1.303344e-09, 1.305358e-09, 
    1.309786e-09, 1.314732e-09, 1.32165e-09, 1.32662e-09, 1.329952e-09, 
    1.327909e-09, 1.329713e-09, 1.327697e-09, 1.326752e-09, 1.33725e-09, 
    1.331354e-09, 1.3402e-09, 1.339711e-09, 1.335707e-09, 1.339766e-09, 
    1.30017e-09, 1.299028e-09, 1.295065e-09, 1.298167e-09, 1.292515e-09, 
    1.295678e-09, 1.297497e-09, 1.304516e-09, 1.306059e-09, 1.307489e-09, 
    1.310314e-09, 1.313939e-09, 1.3203e-09, 1.325834e-09, 1.330888e-09, 
    1.330518e-09, 1.330648e-09, 1.331777e-09, 1.328981e-09, 1.332236e-09, 
    1.332782e-09, 1.331354e-09, 1.339645e-09, 1.337276e-09, 1.3397e-09, 
    1.338158e-09, 1.2994e-09, 1.301321e-09, 1.300283e-09, 1.302235e-09, 
    1.300859e-09, 1.306975e-09, 1.308808e-09, 1.317389e-09, 1.313868e-09, 
    1.319473e-09, 1.314437e-09, 1.315329e-09, 1.319655e-09, 1.314709e-09, 
    1.325529e-09, 1.318193e-09, 1.331821e-09, 1.324494e-09, 1.33228e-09, 
    1.330866e-09, 1.333207e-09, 1.335304e-09, 1.337942e-09, 1.342809e-09, 
    1.341682e-09, 1.345754e-09, 1.304185e-09, 1.306676e-09, 1.306457e-09, 
    1.309065e-09, 1.310994e-09, 1.315175e-09, 1.321882e-09, 1.31936e-09, 
    1.32399e-09, 1.32492e-09, 1.317885e-09, 1.322204e-09, 1.308344e-09, 
    1.310583e-09, 1.30925e-09, 1.304381e-09, 1.31994e-09, 1.311955e-09, 
    1.326703e-09, 1.322376e-09, 1.335005e-09, 1.328723e-09, 1.341062e-09, 
    1.346337e-09, 1.351303e-09, 1.357106e-09, 1.308037e-09, 1.306343e-09, 
    1.309375e-09, 1.31357e-09, 1.317463e-09, 1.322639e-09, 1.323169e-09, 
    1.324139e-09, 1.326651e-09, 1.328763e-09, 1.324445e-09, 1.329292e-09, 
    1.311102e-09, 1.320634e-09, 1.305703e-09, 1.310198e-09, 1.313323e-09, 
    1.311953e-09, 1.319072e-09, 1.32075e-09, 1.327569e-09, 1.324044e-09, 
    1.345035e-09, 1.335747e-09, 1.361526e-09, 1.35432e-09, 1.305752e-09, 
    1.308031e-09, 1.315964e-09, 1.312189e-09, 1.322985e-09, 1.325643e-09, 
    1.327804e-09, 1.330565e-09, 1.330864e-09, 1.3325e-09, 1.329819e-09, 
    1.332394e-09, 1.32265e-09, 1.327005e-09, 1.315057e-09, 1.317965e-09, 
    1.316627e-09, 1.31516e-09, 1.319688e-09, 1.324513e-09, 1.324617e-09, 
    1.326164e-09, 1.330523e-09, 1.323029e-09, 1.346233e-09, 1.331901e-09, 
    1.310516e-09, 1.314906e-09, 1.315534e-09, 1.313833e-09, 1.325376e-09, 
    1.321193e-09, 1.33246e-09, 1.329415e-09, 1.334405e-09, 1.331925e-09, 
    1.331561e-09, 1.328376e-09, 1.326394e-09, 1.321385e-09, 1.31731e-09, 
    1.31408e-09, 1.314831e-09, 1.31838e-09, 1.324808e-09, 1.330891e-09, 
    1.329558e-09, 1.334026e-09, 1.322202e-09, 1.32716e-09, 1.325243e-09, 
    1.33024e-09, 1.319293e-09, 1.328614e-09, 1.31691e-09, 1.317936e-09, 
    1.32111e-09, 1.327496e-09, 1.328909e-09, 1.330417e-09, 1.329487e-09, 
    1.324972e-09, 1.324232e-09, 1.321033e-09, 1.32015e-09, 1.317713e-09, 
    1.315695e-09, 1.317539e-09, 1.319475e-09, 1.324974e-09, 1.32993e-09, 
    1.335334e-09, 1.336656e-09, 1.342971e-09, 1.33783e-09, 1.346313e-09, 
    1.3391e-09, 1.351587e-09, 1.329155e-09, 1.338889e-09, 1.321255e-09, 
    1.323154e-09, 1.32659e-09, 1.334471e-09, 1.330216e-09, 1.335192e-09, 
    1.324203e-09, 1.318502e-09, 1.317028e-09, 1.314276e-09, 1.317091e-09, 
    1.316862e-09, 1.319555e-09, 1.318689e-09, 1.325156e-09, 1.321683e-09, 
    1.331551e-09, 1.335153e-09, 1.345327e-09, 1.351564e-09, 1.357915e-09, 
    1.360719e-09, 1.361572e-09, 1.361929e-09 ;

 SOIL2_HR_S3 =
  9.238458e-11, 9.279509e-11, 9.271529e-11, 9.304642e-11, 9.286274e-11, 
    9.307956e-11, 9.246781e-11, 9.281138e-11, 9.259205e-11, 9.242154e-11, 
    9.368908e-11, 9.30612e-11, 9.434153e-11, 9.394097e-11, 9.494731e-11, 
    9.42792e-11, 9.508206e-11, 9.492807e-11, 9.539163e-11, 9.525882e-11, 
    9.585177e-11, 9.545294e-11, 9.615922e-11, 9.575653e-11, 9.581951e-11, 
    9.543977e-11, 9.318757e-11, 9.36109e-11, 9.316248e-11, 9.322285e-11, 
    9.319576e-11, 9.286653e-11, 9.27006e-11, 9.235322e-11, 9.241628e-11, 
    9.267144e-11, 9.324999e-11, 9.305361e-11, 9.354861e-11, 9.353743e-11, 
    9.40886e-11, 9.384008e-11, 9.476662e-11, 9.450326e-11, 9.526437e-11, 
    9.507294e-11, 9.525537e-11, 9.520006e-11, 9.525609e-11, 9.497535e-11, 
    9.509563e-11, 9.48486e-11, 9.388661e-11, 9.41693e-11, 9.332626e-11, 
    9.281943e-11, 9.248287e-11, 9.224406e-11, 9.227782e-11, 9.234218e-11, 
    9.267294e-11, 9.298396e-11, 9.322101e-11, 9.337957e-11, 9.353583e-11, 
    9.400877e-11, 9.425917e-11, 9.481986e-11, 9.471869e-11, 9.48901e-11, 
    9.50539e-11, 9.532888e-11, 9.528362e-11, 9.540477e-11, 9.48856e-11, 
    9.523063e-11, 9.466106e-11, 9.481683e-11, 9.357824e-11, 9.310659e-11, 
    9.290607e-11, 9.273063e-11, 9.230378e-11, 9.259854e-11, 9.248233e-11, 
    9.275881e-11, 9.293449e-11, 9.284761e-11, 9.338391e-11, 9.31754e-11, 
    9.427401e-11, 9.380076e-11, 9.503479e-11, 9.473946e-11, 9.510558e-11, 
    9.491876e-11, 9.523888e-11, 9.495078e-11, 9.544987e-11, 9.555855e-11, 
    9.548428e-11, 9.576961e-11, 9.49348e-11, 9.525537e-11, 9.284517e-11, 
    9.285934e-11, 9.292536e-11, 9.263515e-11, 9.261739e-11, 9.235148e-11, 
    9.25881e-11, 9.268886e-11, 9.294469e-11, 9.3096e-11, 9.323986e-11, 
    9.355617e-11, 9.390946e-11, 9.440356e-11, 9.47586e-11, 9.49966e-11, 
    9.485067e-11, 9.497951e-11, 9.483547e-11, 9.476797e-11, 9.551782e-11, 
    9.509675e-11, 9.572857e-11, 9.569361e-11, 9.540765e-11, 9.569755e-11, 
    9.286929e-11, 9.278775e-11, 9.250462e-11, 9.272619e-11, 9.232252e-11, 
    9.254846e-11, 9.267838e-11, 9.317973e-11, 9.328992e-11, 9.339207e-11, 
    9.359385e-11, 9.38528e-11, 9.430712e-11, 9.470246e-11, 9.506343e-11, 
    9.503698e-11, 9.504629e-11, 9.512693e-11, 9.492718e-11, 9.515971e-11, 
    9.519874e-11, 9.50967e-11, 9.568893e-11, 9.551972e-11, 9.569287e-11, 
    9.55827e-11, 9.281426e-11, 9.295147e-11, 9.287732e-11, 9.301675e-11, 
    9.291852e-11, 9.335532e-11, 9.34863e-11, 9.409924e-11, 9.38477e-11, 
    9.424807e-11, 9.388837e-11, 9.39521e-11, 9.426111e-11, 9.390781e-11, 
    9.468065e-11, 9.415665e-11, 9.513006e-11, 9.460669e-11, 9.516286e-11, 
    9.506187e-11, 9.522908e-11, 9.537884e-11, 9.556728e-11, 9.591496e-11, 
    9.583445e-11, 9.612525e-11, 9.315605e-11, 9.333403e-11, 9.331837e-11, 
    9.350466e-11, 9.364243e-11, 9.394108e-11, 9.442012e-11, 9.423998e-11, 
    9.457071e-11, 9.463711e-11, 9.413465e-11, 9.444313e-11, 9.345318e-11, 
    9.361308e-11, 9.351788e-11, 9.317008e-11, 9.428146e-11, 9.371105e-11, 
    9.476447e-11, 9.445539e-11, 9.535749e-11, 9.490882e-11, 9.579013e-11, 
    9.616691e-11, 9.652164e-11, 9.693614e-11, 9.343119e-11, 9.331025e-11, 
    9.352683e-11, 9.382645e-11, 9.410454e-11, 9.447424e-11, 9.451208e-11, 
    9.458134e-11, 9.476078e-11, 9.491163e-11, 9.460323e-11, 9.494946e-11, 
    9.365014e-11, 9.433099e-11, 9.326451e-11, 9.35856e-11, 9.38088e-11, 
    9.37109e-11, 9.42194e-11, 9.433924e-11, 9.482633e-11, 9.457454e-11, 
    9.60739e-11, 9.541046e-11, 9.725182e-11, 9.673714e-11, 9.326799e-11, 
    9.343078e-11, 9.399741e-11, 9.37278e-11, 9.449893e-11, 9.468876e-11, 
    9.484311e-11, 9.504039e-11, 9.50617e-11, 9.517859e-11, 9.498704e-11, 
    9.517103e-11, 9.447503e-11, 9.478604e-11, 9.393265e-11, 9.414033e-11, 
    9.404479e-11, 9.393999e-11, 9.426346e-11, 9.460808e-11, 9.461547e-11, 
    9.472597e-11, 9.503735e-11, 9.450207e-11, 9.61595e-11, 9.513578e-11, 
    9.360832e-11, 9.392188e-11, 9.396671e-11, 9.384523e-11, 9.466973e-11, 
    9.437096e-11, 9.517575e-11, 9.495823e-11, 9.531465e-11, 9.513753e-11, 
    9.511147e-11, 9.488401e-11, 9.474239e-11, 9.438465e-11, 9.409361e-11, 
    9.386285e-11, 9.391651e-11, 9.417e-11, 9.462917e-11, 9.506362e-11, 
    9.496844e-11, 9.528756e-11, 9.444302e-11, 9.479711e-11, 9.466024e-11, 
    9.501714e-11, 9.42352e-11, 9.490098e-11, 9.406502e-11, 9.413831e-11, 
    9.436503e-11, 9.482111e-11, 9.492206e-11, 9.50298e-11, 9.496332e-11, 
    9.464083e-11, 9.4588e-11, 9.435952e-11, 9.429642e-11, 9.412236e-11, 
    9.397823e-11, 9.410991e-11, 9.424819e-11, 9.464097e-11, 9.499498e-11, 
    9.538097e-11, 9.547545e-11, 9.592647e-11, 9.555929e-11, 9.616519e-11, 
    9.565002e-11, 9.654191e-11, 9.493961e-11, 9.56349e-11, 9.437535e-11, 
    9.451103e-11, 9.475642e-11, 9.531936e-11, 9.501546e-11, 9.537088e-11, 
    9.458594e-11, 9.417873e-11, 9.407341e-11, 9.387688e-11, 9.407791e-11, 
    9.406156e-11, 9.425393e-11, 9.419211e-11, 9.465401e-11, 9.440589e-11, 
    9.511082e-11, 9.536808e-11, 9.609476e-11, 9.65403e-11, 9.699393e-11, 
    9.719421e-11, 9.725518e-11, 9.728066e-11 ;

 SOIL3C =
  5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611 ;

 SOIL3C_TO_SOIL1C =
  2.55052e-11, 2.561851e-11, 2.559648e-11, 2.568788e-11, 2.563718e-11, 
    2.569703e-11, 2.552817e-11, 2.5623e-11, 2.556247e-11, 2.55154e-11, 
    2.586527e-11, 2.569196e-11, 2.604535e-11, 2.593479e-11, 2.621256e-11, 
    2.602814e-11, 2.624975e-11, 2.620724e-11, 2.633519e-11, 2.629854e-11, 
    2.64622e-11, 2.635211e-11, 2.654706e-11, 2.643591e-11, 2.64533e-11, 
    2.634848e-11, 2.572684e-11, 2.584369e-11, 2.571991e-11, 2.573658e-11, 
    2.57291e-11, 2.563823e-11, 2.559243e-11, 2.549654e-11, 2.551395e-11, 
    2.558438e-11, 2.574407e-11, 2.568986e-11, 2.582649e-11, 2.582341e-11, 
    2.597554e-11, 2.590694e-11, 2.616268e-11, 2.608999e-11, 2.630007e-11, 
    2.624723e-11, 2.629759e-11, 2.628232e-11, 2.629778e-11, 2.622029e-11, 
    2.625349e-11, 2.618531e-11, 2.591979e-11, 2.599781e-11, 2.576512e-11, 
    2.562523e-11, 2.553233e-11, 2.546641e-11, 2.547573e-11, 2.549349e-11, 
    2.558479e-11, 2.567064e-11, 2.573607e-11, 2.577984e-11, 2.582297e-11, 
    2.59535e-11, 2.602262e-11, 2.617738e-11, 2.614945e-11, 2.619677e-11, 
    2.624197e-11, 2.631787e-11, 2.630538e-11, 2.633882e-11, 2.619552e-11, 
    2.629075e-11, 2.613354e-11, 2.617654e-11, 2.583467e-11, 2.570449e-11, 
    2.564914e-11, 2.560072e-11, 2.54829e-11, 2.556426e-11, 2.553218e-11, 
    2.560849e-11, 2.565699e-11, 2.5633e-11, 2.578103e-11, 2.572348e-11, 
    2.602671e-11, 2.589609e-11, 2.62367e-11, 2.615518e-11, 2.625624e-11, 
    2.620467e-11, 2.629303e-11, 2.621351e-11, 2.635127e-11, 2.638127e-11, 
    2.636077e-11, 2.643952e-11, 2.62091e-11, 2.629758e-11, 2.563233e-11, 
    2.563624e-11, 2.565446e-11, 2.557436e-11, 2.556946e-11, 2.549607e-11, 
    2.556137e-11, 2.558919e-11, 2.56598e-11, 2.570156e-11, 2.574127e-11, 
    2.582858e-11, 2.592609e-11, 2.606247e-11, 2.616047e-11, 2.622616e-11, 
    2.618588e-11, 2.622144e-11, 2.618169e-11, 2.616306e-11, 2.637002e-11, 
    2.62538e-11, 2.642819e-11, 2.641854e-11, 2.633962e-11, 2.641963e-11, 
    2.563899e-11, 2.561648e-11, 2.553833e-11, 2.559949e-11, 2.548807e-11, 
    2.555044e-11, 2.558629e-11, 2.572468e-11, 2.575509e-11, 2.578329e-11, 
    2.583898e-11, 2.591045e-11, 2.603585e-11, 2.614497e-11, 2.624461e-11, 
    2.62373e-11, 2.623987e-11, 2.626213e-11, 2.6207e-11, 2.627118e-11, 
    2.628195e-11, 2.625379e-11, 2.641725e-11, 2.637055e-11, 2.641834e-11, 
    2.638793e-11, 2.56238e-11, 2.566167e-11, 2.564121e-11, 2.567969e-11, 
    2.565258e-11, 2.577314e-11, 2.580929e-11, 2.597848e-11, 2.590905e-11, 
    2.601955e-11, 2.592027e-11, 2.593786e-11, 2.602315e-11, 2.592564e-11, 
    2.613895e-11, 2.599432e-11, 2.6263e-11, 2.611854e-11, 2.627205e-11, 
    2.624418e-11, 2.629033e-11, 2.633166e-11, 2.638367e-11, 2.647964e-11, 
    2.645742e-11, 2.653768e-11, 2.571814e-11, 2.576727e-11, 2.576294e-11, 
    2.581436e-11, 2.585239e-11, 2.593482e-11, 2.606704e-11, 2.601732e-11, 
    2.610861e-11, 2.612693e-11, 2.598825e-11, 2.607339e-11, 2.580015e-11, 
    2.584429e-11, 2.581801e-11, 2.572201e-11, 2.602877e-11, 2.587133e-11, 
    2.616209e-11, 2.607678e-11, 2.632577e-11, 2.620193e-11, 2.644518e-11, 
    2.654918e-11, 2.664709e-11, 2.67615e-11, 2.579408e-11, 2.57607e-11, 
    2.582048e-11, 2.590318e-11, 2.597994e-11, 2.608198e-11, 2.609243e-11, 
    2.611154e-11, 2.616107e-11, 2.620271e-11, 2.611758e-11, 2.621315e-11, 
    2.585452e-11, 2.604244e-11, 2.574808e-11, 2.58367e-11, 2.589831e-11, 
    2.587129e-11, 2.601164e-11, 2.604472e-11, 2.617916e-11, 2.610966e-11, 
    2.652351e-11, 2.634039e-11, 2.684863e-11, 2.670657e-11, 2.574904e-11, 
    2.579397e-11, 2.595037e-11, 2.587595e-11, 2.60888e-11, 2.614119e-11, 
    2.618379e-11, 2.623825e-11, 2.624413e-11, 2.627639e-11, 2.622352e-11, 
    2.627431e-11, 2.60822e-11, 2.616804e-11, 2.593249e-11, 2.598982e-11, 
    2.596345e-11, 2.593452e-11, 2.60238e-11, 2.611892e-11, 2.612096e-11, 
    2.615146e-11, 2.623741e-11, 2.608966e-11, 2.654713e-11, 2.626458e-11, 
    2.584297e-11, 2.592952e-11, 2.594189e-11, 2.590836e-11, 2.613594e-11, 
    2.605347e-11, 2.627561e-11, 2.621557e-11, 2.631394e-11, 2.626506e-11, 
    2.625787e-11, 2.619508e-11, 2.6156e-11, 2.605725e-11, 2.597692e-11, 
    2.591323e-11, 2.592804e-11, 2.5998e-11, 2.612474e-11, 2.624466e-11, 
    2.621839e-11, 2.630647e-11, 2.607336e-11, 2.61711e-11, 2.613332e-11, 
    2.623183e-11, 2.6016e-11, 2.619977e-11, 2.596903e-11, 2.598926e-11, 
    2.605184e-11, 2.617772e-11, 2.620559e-11, 2.623532e-11, 2.621697e-11, 
    2.612796e-11, 2.611338e-11, 2.605032e-11, 2.60329e-11, 2.598485e-11, 
    2.594508e-11, 2.598142e-11, 2.601959e-11, 2.6128e-11, 2.622571e-11, 
    2.633225e-11, 2.635833e-11, 2.648282e-11, 2.638147e-11, 2.654871e-11, 
    2.640651e-11, 2.665269e-11, 2.621043e-11, 2.640234e-11, 2.605469e-11, 
    2.609214e-11, 2.615987e-11, 2.631525e-11, 2.623137e-11, 2.632947e-11, 
    2.611281e-11, 2.600042e-11, 2.597134e-11, 2.59171e-11, 2.597259e-11, 
    2.596807e-11, 2.602117e-11, 2.600411e-11, 2.61316e-11, 2.606312e-11, 
    2.625768e-11, 2.632869e-11, 2.652927e-11, 2.665224e-11, 2.677745e-11, 
    2.683273e-11, 2.684956e-11, 2.685659e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  1.003089e-36, -2.055969e-20, -1.003089e-36, -2.569961e-21, -1.798972e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 
    -1.28498e-20, -1.027984e-20, -1.798972e-20, 7.709882e-21, -2.312965e-20, 
    7.709882e-21, 2.569961e-21, 1.027984e-20, -1.28498e-20, 2.569961e-21, 
    7.709882e-21, 1.003089e-36, -7.709882e-21, 0, -5.139921e-21, 
    -1.28498e-20, 1.28498e-20, -1.027984e-20, -7.709882e-21, 1.798972e-20, 
    -5.139921e-21, 1.003089e-36, -5.139921e-21, 5.139921e-21, -1.541976e-20, 
    -2.569961e-21, -1.541976e-20, 7.709882e-21, -1.027984e-20, -1.28498e-20, 
    2.569961e-21, -7.709882e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 7.709882e-21, -1.027984e-20, 1.003089e-36, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, -7.709882e-21, -2.312965e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -2.569961e-21, 1.027984e-20, 5.139921e-21, 1.027984e-20, 1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -1.798972e-20, 1.027984e-20, 
    1.027984e-20, -1.003089e-36, -1.28498e-20, -1.003089e-36, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 
    -1.541976e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -1.003089e-36, -2.569961e-21, -2.569961e-21, -1.027984e-20, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, 2.055969e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 0, -1.541976e-20, -2.569961e-21, 
    5.139921e-21, 1.003089e-36, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -1.027984e-20, -1.541976e-20, -1.798972e-20, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, 1.798972e-20, 5.139921e-21, 
    1.027984e-20, 0, 2.569961e-21, 0, 2.569961e-21, -3.083953e-20, 
    -7.709882e-21, 5.139921e-21, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -1.28498e-20, 1.28498e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 1.003089e-36, -1.541976e-20, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, 1.003089e-36, 
    1.28498e-20, 2.569961e-21, 1.027984e-20, -1.027984e-20, 1.28498e-20, 
    -2.569961e-21, -1.28498e-20, -1.541976e-20, 1.28498e-20, -1.798972e-20, 
    -1.798972e-20, 1.003089e-36, 5.139921e-21, -7.709882e-21, 1.541976e-20, 
    7.709882e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, -1.28498e-20, 
    -1.541976e-20, 5.139921e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    1.28498e-20, 2.569961e-21, -5.139921e-21, 1.541976e-20, -7.709882e-21, 
    1.541976e-20, 2.569961e-21, 2.569961e-21, -1.027984e-20, 7.709882e-21, 
    1.28498e-20, 1.541976e-20, 3.083953e-20, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 1.28498e-20, 1.027984e-20, -1.28498e-20, -2.569961e-21, 
    -1.027984e-20, -1.003089e-36, 1.027984e-20, -1.541976e-20, 7.709882e-21, 
    -2.569961e-21, -1.798972e-20, 7.709882e-21, -7.709882e-21, -1.28498e-20, 
    -1.541976e-20, 1.28498e-20, -1.027984e-20, -2.312965e-20, 5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -1.28498e-20, 0, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    1.003089e-36, -1.027984e-20, 7.709882e-21, 2.569961e-21, -1.541976e-20, 
    -1.027984e-20, 2.055969e-20, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 1.541976e-20, 
    -1.798972e-20, 5.139921e-21, 1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, -1.541976e-20, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -1.541976e-20, 7.709882e-21, 1.003089e-36, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, -1.28498e-20, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 1.28498e-20, 1.003089e-36, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -1.541976e-20, 1.28498e-20, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 1.003089e-36, 1.027984e-20, 1.003089e-36, 2.826957e-20, 
    -2.569961e-21, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 
    1.003089e-36, -1.027984e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -1.027984e-20, -1.28498e-20, -7.709882e-21, 7.709882e-21, 0, 
    1.003089e-36, 1.28498e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, -1.003089e-36, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, 2.569961e-21,
  2.569961e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 0, -5.139921e-21, 
    5.139921e-21, 0, -1.28498e-20, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, 2.569961e-21, 1.003089e-36, -5.139921e-21, 
    1.027984e-20, -7.709882e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, 0, 0, -1.003089e-36, -5.139921e-21, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 0, 
    -1.027984e-20, 0, 0, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, 0, 5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, 2.569961e-21, -1.28498e-20, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, -7.709882e-21, 2.569961e-21, 1.003089e-36, 2.569961e-21, 
    -1.28498e-20, 0, -1.003089e-36, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 7.709882e-21, 0, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, 1.798972e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, -1.027984e-20, 2.569961e-21, -1.541976e-20, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, 1.027984e-20, 0, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -1.027984e-20, 1.027984e-20, 1.28498e-20, -1.798972e-20, -7.709882e-21, 
    -1.28498e-20, -5.139921e-21, -7.709882e-21, 0, -5.139921e-21, 0, 
    -7.709882e-21, -5.139921e-21, 1.28498e-20, -2.569961e-21, 1.28498e-20, 
    2.569961e-21, -2.569961e-21, -1.541976e-20, -2.569961e-21, 0, 0, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -1.003089e-36, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 0, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 0, 5.139921e-21, 
    5.139921e-21, -1.798972e-20, 5.139921e-21, 1.541976e-20, 0, 
    -5.139921e-21, 0, 0, -7.709882e-21, 2.569961e-21, -1.003089e-36, 
    -1.541976e-20, -7.709882e-21, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 0, 2.569961e-21, -5.139921e-21, 1.28498e-20, 7.709882e-21, 
    -7.709882e-21, -1.541976e-20, 0, 1.28498e-20, 1.027984e-20, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, 1.28498e-20, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 7.709882e-21, 1.003089e-36, -7.709882e-21, 0, 0, 
    2.569961e-21, 1.798972e-20, -1.003089e-36, -1.027984e-20, 2.569961e-21, 
    1.027984e-20, -1.28498e-20, 7.709882e-21, 0, -1.541976e-20, 5.139921e-21, 
    -1.027984e-20, -1.003089e-36, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 1.003089e-36, -1.027984e-20, 0, 
    5.139921e-21, 0, -1.027984e-20, -5.139921e-21, 0, -5.139921e-21, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, -7.709882e-21, 1.003089e-36, 
    7.709882e-21, -5.139921e-21, -1.28498e-20, -1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 1.541976e-20, 2.569961e-21, 
    5.139921e-21, -1.28498e-20, 0, -1.027984e-20, -2.569961e-21, 1.28498e-20, 
    -1.003089e-36, 1.027984e-20, -2.569961e-21, -1.541976e-20, -7.709882e-21, 
    0, 0, 7.709882e-21, 2.569961e-21, -7.709882e-21, 2.312965e-20, 
    1.027984e-20, -1.28498e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    0, -7.709882e-21, -1.027984e-20, 1.003089e-36, -7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 0, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.003089e-36, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -1.28498e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 0, -2.569961e-21, 2.055969e-20, 
    5.139921e-21, 7.709882e-21, 1.541976e-20, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -2.055969e-20, 5.139921e-21, 0, 
    5.139921e-21, -1.28498e-20, -7.709882e-21, -1.28498e-20, 5.139921e-21, 
    1.003089e-36,
  -2.569961e-21, 1.027984e-20, 2.569961e-21, 7.709882e-21, 1.28498e-20, 
    2.569961e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, -1.003089e-36, 
    0, -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 0, 
    1.798972e-20, 1.027984e-20, -2.312965e-20, 7.709882e-21, 1.798972e-20, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    1.027984e-20, -1.027984e-20, 1.541976e-20, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    -2.569961e-21, -2.055969e-20, -2.569961e-21, -1.003089e-36, 
    -1.003089e-36, -5.139921e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -1.798972e-20, 1.027984e-20, -7.709882e-21, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, -1.003089e-36, -1.003089e-36, 0, 1.003089e-36, 
    7.709882e-21, 1.541976e-20, -7.709882e-21, 2.569961e-21, 1.027984e-20, 
    -7.709882e-21, -1.003089e-36, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.003089e-36, 0, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    0, 2.055969e-20, 0, -7.709882e-21, 1.798972e-20, -1.798972e-20, 
    -7.709882e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.541976e-20, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, 1.541976e-20, 5.139921e-21, 
    2.569961e-21, 0, 5.139921e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, 0, 2.569961e-21, 1.027984e-20, 1.027984e-20, 
    2.569961e-21, 1.28498e-20, 7.709882e-21, 5.139921e-21, 1.003089e-36, 
    7.709882e-21, -2.569961e-21, -1.798972e-20, -1.28498e-20, 1.28498e-20, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, 0, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 1.28498e-20, -1.003089e-36, -2.569961e-21, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 7.709882e-21, -1.28498e-20, 
    -2.569961e-21, -1.28498e-20, 0, 0, 5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -2.569961e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    -1.798972e-20, 1.003089e-36, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    7.709882e-21, 5.139921e-21, 1.027984e-20, -7.709882e-21, 1.28498e-20, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    7.709882e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 0, 
    1.027984e-20, -7.709882e-21, 1.003089e-36, 1.003089e-36, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -2.569961e-21, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, -1.003089e-36, 5.139921e-21, 1.541976e-20, 
    -2.569961e-21, 1.003089e-36, -1.541976e-20, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 1.027984e-20, 1.027984e-20, 7.709882e-21, 
    -7.709882e-21, 1.28498e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, 2.569961e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, 0, 1.28498e-20, 
    -2.055969e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.541976e-20, 1.28498e-20, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    2.569961e-21, -7.709882e-21, -1.28498e-20, 2.569961e-21, 1.28498e-20, 
    -1.798972e-20, -7.709882e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, 0, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -1.003089e-36, -5.139921e-21, -1.541976e-20, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    5.139921e-21, 1.28498e-20, -7.709882e-21, 2.569961e-21, 0, -1.541976e-20, 
    0, -2.569961e-21, -2.312965e-20, -2.569961e-21, -1.003089e-36, 
    5.139921e-21, -1.027984e-20, -1.003089e-36, 0, -5.139921e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 1.541976e-20, -2.569961e-21, 
    -2.569961e-21, 0, 1.003089e-36, -1.003089e-36, 0, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 0,
  0, -2.569961e-21, -1.027984e-20, -1.28498e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    1.28498e-20, 1.003089e-36, -2.569961e-21, 5.139921e-21, -1.28498e-20, 
    -5.139921e-21, -1.28498e-20, 2.569961e-21, -1.003089e-36, 1.28498e-20, 
    2.569961e-21, 1.28498e-20, 0, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    7.709882e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -1.541976e-20, -2.569961e-21, 
    -1.541976e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.28498e-20, -2.569961e-21, 1.003089e-36, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 0, 
    1.28498e-20, 7.709882e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, 
    1.027984e-20, 5.139921e-21, 1.28498e-20, 2.569961e-21, -1.003089e-36, 
    2.569961e-21, 1.28498e-20, -7.709882e-21, 2.569961e-21, 7.709882e-21, 
    -1.28498e-20, 1.28498e-20, -2.569961e-21, 1.027984e-20, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -1.003089e-36, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, -1.027984e-20, 
    -1.003089e-36, 1.541976e-20, -2.569961e-20, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 2.055969e-20, 
    -7.709882e-21, -2.569961e-21, 1.541976e-20, 0, 0, 2.569961e-21, 
    -7.709882e-21, -1.541976e-20, -1.027984e-20, -1.28498e-20, -1.28498e-20, 
    5.139921e-21, 1.027984e-20, -1.28498e-20, 2.569961e-21, 2.569961e-21, 0, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -1.541976e-20, -1.28498e-20, 5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -1.027984e-20, -1.798972e-20, 2.055969e-20, -1.28498e-20, -1.28498e-20, 
    1.541976e-20, -2.569961e-21, -1.541976e-20, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 1.28498e-20, 1.003089e-36, 1.541976e-20, -2.312965e-20, 
    1.003089e-36, -1.541976e-20, 2.569961e-21, -1.027984e-20, 7.709882e-21, 
    0, -2.569961e-21, 0, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, 1.798972e-20, -1.541976e-20, 2.312965e-20, -1.28498e-20, 
    2.569961e-21, 0, 2.569961e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, -2.569961e-20, 
    3.009266e-36, 5.139921e-21, 1.003089e-36, 1.541976e-20, -2.569961e-21, 
    -1.28498e-20, -1.027984e-20, -2.312965e-20, -2.569961e-21, -1.798972e-20, 
    1.027984e-20, -7.709882e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, 1.003089e-36, 2.569961e-21, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, 7.709882e-21, 1.003089e-36, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, 2.569961e-21, 1.541976e-20, 2.312965e-20, -5.139921e-21, 
    -2.055969e-20, -2.055969e-20, -1.541976e-20, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, -5.139921e-21, 
    1.541976e-20, -7.709882e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 1.003089e-36, 5.139921e-21, 1.798972e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -1.504633e-36, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, 0, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 1.541976e-20, -1.027984e-20, 2.569961e-21, 
    0, 0, 0, -1.003089e-36, 1.003089e-36, -2.569961e-21, 1.541976e-20, 
    1.027984e-20, 5.015443e-37, 0, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.28498e-20, -7.709882e-21, -1.541976e-20, 0, 5.139921e-21, 
    -2.569961e-21, -1.541976e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    7.709882e-21, -1.003089e-36, 1.027984e-20, 1.28498e-20, 1.28498e-20, 
    1.003089e-36, -5.139921e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, 7.709882e-21, -1.027984e-20, -1.798972e-20, 1.027984e-20, 
    1.28498e-20, 1.798972e-20, -2.312965e-20, 5.139921e-21, 7.709882e-21, 0, 
    -1.027984e-20, 7.709882e-21, 0, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 
    0, -2.569961e-21, -1.28498e-20, 2.055969e-20, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 1.541976e-20,
  2.569961e-21, 5.139921e-21, 1.28498e-20, -1.027984e-20, -2.569961e-21, 
    1.28498e-20, -5.139921e-21, 1.28498e-20, 2.569961e-20, -2.569961e-21, 
    -2.055969e-20, 7.709882e-21, -2.569961e-20, -1.28498e-20, -1.28498e-20, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    0, -1.027984e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    1.798972e-20, 5.139921e-21, -2.569961e-21, 2.569961e-21, 1.28498e-20, 
    -1.027984e-20, -2.569961e-21, 2.569961e-21, -1.027984e-20, 0, 
    5.139921e-21, -5.139921e-21, 7.709882e-21, 1.28498e-20, -5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 1.003089e-36, -1.027984e-20, -2.569961e-21, 
    -1.027984e-20, 1.003089e-36, 7.709882e-21, -7.709882e-21, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, -1.28498e-20, 0, 5.139921e-21, 1.798972e-20, 
    1.28498e-20, 1.541976e-20, -1.027984e-20, -7.709882e-21, 1.541976e-20, 
    -1.28498e-20, 1.027984e-20, -2.569961e-21, -7.709882e-21, 0, 
    1.541976e-20, 5.139921e-21, 2.569961e-21, 0, -2.312965e-20, 
    -2.569961e-21, -1.027984e-20, 1.027984e-20, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, -1.027984e-20, -1.027984e-20, -1.541976e-20, 7.709882e-21, 
    1.541976e-20, -2.312965e-20, -1.003089e-36, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, 1.541976e-20, 2.569961e-21, 5.139921e-21, 1.28498e-20, 
    2.569961e-20, 7.709882e-21, 2.569961e-21, -1.027984e-20, -5.139921e-21, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 1.003089e-36, 
    -1.28498e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 1.541976e-20, 
    2.055969e-20, -1.798972e-20, 1.027984e-20, 1.541976e-20, 2.569961e-21, 
    -2.055969e-20, -1.027984e-20, 7.709882e-21, 5.139921e-21, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 0, -1.541976e-20, 
    1.541976e-20, -1.28498e-20, -1.003089e-36, -1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, 1.28498e-20, -1.541976e-20, 
    -5.139921e-21, 0, -7.709882e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, -1.541976e-20, 1.027984e-20, 1.28498e-20, 1.28498e-20, 
    2.055969e-20, 1.28498e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, -2.055969e-20, 2.055969e-20, 
    7.709882e-21, -1.798972e-20, 0, 5.139921e-21, 7.709882e-21, 0, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 1.798972e-20, 
    1.541976e-20, -2.569961e-21, -1.798972e-20, 2.569961e-21, 0, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.28498e-20, 2.055969e-20, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, 1.798972e-20, 1.027984e-20, 
    -1.28498e-20, -1.027984e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -1.003089e-36, -7.709882e-21, 2.055969e-20, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    1.798972e-20, 5.139921e-21, -7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, 1.28498e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 1.798972e-20, -1.027984e-20, -1.027984e-20, -2.569961e-21, 
    -1.027984e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    1.798972e-20, -1.798972e-20, 0, -1.28498e-20, 0, -1.798972e-20, 
    -1.027984e-20, -2.569961e-21, 1.541976e-20, 5.139921e-21, 0, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 1.003089e-36, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -1.541976e-20, -1.027984e-20, 7.709882e-21, 
    1.003089e-36, 7.709882e-21, 1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -7.709882e-21, -1.003089e-36, 7.709882e-21, 2.312965e-20, 1.541976e-20, 
    -1.027984e-20, 2.569961e-21, 1.003089e-36, 1.798972e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    0, -2.569961e-21, 2.055969e-20, -1.003089e-36, 1.798972e-20, 
    -1.541976e-20, -1.027984e-20, -5.139921e-21, 1.798972e-20, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 1.28498e-20, 1.027984e-20, 
    1.541976e-20, -1.541976e-20, 1.541976e-20, -7.709882e-21, -5.139921e-21, 
    7.709882e-21, 1.027984e-20, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, -1.798972e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, -1.003089e-36, 1.541976e-20, 
    5.139921e-21, -2.312965e-20, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    0, -5.139921e-21, 2.569961e-21, -2.312965e-20, -2.312965e-20, 
    1.003089e-36, -2.312965e-20, 0, -5.139921e-21, -5.139921e-21, 
    2.569961e-20, -1.003089e-36, 5.139921e-21, 1.541976e-20, 2.569961e-21, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, -1.28498e-20, -1.003089e-36, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -1.541976e-20, 1.003089e-36, 5.139921e-21, 
    -2.312965e-20, -1.798972e-20, 0, 1.027984e-20, -7.709882e-21,
  6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.152565e-12, 5.175456e-12, 5.171006e-12, 5.18947e-12, 5.179229e-12, 
    5.191318e-12, 5.157207e-12, 5.176365e-12, 5.164135e-12, 5.154627e-12, 
    5.225306e-12, 5.190295e-12, 5.261687e-12, 5.239352e-12, 5.295466e-12, 
    5.258211e-12, 5.302979e-12, 5.294393e-12, 5.320241e-12, 5.312836e-12, 
    5.345899e-12, 5.323659e-12, 5.363042e-12, 5.340589e-12, 5.3441e-12, 
    5.322926e-12, 5.197341e-12, 5.220947e-12, 5.195942e-12, 5.199308e-12, 
    5.197798e-12, 5.179439e-12, 5.170188e-12, 5.150817e-12, 5.154334e-12, 
    5.168561e-12, 5.200822e-12, 5.189871e-12, 5.217474e-12, 5.21685e-12, 
    5.247584e-12, 5.233726e-12, 5.28539e-12, 5.270705e-12, 5.313145e-12, 
    5.302471e-12, 5.312644e-12, 5.309559e-12, 5.312683e-12, 5.297029e-12, 
    5.303736e-12, 5.289962e-12, 5.236321e-12, 5.252083e-12, 5.205075e-12, 
    5.176813e-12, 5.158047e-12, 5.14473e-12, 5.146612e-12, 5.150201e-12, 
    5.168645e-12, 5.185988e-12, 5.199206e-12, 5.208048e-12, 5.216761e-12, 
    5.243132e-12, 5.257095e-12, 5.288359e-12, 5.282718e-12, 5.292276e-12, 
    5.301409e-12, 5.316742e-12, 5.314219e-12, 5.320974e-12, 5.292025e-12, 
    5.311264e-12, 5.279504e-12, 5.28819e-12, 5.219125e-12, 5.192826e-12, 
    5.181645e-12, 5.171862e-12, 5.14806e-12, 5.164496e-12, 5.158017e-12, 
    5.173433e-12, 5.18323e-12, 5.178385e-12, 5.20829e-12, 5.196663e-12, 
    5.257922e-12, 5.231534e-12, 5.300343e-12, 5.283876e-12, 5.304291e-12, 
    5.293874e-12, 5.311724e-12, 5.295659e-12, 5.323489e-12, 5.329549e-12, 
    5.325408e-12, 5.341318e-12, 5.294768e-12, 5.312643e-12, 5.178249e-12, 
    5.179039e-12, 5.18272e-12, 5.166537e-12, 5.165548e-12, 5.15072e-12, 
    5.163914e-12, 5.169532e-12, 5.183798e-12, 5.192235e-12, 5.200257e-12, 
    5.217895e-12, 5.237595e-12, 5.265146e-12, 5.284943e-12, 5.298214e-12, 
    5.290077e-12, 5.297261e-12, 5.28923e-12, 5.285466e-12, 5.327278e-12, 
    5.303799e-12, 5.339029e-12, 5.33708e-12, 5.321135e-12, 5.337299e-12, 
    5.179594e-12, 5.175047e-12, 5.159259e-12, 5.171614e-12, 5.149106e-12, 
    5.161704e-12, 5.168948e-12, 5.196905e-12, 5.203048e-12, 5.208744e-12, 
    5.219995e-12, 5.234435e-12, 5.259768e-12, 5.281813e-12, 5.30194e-12, 
    5.300466e-12, 5.300985e-12, 5.305481e-12, 5.294344e-12, 5.30731e-12, 
    5.309485e-12, 5.303796e-12, 5.336819e-12, 5.327384e-12, 5.337038e-12, 
    5.330895e-12, 5.176525e-12, 5.184176e-12, 5.180042e-12, 5.187816e-12, 
    5.182339e-12, 5.206695e-12, 5.213999e-12, 5.248177e-12, 5.234151e-12, 
    5.256476e-12, 5.236419e-12, 5.239972e-12, 5.257202e-12, 5.237503e-12, 
    5.280596e-12, 5.251378e-12, 5.305656e-12, 5.276472e-12, 5.307484e-12, 
    5.301854e-12, 5.311178e-12, 5.319528e-12, 5.330035e-12, 5.349422e-12, 
    5.344933e-12, 5.361148e-12, 5.195584e-12, 5.205508e-12, 5.204635e-12, 
    5.215022e-12, 5.222705e-12, 5.239358e-12, 5.266069e-12, 5.256024e-12, 
    5.274466e-12, 5.278169e-12, 5.250151e-12, 5.267352e-12, 5.212151e-12, 
    5.221068e-12, 5.21576e-12, 5.196366e-12, 5.258338e-12, 5.226531e-12, 
    5.28527e-12, 5.268036e-12, 5.318337e-12, 5.29332e-12, 5.342462e-12, 
    5.363471e-12, 5.383251e-12, 5.406363e-12, 5.210926e-12, 5.204182e-12, 
    5.216258e-12, 5.232966e-12, 5.248472e-12, 5.269087e-12, 5.271197e-12, 
    5.275059e-12, 5.285064e-12, 5.293477e-12, 5.276279e-12, 5.295585e-12, 
    5.223135e-12, 5.261099e-12, 5.201632e-12, 5.219536e-12, 5.231982e-12, 
    5.226523e-12, 5.254877e-12, 5.26156e-12, 5.28872e-12, 5.27468e-12, 
    5.358285e-12, 5.321291e-12, 5.423966e-12, 5.395267e-12, 5.201826e-12, 
    5.210903e-12, 5.242499e-12, 5.227465e-12, 5.270464e-12, 5.281049e-12, 
    5.289655e-12, 5.300656e-12, 5.301844e-12, 5.308362e-12, 5.297681e-12, 
    5.307941e-12, 5.269131e-12, 5.286473e-12, 5.238888e-12, 5.250468e-12, 
    5.245141e-12, 5.239297e-12, 5.257334e-12, 5.27655e-12, 5.276962e-12, 
    5.283124e-12, 5.300487e-12, 5.270639e-12, 5.363058e-12, 5.305975e-12, 
    5.220802e-12, 5.238287e-12, 5.240787e-12, 5.234013e-12, 5.279988e-12, 
    5.263328e-12, 5.308204e-12, 5.296075e-12, 5.315948e-12, 5.306072e-12, 
    5.304619e-12, 5.291936e-12, 5.28404e-12, 5.264092e-12, 5.247862e-12, 
    5.234996e-12, 5.237988e-12, 5.252122e-12, 5.277726e-12, 5.301951e-12, 
    5.296644e-12, 5.314438e-12, 5.267346e-12, 5.287091e-12, 5.279459e-12, 
    5.299359e-12, 5.255758e-12, 5.292882e-12, 5.246269e-12, 5.250355e-12, 
    5.262998e-12, 5.288429e-12, 5.294058e-12, 5.300066e-12, 5.296358e-12, 
    5.278376e-12, 5.275431e-12, 5.26269e-12, 5.259172e-12, 5.249466e-12, 
    5.241429e-12, 5.248771e-12, 5.256482e-12, 5.278384e-12, 5.298123e-12, 
    5.319647e-12, 5.324915e-12, 5.350064e-12, 5.32959e-12, 5.363376e-12, 
    5.334649e-12, 5.384381e-12, 5.295036e-12, 5.333806e-12, 5.263573e-12, 
    5.271139e-12, 5.284822e-12, 5.316211e-12, 5.299266e-12, 5.319084e-12, 
    5.275315e-12, 5.25261e-12, 5.246737e-12, 5.235778e-12, 5.246987e-12, 
    5.246075e-12, 5.256802e-12, 5.253355e-12, 5.279111e-12, 5.265276e-12, 
    5.304583e-12, 5.318928e-12, 5.359448e-12, 5.384292e-12, 5.409586e-12, 
    5.420754e-12, 5.424152e-12, 5.425574e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818189, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 
    1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818189, 1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818189, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.117302e-11, 3.131151e-11, 3.128459e-11, 3.13963e-11, 3.133433e-11, 
    3.140748e-11, 3.12011e-11, 3.1317e-11, 3.124302e-11, 3.118549e-11, 
    3.16131e-11, 3.140128e-11, 3.183321e-11, 3.169808e-11, 3.203757e-11, 
    3.181218e-11, 3.208303e-11, 3.203108e-11, 3.218746e-11, 3.214266e-11, 
    3.234269e-11, 3.220814e-11, 3.244641e-11, 3.231056e-11, 3.23318e-11, 
    3.22037e-11, 3.144391e-11, 3.158673e-11, 3.143545e-11, 3.145581e-11, 
    3.144668e-11, 3.133561e-11, 3.127964e-11, 3.116244e-11, 3.118372e-11, 
    3.12698e-11, 3.146497e-11, 3.139872e-11, 3.156572e-11, 3.156194e-11, 
    3.174788e-11, 3.166404e-11, 3.197661e-11, 3.188777e-11, 3.214453e-11, 
    3.207995e-11, 3.214149e-11, 3.212283e-11, 3.214173e-11, 3.204702e-11, 
    3.20876e-11, 3.200427e-11, 3.167974e-11, 3.17751e-11, 3.14907e-11, 
    3.131972e-11, 3.120618e-11, 3.112562e-11, 3.113701e-11, 3.115872e-11, 
    3.12703e-11, 3.137523e-11, 3.14552e-11, 3.150869e-11, 3.15614e-11, 
    3.172095e-11, 3.180542e-11, 3.199457e-11, 3.196044e-11, 3.201827e-11, 
    3.207352e-11, 3.216629e-11, 3.215102e-11, 3.219189e-11, 3.201675e-11, 
    3.213314e-11, 3.1941e-11, 3.199355e-11, 3.157571e-11, 3.14166e-11, 
    3.134895e-11, 3.128976e-11, 3.114576e-11, 3.12452e-11, 3.1206e-11, 
    3.129927e-11, 3.135854e-11, 3.132923e-11, 3.151015e-11, 3.143981e-11, 
    3.181043e-11, 3.165078e-11, 3.206708e-11, 3.196745e-11, 3.209096e-11, 
    3.202794e-11, 3.213593e-11, 3.203874e-11, 3.220711e-11, 3.224377e-11, 
    3.221871e-11, 3.231497e-11, 3.203335e-11, 3.214149e-11, 3.132841e-11, 
    3.133319e-11, 3.135546e-11, 3.125755e-11, 3.125156e-11, 3.116186e-11, 
    3.124168e-11, 3.127567e-11, 3.136198e-11, 3.141302e-11, 3.146156e-11, 
    3.156826e-11, 3.168745e-11, 3.185413e-11, 3.197391e-11, 3.20542e-11, 
    3.200496e-11, 3.204843e-11, 3.199984e-11, 3.197707e-11, 3.223003e-11, 
    3.208798e-11, 3.230113e-11, 3.228933e-11, 3.219287e-11, 3.229066e-11, 
    3.133654e-11, 3.130903e-11, 3.121352e-11, 3.128827e-11, 3.115209e-11, 
    3.122831e-11, 3.127214e-11, 3.144127e-11, 3.147844e-11, 3.15129e-11, 
    3.158097e-11, 3.166833e-11, 3.18216e-11, 3.195497e-11, 3.207674e-11, 
    3.206782e-11, 3.207096e-11, 3.209816e-11, 3.203078e-11, 3.210922e-11, 
    3.212239e-11, 3.208796e-11, 3.228775e-11, 3.223067e-11, 3.228908e-11, 
    3.225192e-11, 3.131798e-11, 3.136427e-11, 3.133925e-11, 3.138629e-11, 
    3.135315e-11, 3.150051e-11, 3.154469e-11, 3.175147e-11, 3.166661e-11, 
    3.180168e-11, 3.168033e-11, 3.170183e-11, 3.180608e-11, 3.168689e-11, 
    3.194761e-11, 3.177084e-11, 3.209922e-11, 3.192266e-11, 3.211028e-11, 
    3.207621e-11, 3.213262e-11, 3.218315e-11, 3.224671e-11, 3.2364e-11, 
    3.233685e-11, 3.243494e-11, 3.143328e-11, 3.149333e-11, 3.148804e-11, 
    3.155089e-11, 3.159736e-11, 3.169812e-11, 3.185972e-11, 3.179895e-11, 
    3.191052e-11, 3.193292e-11, 3.176341e-11, 3.186748e-11, 3.153352e-11, 
    3.158746e-11, 3.155535e-11, 3.143802e-11, 3.181294e-11, 3.162051e-11, 
    3.197588e-11, 3.187162e-11, 3.217594e-11, 3.202458e-11, 3.232189e-11, 
    3.2449e-11, 3.256867e-11, 3.27085e-11, 3.15261e-11, 3.14853e-11, 
    3.155836e-11, 3.165945e-11, 3.175326e-11, 3.187798e-11, 3.189074e-11, 
    3.191411e-11, 3.197464e-11, 3.202553e-11, 3.192149e-11, 3.203829e-11, 
    3.159997e-11, 3.182965e-11, 3.146987e-11, 3.157819e-11, 3.165349e-11, 
    3.162046e-11, 3.1792e-11, 3.183244e-11, 3.199675e-11, 3.191181e-11, 
    3.241762e-11, 3.219381e-11, 3.281499e-11, 3.264137e-11, 3.147104e-11, 
    3.152596e-11, 3.171712e-11, 3.162616e-11, 3.188631e-11, 3.195035e-11, 
    3.200241e-11, 3.206897e-11, 3.207616e-11, 3.211559e-11, 3.205097e-11, 
    3.211304e-11, 3.187824e-11, 3.198316e-11, 3.169527e-11, 3.176533e-11, 
    3.17331e-11, 3.169775e-11, 3.180687e-11, 3.192313e-11, 3.192562e-11, 
    3.19629e-11, 3.206794e-11, 3.188736e-11, 3.24465e-11, 3.210115e-11, 
    3.158586e-11, 3.169164e-11, 3.170676e-11, 3.166578e-11, 3.194393e-11, 
    3.184314e-11, 3.211463e-11, 3.204125e-11, 3.216149e-11, 3.210174e-11, 
    3.209295e-11, 3.201621e-11, 3.196844e-11, 3.184775e-11, 3.174957e-11, 
    3.167172e-11, 3.168982e-11, 3.177534e-11, 3.193024e-11, 3.20768e-11, 
    3.20447e-11, 3.215235e-11, 3.186744e-11, 3.19869e-11, 3.194072e-11, 
    3.206112e-11, 3.179733e-11, 3.202194e-11, 3.173992e-11, 3.176465e-11, 
    3.184113e-11, 3.199499e-11, 3.202905e-11, 3.20654e-11, 3.204297e-11, 
    3.193418e-11, 3.191635e-11, 3.183928e-11, 3.181799e-11, 3.175927e-11, 
    3.171065e-11, 3.175507e-11, 3.180172e-11, 3.193422e-11, 3.205365e-11, 
    3.218386e-11, 3.221574e-11, 3.236789e-11, 3.224402e-11, 3.244842e-11, 
    3.227463e-11, 3.25755e-11, 3.203497e-11, 3.226952e-11, 3.184462e-11, 
    3.189039e-11, 3.197317e-11, 3.216308e-11, 3.206056e-11, 3.218046e-11, 
    3.191566e-11, 3.177829e-11, 3.174275e-11, 3.167645e-11, 3.174427e-11, 
    3.173876e-11, 3.180365e-11, 3.17828e-11, 3.193862e-11, 3.185492e-11, 
    3.209272e-11, 3.217952e-11, 3.242466e-11, 3.257496e-11, 3.272799e-11, 
    3.279556e-11, 3.281612e-11, 3.282472e-11 ;

 SOILC =
  17.3448, 17.34479, 17.34479, 17.34478, 17.34479, 17.34478, 17.3448, 
    17.34479, 17.3448, 17.3448, 17.34476, 17.34478, 17.34474, 17.34475, 
    17.34472, 17.34474, 17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34468, 17.3447, 17.34469, 17.34471, 17.34478, 17.34476, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.34479, 17.3448, 17.3448, 
    17.3448, 17.34478, 17.34478, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34471, 17.34472, 17.34471, 17.34471, 17.34471, 
    17.34472, 17.34472, 17.34472, 17.34476, 17.34475, 17.34477, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 
    17.34477, 17.34477, 17.34475, 17.34474, 17.34472, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.34471, 17.34472, 17.34471, 17.34473, 
    17.34472, 17.34476, 17.34478, 17.34479, 17.34479, 17.34481, 17.3448, 
    17.3448, 17.34479, 17.34479, 17.34479, 17.34477, 17.34478, 17.34474, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34472, 17.34471, 17.34472, 
    17.34471, 17.3447, 17.3447, 17.34469, 17.34472, 17.34471, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.3448, 17.3448, 17.34479, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34472, 17.34473, 17.3447, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.3448, 17.34479, 17.34478, 17.34477, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34472, 17.3447, 17.3447, 
    17.3447, 17.3447, 17.34479, 17.34479, 17.34479, 17.34478, 17.34479, 
    17.34477, 17.34477, 17.34475, 17.34476, 17.34474, 17.34476, 17.34475, 
    17.34474, 17.34476, 17.34473, 17.34475, 17.34472, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.34469, 17.34469, 17.34468, 
    17.34478, 17.34477, 17.34477, 17.34477, 17.34476, 17.34475, 17.34474, 
    17.34474, 17.34473, 17.34473, 17.34475, 17.34474, 17.34477, 17.34476, 
    17.34477, 17.34478, 17.34474, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34472, 17.34469, 17.34468, 17.34467, 17.34466, 17.34477, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34476, 17.34474, 17.34478, 17.34476, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34472, 17.34473, 17.34468, 
    17.34471, 17.34465, 17.34466, 17.34478, 17.34477, 17.34475, 17.34476, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34471, 17.34472, 
    17.34471, 17.34474, 17.34473, 17.34475, 17.34475, 17.34475, 17.34475, 
    17.34474, 17.34473, 17.34473, 17.34473, 17.34472, 17.34474, 17.34468, 
    17.34472, 17.34476, 17.34476, 17.34475, 17.34476, 17.34473, 17.34474, 
    17.34471, 17.34472, 17.34471, 17.34472, 17.34472, 17.34472, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34474, 17.34473, 17.34473, 17.34472, 17.34474, 
    17.34472, 17.34475, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 
    17.34475, 17.34474, 17.34473, 17.34472, 17.34471, 17.3447, 17.34469, 
    17.3447, 17.34468, 17.3447, 17.34467, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34473, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34468, 17.34467, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 SOILC_HR =
  6.194319e-08, 6.221824e-08, 6.216477e-08, 6.238663e-08, 6.226357e-08, 
    6.240884e-08, 6.199895e-08, 6.222916e-08, 6.20822e-08, 6.196796e-08, 
    6.281724e-08, 6.239654e-08, 6.325438e-08, 6.2986e-08, 6.366027e-08, 
    6.321261e-08, 6.375054e-08, 6.364737e-08, 6.395796e-08, 6.386897e-08, 
    6.426626e-08, 6.399903e-08, 6.447225e-08, 6.420245e-08, 6.424465e-08, 
    6.399021e-08, 6.248121e-08, 6.276485e-08, 6.24644e-08, 6.250485e-08, 
    6.24867e-08, 6.22661e-08, 6.215493e-08, 6.192218e-08, 6.196444e-08, 
    6.213539e-08, 6.252303e-08, 6.239145e-08, 6.272312e-08, 6.271563e-08, 
    6.308491e-08, 6.29184e-08, 6.35392e-08, 6.336274e-08, 6.387269e-08, 
    6.374443e-08, 6.386666e-08, 6.38296e-08, 6.386715e-08, 6.367905e-08, 
    6.375964e-08, 6.359412e-08, 6.294958e-08, 6.313898e-08, 6.257413e-08, 
    6.223455e-08, 6.200905e-08, 6.184904e-08, 6.187166e-08, 6.191478e-08, 
    6.213639e-08, 6.234479e-08, 6.250362e-08, 6.260986e-08, 6.271455e-08, 
    6.303143e-08, 6.31992e-08, 6.357487e-08, 6.350708e-08, 6.362193e-08, 
    6.373168e-08, 6.391591e-08, 6.388559e-08, 6.396677e-08, 6.361891e-08, 
    6.385008e-08, 6.346847e-08, 6.357283e-08, 6.274296e-08, 6.242695e-08, 
    6.22926e-08, 6.217505e-08, 6.188905e-08, 6.208655e-08, 6.200869e-08, 
    6.219393e-08, 6.231164e-08, 6.225343e-08, 6.261276e-08, 6.247306e-08, 
    6.320914e-08, 6.289206e-08, 6.371887e-08, 6.352099e-08, 6.37663e-08, 
    6.364113e-08, 6.385561e-08, 6.366258e-08, 6.399698e-08, 6.406979e-08, 
    6.402004e-08, 6.421121e-08, 6.365187e-08, 6.386666e-08, 6.225179e-08, 
    6.226129e-08, 6.230552e-08, 6.211108e-08, 6.209918e-08, 6.192101e-08, 
    6.207955e-08, 6.214706e-08, 6.231847e-08, 6.241986e-08, 6.251624e-08, 
    6.272818e-08, 6.296489e-08, 6.329594e-08, 6.353382e-08, 6.369329e-08, 
    6.359551e-08, 6.368183e-08, 6.358533e-08, 6.35401e-08, 6.404251e-08, 
    6.376038e-08, 6.418371e-08, 6.416029e-08, 6.39687e-08, 6.416293e-08, 
    6.226796e-08, 6.221332e-08, 6.202362e-08, 6.217208e-08, 6.190162e-08, 
    6.2053e-08, 6.214005e-08, 6.247596e-08, 6.254979e-08, 6.261823e-08, 
    6.275342e-08, 6.292692e-08, 6.323132e-08, 6.349621e-08, 6.373806e-08, 
    6.372034e-08, 6.372658e-08, 6.37806e-08, 6.364677e-08, 6.380257e-08, 
    6.382872e-08, 6.376035e-08, 6.415715e-08, 6.404378e-08, 6.415979e-08, 
    6.408597e-08, 6.223108e-08, 6.232302e-08, 6.227334e-08, 6.236676e-08, 
    6.230094e-08, 6.259361e-08, 6.268137e-08, 6.309205e-08, 6.29235e-08, 
    6.319176e-08, 6.295076e-08, 6.299346e-08, 6.32005e-08, 6.296379e-08, 
    6.348159e-08, 6.313051e-08, 6.37827e-08, 6.343204e-08, 6.380468e-08, 
    6.373701e-08, 6.384905e-08, 6.394939e-08, 6.407564e-08, 6.430859e-08, 
    6.425465e-08, 6.444949e-08, 6.246009e-08, 6.257934e-08, 6.256885e-08, 
    6.269367e-08, 6.278598e-08, 6.298608e-08, 6.330703e-08, 6.318634e-08, 
    6.340794e-08, 6.345242e-08, 6.311577e-08, 6.332245e-08, 6.265917e-08, 
    6.276631e-08, 6.270252e-08, 6.24695e-08, 6.321414e-08, 6.283195e-08, 
    6.353775e-08, 6.333067e-08, 6.393508e-08, 6.363447e-08, 6.422496e-08, 
    6.44774e-08, 6.471507e-08, 6.499279e-08, 6.264444e-08, 6.256341e-08, 
    6.270852e-08, 6.290927e-08, 6.309559e-08, 6.334329e-08, 6.336865e-08, 
    6.341506e-08, 6.353527e-08, 6.363636e-08, 6.342972e-08, 6.366169e-08, 
    6.279114e-08, 6.324732e-08, 6.253276e-08, 6.274789e-08, 6.289744e-08, 
    6.283185e-08, 6.317255e-08, 6.325285e-08, 6.35792e-08, 6.34105e-08, 
    6.441508e-08, 6.397057e-08, 6.52043e-08, 6.485946e-08, 6.253509e-08, 
    6.264417e-08, 6.302381e-08, 6.284317e-08, 6.335984e-08, 6.348703e-08, 
    6.359044e-08, 6.372262e-08, 6.37369e-08, 6.381522e-08, 6.368688e-08, 
    6.381016e-08, 6.334383e-08, 6.355221e-08, 6.298043e-08, 6.311958e-08, 
    6.305557e-08, 6.298534e-08, 6.320207e-08, 6.343297e-08, 6.343792e-08, 
    6.351196e-08, 6.372059e-08, 6.336194e-08, 6.447243e-08, 6.378654e-08, 
    6.276311e-08, 6.297321e-08, 6.300324e-08, 6.292185e-08, 6.347427e-08, 
    6.32741e-08, 6.381332e-08, 6.366758e-08, 6.390638e-08, 6.378771e-08, 
    6.377025e-08, 6.361785e-08, 6.352296e-08, 6.328327e-08, 6.308827e-08, 
    6.293366e-08, 6.296961e-08, 6.313945e-08, 6.34471e-08, 6.373818e-08, 
    6.367442e-08, 6.388823e-08, 6.332237e-08, 6.355963e-08, 6.346792e-08, 
    6.370704e-08, 6.318313e-08, 6.362922e-08, 6.306912e-08, 6.311822e-08, 
    6.327013e-08, 6.35757e-08, 6.364334e-08, 6.371553e-08, 6.367099e-08, 
    6.345491e-08, 6.341952e-08, 6.326643e-08, 6.322416e-08, 6.310753e-08, 
    6.301097e-08, 6.309919e-08, 6.319184e-08, 6.3455e-08, 6.369219e-08, 
    6.395081e-08, 6.401412e-08, 6.43163e-08, 6.407029e-08, 6.447625e-08, 
    6.413108e-08, 6.472865e-08, 6.36551e-08, 6.412095e-08, 6.327704e-08, 
    6.336795e-08, 6.353237e-08, 6.390953e-08, 6.370593e-08, 6.394406e-08, 
    6.341813e-08, 6.314531e-08, 6.307474e-08, 6.294306e-08, 6.307775e-08, 
    6.306679e-08, 6.319569e-08, 6.315427e-08, 6.346375e-08, 6.329751e-08, 
    6.376981e-08, 6.394218e-08, 6.442907e-08, 6.472758e-08, 6.503151e-08, 
    6.51657e-08, 6.520654e-08, 6.522362e-08 ;

 SOILC_LOSS =
  6.194319e-08, 6.221824e-08, 6.216477e-08, 6.238663e-08, 6.226357e-08, 
    6.240884e-08, 6.199895e-08, 6.222916e-08, 6.20822e-08, 6.196796e-08, 
    6.281724e-08, 6.239654e-08, 6.325438e-08, 6.2986e-08, 6.366027e-08, 
    6.321261e-08, 6.375054e-08, 6.364737e-08, 6.395796e-08, 6.386897e-08, 
    6.426626e-08, 6.399903e-08, 6.447225e-08, 6.420245e-08, 6.424465e-08, 
    6.399021e-08, 6.248121e-08, 6.276485e-08, 6.24644e-08, 6.250485e-08, 
    6.24867e-08, 6.22661e-08, 6.215493e-08, 6.192218e-08, 6.196444e-08, 
    6.213539e-08, 6.252303e-08, 6.239145e-08, 6.272312e-08, 6.271563e-08, 
    6.308491e-08, 6.29184e-08, 6.35392e-08, 6.336274e-08, 6.387269e-08, 
    6.374443e-08, 6.386666e-08, 6.38296e-08, 6.386715e-08, 6.367905e-08, 
    6.375964e-08, 6.359412e-08, 6.294958e-08, 6.313898e-08, 6.257413e-08, 
    6.223455e-08, 6.200905e-08, 6.184904e-08, 6.187166e-08, 6.191478e-08, 
    6.213639e-08, 6.234479e-08, 6.250362e-08, 6.260986e-08, 6.271455e-08, 
    6.303143e-08, 6.31992e-08, 6.357487e-08, 6.350708e-08, 6.362193e-08, 
    6.373168e-08, 6.391591e-08, 6.388559e-08, 6.396677e-08, 6.361891e-08, 
    6.385008e-08, 6.346847e-08, 6.357283e-08, 6.274296e-08, 6.242695e-08, 
    6.22926e-08, 6.217505e-08, 6.188905e-08, 6.208655e-08, 6.200869e-08, 
    6.219393e-08, 6.231164e-08, 6.225343e-08, 6.261276e-08, 6.247306e-08, 
    6.320914e-08, 6.289206e-08, 6.371887e-08, 6.352099e-08, 6.37663e-08, 
    6.364113e-08, 6.385561e-08, 6.366258e-08, 6.399698e-08, 6.406979e-08, 
    6.402004e-08, 6.421121e-08, 6.365187e-08, 6.386666e-08, 6.225179e-08, 
    6.226129e-08, 6.230552e-08, 6.211108e-08, 6.209918e-08, 6.192101e-08, 
    6.207955e-08, 6.214706e-08, 6.231847e-08, 6.241986e-08, 6.251624e-08, 
    6.272818e-08, 6.296489e-08, 6.329594e-08, 6.353382e-08, 6.369329e-08, 
    6.359551e-08, 6.368183e-08, 6.358533e-08, 6.35401e-08, 6.404251e-08, 
    6.376038e-08, 6.418371e-08, 6.416029e-08, 6.39687e-08, 6.416293e-08, 
    6.226796e-08, 6.221332e-08, 6.202362e-08, 6.217208e-08, 6.190162e-08, 
    6.2053e-08, 6.214005e-08, 6.247596e-08, 6.254979e-08, 6.261823e-08, 
    6.275342e-08, 6.292692e-08, 6.323132e-08, 6.349621e-08, 6.373806e-08, 
    6.372034e-08, 6.372658e-08, 6.37806e-08, 6.364677e-08, 6.380257e-08, 
    6.382872e-08, 6.376035e-08, 6.415715e-08, 6.404378e-08, 6.415979e-08, 
    6.408597e-08, 6.223108e-08, 6.232302e-08, 6.227334e-08, 6.236676e-08, 
    6.230094e-08, 6.259361e-08, 6.268137e-08, 6.309205e-08, 6.29235e-08, 
    6.319176e-08, 6.295076e-08, 6.299346e-08, 6.32005e-08, 6.296379e-08, 
    6.348159e-08, 6.313051e-08, 6.37827e-08, 6.343204e-08, 6.380468e-08, 
    6.373701e-08, 6.384905e-08, 6.394939e-08, 6.407564e-08, 6.430859e-08, 
    6.425465e-08, 6.444949e-08, 6.246009e-08, 6.257934e-08, 6.256885e-08, 
    6.269367e-08, 6.278598e-08, 6.298608e-08, 6.330703e-08, 6.318634e-08, 
    6.340794e-08, 6.345242e-08, 6.311577e-08, 6.332245e-08, 6.265917e-08, 
    6.276631e-08, 6.270252e-08, 6.24695e-08, 6.321414e-08, 6.283195e-08, 
    6.353775e-08, 6.333067e-08, 6.393508e-08, 6.363447e-08, 6.422496e-08, 
    6.44774e-08, 6.471507e-08, 6.499279e-08, 6.264444e-08, 6.256341e-08, 
    6.270852e-08, 6.290927e-08, 6.309559e-08, 6.334329e-08, 6.336865e-08, 
    6.341506e-08, 6.353527e-08, 6.363636e-08, 6.342972e-08, 6.366169e-08, 
    6.279114e-08, 6.324732e-08, 6.253276e-08, 6.274789e-08, 6.289744e-08, 
    6.283185e-08, 6.317255e-08, 6.325285e-08, 6.35792e-08, 6.34105e-08, 
    6.441508e-08, 6.397057e-08, 6.52043e-08, 6.485946e-08, 6.253509e-08, 
    6.264417e-08, 6.302381e-08, 6.284317e-08, 6.335984e-08, 6.348703e-08, 
    6.359044e-08, 6.372262e-08, 6.37369e-08, 6.381522e-08, 6.368688e-08, 
    6.381016e-08, 6.334383e-08, 6.355221e-08, 6.298043e-08, 6.311958e-08, 
    6.305557e-08, 6.298534e-08, 6.320207e-08, 6.343297e-08, 6.343792e-08, 
    6.351196e-08, 6.372059e-08, 6.336194e-08, 6.447243e-08, 6.378654e-08, 
    6.276311e-08, 6.297321e-08, 6.300324e-08, 6.292185e-08, 6.347427e-08, 
    6.32741e-08, 6.381332e-08, 6.366758e-08, 6.390638e-08, 6.378771e-08, 
    6.377025e-08, 6.361785e-08, 6.352296e-08, 6.328327e-08, 6.308827e-08, 
    6.293366e-08, 6.296961e-08, 6.313945e-08, 6.34471e-08, 6.373818e-08, 
    6.367442e-08, 6.388823e-08, 6.332237e-08, 6.355963e-08, 6.346792e-08, 
    6.370704e-08, 6.318313e-08, 6.362922e-08, 6.306912e-08, 6.311822e-08, 
    6.327013e-08, 6.35757e-08, 6.364334e-08, 6.371553e-08, 6.367099e-08, 
    6.345491e-08, 6.341952e-08, 6.326643e-08, 6.322416e-08, 6.310753e-08, 
    6.301097e-08, 6.309919e-08, 6.319184e-08, 6.3455e-08, 6.369219e-08, 
    6.395081e-08, 6.401412e-08, 6.43163e-08, 6.407029e-08, 6.447625e-08, 
    6.413108e-08, 6.472865e-08, 6.36551e-08, 6.412095e-08, 6.327704e-08, 
    6.336795e-08, 6.353237e-08, 6.390953e-08, 6.370593e-08, 6.394406e-08, 
    6.341813e-08, 6.314531e-08, 6.307474e-08, 6.294306e-08, 6.307775e-08, 
    6.306679e-08, 6.319569e-08, 6.315427e-08, 6.346375e-08, 6.329751e-08, 
    6.376981e-08, 6.394218e-08, 6.442907e-08, 6.472758e-08, 6.503151e-08, 
    6.51657e-08, 6.520654e-08, 6.522362e-08 ;

 SOILICE =
  95.12831, 95.56489, 95.47991, 95.83276, 95.63691, 95.86811, 95.21671, 
    95.58227, 95.34879, 95.16753, 96.51984, 95.84852, 97.21997, 96.78965, 
    97.87275, 97.15296, 98.01825, 97.85188, 98.353, 98.20927, 98.852, 
    98.41936, 99.18605, 98.74854, 98.81693, 98.40512, 95.98334, 96.43613, 
    95.95657, 96.02104, 95.9921, 95.64097, 95.46436, 95.09496, 95.16195, 
    95.43327, 96.05004, 95.84037, 96.36922, 96.35725, 96.94808, 96.68143, 
    97.67769, 97.3939, 98.21527, 98.00833, 98.20555, 98.14572, 98.20634, 
    97.90293, 98.03286, 97.76611, 96.73134, 97.03478, 96.1315, 95.5909, 
    95.23273, 94.9791, 95.01493, 95.08327, 95.43486, 95.76611, 96.01903, 
    96.18844, 96.35554, 96.86253, 97.13141, 97.73516, 97.62599, 97.81094, 
    97.98775, 98.2851, 98.23611, 98.36726, 97.80602, 98.17883, 97.56385, 
    97.73183, 96.40117, 95.8969, 95.6832, 95.49625, 95.04249, 95.35571, 
    95.23217, 95.52621, 95.71337, 95.62077, 96.19308, 95.97034, 97.14736, 
    96.63931, 97.96712, 97.64839, 98.0436, 97.8418, 98.18774, 97.87637, 
    98.41608, 98.53384, 98.45336, 98.76269, 97.85913, 98.20557, 95.61819, 
    95.63329, 95.70363, 95.39465, 95.37576, 95.09313, 95.34458, 95.45179, 
    95.72421, 95.8856, 96.03917, 96.37733, 96.75587, 97.28666, 97.66904, 
    97.92586, 97.76832, 97.90739, 97.75194, 97.67912, 98.48972, 98.03408, 
    98.71816, 98.68023, 98.37038, 98.6845, 95.64389, 95.55701, 95.25584, 
    95.49149, 95.06239, 95.30245, 95.44067, 95.97503, 96.09264, 96.20182, 
    96.41764, 96.69506, 97.18291, 97.60854, 97.99804, 97.96947, 97.97952, 
    98.06667, 97.85091, 98.10212, 98.14433, 98.034, 98.67516, 98.49173, 
    98.67943, 98.55997, 95.58524, 95.73146, 95.65244, 95.80108, 95.69636, 
    96.1626, 96.30265, 96.95959, 96.68961, 97.11945, 96.7332, 96.80158, 
    97.13356, 96.75404, 97.58508, 97.02126, 98.07006, 97.50543, 98.10551, 
    97.99635, 98.1771, 98.33917, 98.54326, 98.92053, 98.83308, 99.14906, 
    95.94968, 96.13981, 96.12303, 96.3222, 96.46967, 96.78973, 97.30444, 
    97.11069, 97.46653, 97.53807, 96.99751, 97.32922, 96.26716, 96.43831, 
    96.33636, 95.96469, 97.15536, 96.54321, 97.67537, 97.34239, 98.31606, 
    97.83115, 98.78497, 99.19449, 99.58063, 100.0332, 96.24364, 96.11434, 
    96.3459, 96.66689, 96.96519, 97.36269, 97.40339, 97.478, 97.67136, 
    97.83412, 97.50163, 97.87495, 96.4781, 97.20859, 96.06551, 96.40891, 
    96.64793, 96.543, 97.08855, 97.21741, 97.74212, 97.47064, 99.09335, 
    98.37347, 100.3784, 99.8158, 96.0692, 96.24318, 96.85022, 96.5611, 
    97.38924, 97.59375, 97.76016, 97.97319, 97.99618, 98.12254, 97.91553, 
    98.11434, 97.36353, 97.69862, 96.78068, 97.00364, 96.90102, 96.78855, 
    97.13592, 97.50687, 97.51474, 97.63388, 97.97018, 97.3926, 99.1866, 
    98.07648, 96.43311, 96.76923, 96.81724, 96.68692, 97.57323, 97.25154, 
    98.11945, 97.88442, 98.26967, 98.07812, 98.04996, 97.80431, 97.65157, 
    97.26629, 96.95347, 96.70581, 96.76336, 97.03552, 97.52957, 97.99828, 
    97.89551, 98.24036, 97.32905, 97.71059, 97.56304, 97.94805, 97.10555, 
    97.82288, 96.92273, 97.00143, 97.24516, 97.73654, 97.84538, 97.96175, 
    97.88992, 97.54212, 97.48518, 97.23922, 97.1714, 96.98429, 96.82957, 
    96.97094, 97.11954, 97.54224, 97.92413, 98.34149, 98.44376, 98.93317, 
    98.53474, 99.19281, 98.63329, 99.60297, 97.86446, 98.61674, 97.25624, 
    97.40225, 97.66676, 98.27488, 97.94624, 98.33062, 97.48295, 97.04494, 
    96.93174, 96.72086, 96.93657, 96.91901, 97.12566, 97.05923, 97.5563, 
    97.2891, 98.04927, 98.32757, 99.11593, 99.60108, 100.0962, 100.3153, 
    100.3821, 100.41,
  94.75558, 95.22529, 95.13383, 95.51356, 95.30276, 95.55161, 94.85065, 
    95.244, 94.99275, 94.79774, 96.25324, 95.53051, 96.99527, 96.54363, 
    97.67678, 96.92535, 97.82872, 97.65495, 98.17826, 98.02816, 98.69962, 
    98.24759, 99.04862, 98.5915, 98.66296, 98.23272, 95.67559, 96.16311, 
    95.64678, 95.71619, 95.68502, 95.30715, 95.11714, 94.71967, 94.79173, 
    95.08367, 95.74741, 95.52171, 96.09095, 96.07806, 96.71143, 96.42709, 
    97.47306, 97.17677, 98.03442, 97.81831, 98.02428, 97.96178, 98.02509, 
    97.70825, 97.84393, 97.56538, 96.48084, 96.80194, 95.83508, 95.25333, 
    94.8679, 94.59504, 94.63359, 94.70712, 95.08538, 95.4418, 95.71399, 
    95.89635, 96.07622, 96.62218, 96.90282, 97.5331, 97.41908, 97.61221, 
    97.79682, 98.10736, 98.05619, 98.19318, 97.60705, 97.99638, 97.35419, 
    97.52959, 96.12549, 95.58256, 95.35264, 95.15142, 94.66324, 95.00022, 
    94.8673, 95.18365, 95.38505, 95.28539, 95.90134, 95.6616, 96.91947, 
    96.38177, 97.77528, 97.44247, 97.85514, 97.64441, 98.00568, 97.6805, 
    98.24416, 98.3672, 98.28312, 98.60624, 97.6625, 98.02431, 95.28262, 
    95.29887, 95.37456, 95.04212, 95.02179, 94.71771, 94.98822, 95.10358, 
    95.39671, 95.5704, 95.73569, 96.09969, 96.50728, 97.06485, 97.46402, 
    97.73218, 97.56767, 97.7129, 97.55057, 97.47453, 98.32111, 97.84522, 
    98.55972, 98.5201, 98.19645, 98.52456, 95.31027, 95.21678, 94.89275, 
    95.14628, 94.68462, 94.94291, 95.09164, 95.66667, 95.79322, 95.91076, 
    96.14307, 96.44177, 96.95654, 97.40088, 97.80755, 97.77771, 97.78822, 
    97.87923, 97.65392, 97.91625, 97.96036, 97.84512, 98.51479, 98.32318, 
    98.51925, 98.39445, 95.24716, 95.40451, 95.31947, 95.47945, 95.36675, 
    95.86857, 96.01934, 96.72348, 96.43591, 96.89031, 96.48284, 96.55648, 
    96.90512, 96.50526, 97.37642, 96.78787, 97.88277, 97.2933, 97.91979, 
    97.80579, 97.99455, 98.16385, 98.37701, 98.77119, 98.6798, 99.00994, 
    95.63936, 95.84402, 95.82594, 96.04034, 96.19911, 96.5437, 97.0834, 
    96.88113, 97.25259, 97.32729, 96.76299, 97.10928, 95.98111, 96.16538, 
    96.0556, 95.65553, 96.92781, 96.27832, 97.47064, 97.123, 98.13971, 
    97.63333, 98.62954, 99.05749, 99.46096, 99.9341, 95.95577, 95.81658, 
    96.06584, 96.41147, 96.72929, 97.1442, 97.18668, 97.26456, 97.46643, 
    97.63639, 97.28927, 97.67902, 96.20827, 96.98336, 95.76405, 96.13374, 
    96.39104, 96.27805, 96.85801, 96.99252, 97.54035, 97.25688, 98.95183, 
    98.19972, 100.295, 99.70683, 95.768, 95.95526, 96.60886, 96.29753, 
    97.1719, 97.38542, 97.55915, 97.78162, 97.80561, 97.93759, 97.72139, 
    97.92902, 97.14508, 97.49491, 96.53394, 96.76941, 96.66228, 96.54243, 
    96.90746, 97.29475, 97.30293, 97.42734, 97.77866, 97.17541, 99.04936, 
    97.88965, 96.15973, 96.52168, 96.57333, 96.433, 97.36401, 97.02817, 
    97.93436, 97.6889, 98.09124, 97.8912, 97.86179, 97.60526, 97.44578, 
    97.04357, 96.71705, 96.45333, 96.5153, 96.8027, 97.31844, 97.80784, 
    97.70052, 98.06062, 97.10907, 97.50743, 97.35338, 97.75536, 96.87579, 
    97.62482, 96.68494, 96.7671, 97.02151, 97.53457, 97.64813, 97.76969, 
    97.69465, 97.33154, 97.27208, 97.01529, 96.94452, 96.7492, 96.5866, 
    96.73528, 96.8904, 97.33164, 97.73041, 98.16628, 98.27308, 98.78448, 
    98.36821, 99.05587, 98.47128, 99.48445, 97.66817, 98.45389, 97.03306, 
    97.18549, 97.46169, 98.09676, 97.75346, 98.15496, 97.26974, 96.81256, 
    96.69435, 96.46955, 96.69939, 96.68106, 96.89676, 96.82741, 97.34631, 
    97.06736, 97.86108, 98.15176, 98.97535, 99.48239, 99.99995, 100.229, 
    100.2988, 100.328,
  128.9624, 129.6492, 129.5154, 130.0708, 129.7625, 130.1264, 129.1014, 
    129.6765, 129.3091, 129.0241, 131.153, 130.0956, 132.2566, 131.5781, 
    133.2867, 132.151, 133.5165, 133.2538, 134.0452, 133.8181, 134.8339, 
    134.15, 135.3622, 134.6703, 134.7784, 134.1275, 130.3078, 131.0211, 
    130.2656, 130.3672, 130.3216, 129.7689, 129.491, 128.9099, 129.0153, 
    129.4421, 130.4128, 130.0827, 130.9155, 130.8967, 131.8278, 131.4075, 
    132.9788, 132.5309, 133.8276, 133.5008, 133.8122, 133.7177, 133.8135, 
    133.3344, 133.5395, 133.1183, 131.4861, 131.9646, 130.5411, 129.6902, 
    129.1266, 128.7278, 128.7841, 128.8916, 129.4446, 129.9658, 130.364, 
    130.6308, 130.8939, 131.6931, 132.117, 133.0695, 132.8972, 133.1891, 
    133.4683, 133.9379, 133.8605, 134.0677, 133.1813, 133.7701, 132.7991, 
    133.0642, 130.966, 130.1717, 129.8354, 129.5412, 128.8274, 129.3201, 
    129.1257, 129.5883, 129.8828, 129.7371, 130.638, 130.2873, 132.1421, 
    131.3411, 133.4357, 132.9325, 133.5565, 133.2378, 133.7841, 133.2924, 
    134.1448, 134.3309, 134.2038, 134.6926, 133.2652, 133.8123, 129.733, 
    129.7568, 129.8675, 129.3813, 129.3516, 128.9071, 129.3025, 129.4712, 
    129.8999, 130.1539, 130.3957, 130.9283, 131.5248, 132.3618, 132.9651, 
    133.3705, 133.1218, 133.3414, 133.096, 132.981, 134.2612, 133.5414, 
    134.6222, 134.5623, 134.0726, 134.569, 129.7735, 129.6367, 129.1629, 
    129.5336, 128.8587, 129.2363, 129.4537, 130.2947, 130.4799, 130.6518, 
    130.9918, 131.429, 132.1981, 132.8697, 133.4845, 133.4394, 133.4553, 
    133.5929, 133.2522, 133.6489, 133.7156, 133.5413, 134.5542, 134.2644, 
    134.561, 134.3722, 129.6812, 129.9113, 129.7869, 130.0209, 129.856, 
    130.5901, 130.8107, 131.846, 131.4204, 132.0981, 131.4891, 131.5969, 
    132.1204, 131.5219, 132.8327, 131.9433, 133.5982, 132.707, 133.6542, 
    133.4818, 133.7673, 134.0233, 134.3458, 134.9422, 134.8039, 135.3036, 
    130.2548, 130.5542, 130.5277, 130.8414, 131.0738, 131.5782, 132.3898, 
    132.0842, 132.6455, 132.7584, 131.9057, 132.4289, 130.7548, 131.0244, 
    130.8638, 130.2784, 132.1547, 131.1897, 132.9751, 132.4497, 133.9868, 
    133.2211, 134.7279, 135.3755, 135.9865, 136.7031, 130.7177, 130.5141, 
    130.8788, 131.3846, 131.8548, 132.4817, 132.5459, 132.6636, 132.9688, 
    133.2257, 132.701, 133.2901, 131.0872, 132.2387, 130.4372, 130.9781, 
    131.3547, 131.1893, 132.0493, 132.2525, 133.0805, 132.652, 135.2156, 
    134.0776, 137.25, 136.3588, 130.443, 130.717, 131.6736, 131.2178, 
    132.5236, 132.8463, 133.1089, 133.4453, 133.4816, 133.6811, 133.3542, 
    133.6682, 132.483, 133.0118, 131.5639, 131.9154, 131.7536, 131.5763, 
    132.124, 132.7092, 132.7216, 132.9097, 133.4407, 132.5289, 135.3632, 
    133.6086, 131.0162, 131.5459, 131.6215, 131.4161, 132.8139, 132.3064, 
    133.6762, 133.3051, 133.9135, 133.611, 133.5665, 133.1786, 132.9375, 
    132.3297, 131.8363, 131.4459, 131.5366, 131.9657, 132.745, 133.4849, 
    133.3226, 133.8672, 132.4286, 133.0307, 132.7979, 133.4056, 132.0761, 
    133.2081, 131.7878, 131.9119, 132.2963, 133.0717, 133.2435, 133.4272, 
    133.3138, 132.7648, 132.675, 132.2869, 132.18, 131.8849, 131.641, 
    131.8639, 132.0982, 132.765, 133.3678, 134.027, 134.1886, 134.9623, 
    134.3324, 135.373, 134.4883, 136.022, 133.2737, 134.4621, 132.3138, 
    132.5441, 132.9616, 133.9218, 133.4027, 134.0099, 132.6714, 131.9806, 
    131.802, 131.4696, 131.8096, 131.782, 132.1078, 132.0031, 132.7872, 
    132.3656, 133.5654, 134.005, 135.2512, 136.0189, 136.8029, 137.15, 
    137.2557, 137.3,
  194.2189, 195.2933, 195.0842, 195.9527, 195.4705, 196.0398, 194.437, 
    195.3361, 194.7617, 194.3161, 197.6465, 195.9915, 199.3758, 198.3124, 
    200.9915, 199.2102, 201.3521, 200.9398, 202.1822, 201.8257, 203.4213, 
    202.3469, 204.2518, 203.1642, 203.3342, 202.3115, 196.3236, 197.44, 
    196.2576, 196.4165, 196.3452, 195.4806, 195.046, 194.134, 194.3024, 
    194.9695, 196.4879, 195.9714, 197.2748, 197.2453, 198.7038, 198.0452, 
    200.5084, 199.806, 201.8405, 201.3275, 201.8164, 201.6681, 201.8184, 
    201.0663, 201.3883, 200.7273, 198.1684, 198.918, 196.6887, 195.3574, 
    194.4764, 193.8394, 193.9305, 194.1043, 194.9734, 195.7886, 196.4115, 
    196.829, 197.241, 198.4925, 199.1569, 200.6507, 200.3804, 200.8384, 
    201.2765, 202.0137, 201.8922, 202.2176, 200.8262, 201.7502, 200.2265, 
    200.6424, 197.3537, 196.1106, 195.5845, 195.1244, 194.0006, 194.7788, 
    194.475, 195.1982, 195.6587, 195.4308, 196.8405, 196.2915, 199.1963, 
    197.9413, 201.2253, 200.4358, 201.4149, 200.9148, 201.7723, 201.0004, 
    202.3387, 202.6311, 202.4313, 203.1993, 200.9577, 201.8165, 195.4245, 
    195.4616, 195.6348, 194.8746, 194.8281, 194.1294, 194.7514, 195.0151, 
    195.6854, 196.0828, 196.4612, 197.2948, 198.229, 199.5407, 200.4869, 
    201.1231, 200.7328, 201.0773, 200.6922, 200.5119, 202.5215, 201.3913, 
    203.0887, 202.9945, 202.2253, 203.0051, 195.4877, 195.2739, 194.5332, 
    195.1127, 194.0512, 194.6478, 194.9877, 196.3031, 196.5929, 196.862, 
    197.3942, 198.0789, 199.2842, 200.3372, 201.3019, 201.2311, 201.2561, 
    201.4721, 200.9374, 201.56, 201.6646, 201.3911, 202.9819, 202.5265, 
    202.9925, 202.6959, 195.3434, 195.7033, 195.5088, 195.8747, 195.6169, 
    196.7654, 197.1107, 198.7322, 198.0654, 199.1273, 198.173, 198.3419, 
    199.1622, 198.2245, 200.2791, 198.8846, 201.4805, 200.082, 201.5684, 
    201.2978, 201.7459, 202.1479, 202.6544, 203.5916, 203.3743, 204.1598, 
    196.2407, 196.7092, 196.6678, 197.1588, 197.5226, 198.3126, 199.5847, 
    199.1056, 199.9857, 200.1627, 198.8259, 199.646, 197.0231, 197.4453, 
    197.1938, 196.2776, 199.2161, 197.7041, 200.5026, 199.6785, 202.0906, 
    200.8885, 203.2547, 204.2728, 205.2339, 206.3619, 196.9651, 196.6464, 
    197.2173, 198.0093, 198.746, 199.7288, 199.8294, 200.0141, 200.4927, 
    200.8958, 200.0726, 200.9969, 197.5435, 199.3477, 196.5261, 197.3727, 
    197.9625, 197.7035, 199.0509, 199.3694, 200.6679, 199.9958, 204.0213, 
    202.233, 207.2234, 205.8199, 196.5351, 196.964, 198.462, 197.7482, 
    199.7944, 200.3006, 200.7126, 201.2404, 201.2973, 201.6106, 201.0975, 
    201.5903, 199.7309, 200.5602, 198.2902, 198.841, 198.5875, 198.3097, 
    199.168, 200.0855, 200.105, 200.3999, 201.2331, 199.8027, 204.2533, 
    201.4965, 197.4324, 198.2621, 198.3806, 198.0587, 200.2498, 199.4539, 
    201.6029, 201.0204, 201.9755, 201.5005, 201.4307, 200.8219, 200.4437, 
    199.4903, 198.7171, 198.1054, 198.2475, 198.9198, 200.1417, 201.3026, 
    201.0479, 201.9028, 199.6455, 200.5899, 200.2245, 201.1781, 199.0929, 
    200.8681, 198.6411, 198.8356, 199.4381, 200.6541, 200.9237, 201.2121, 
    201.034, 200.1728, 200.0318, 199.4234, 199.2557, 198.7932, 198.411, 
    198.7602, 199.1275, 200.173, 201.1188, 202.1537, 202.4074, 203.6231, 
    202.6333, 204.2688, 202.8781, 205.2897, 200.971, 202.8369, 199.4655, 
    199.8266, 200.4813, 201.9884, 201.1736, 202.1267, 200.0263, 198.9431, 
    198.6634, 198.1426, 198.6753, 198.6319, 199.1426, 198.9784, 200.2078, 
    199.5467, 201.429, 202.1191, 204.0774, 205.2849, 206.5191, 207.0659, 
    207.2325, 207.3022,
  318.6083, 320.4049, 320.0548, 321.5094, 320.7017, 321.6553, 318.9716, 
    320.4765, 319.515, 318.7695, 324.3503, 321.5744, 327.2197, 325.4688, 
    329.848, 326.9504, 330.4352, 329.7638, 331.7881, 331.2069, 333.8099, 
    332.0567, 335.1668, 333.3903, 333.6677, 331.9991, 322.131, 324.0035, 
    322.0204, 322.2867, 322.1672, 320.7184, 319.9908, 318.4712, 318.7465, 
    319.8628, 322.4066, 321.5408, 323.7265, 323.677, 326.1265, 325.0199, 
    329.0616, 327.919, 331.2312, 330.3952, 331.1919, 330.9501, 331.1951, 
    329.9698, 330.4942, 329.4179, 325.2269, 326.4759, 322.7432, 320.512, 
    319.0375, 317.9952, 318.1424, 318.4232, 319.8693, 321.2344, 322.2784, 
    322.9786, 323.6699, 325.7713, 326.8639, 329.2932, 328.8533, 329.5987, 
    330.3121, 331.5135, 331.3154, 331.8458, 329.5789, 331.0839, 328.603, 
    329.2798, 323.8588, 321.7741, 320.8925, 320.1221, 318.2556, 319.5435, 
    319.0352, 320.2455, 321.0169, 320.6352, 322.9978, 322.0773, 326.9279, 
    324.8453, 330.2288, 328.9435, 330.5376, 329.7232, 331.1199, 329.8626, 
    332.0434, 332.5202, 332.1943, 333.4476, 329.7931, 331.192, 320.6245, 
    320.6867, 320.9767, 319.7038, 319.626, 318.4637, 319.4977, 319.939, 
    321.0616, 321.7275, 322.3617, 323.7601, 325.3287, 327.4877, 329.0267, 
    330.0623, 329.4268, 329.9878, 329.3608, 329.0673, 332.3415, 330.4991, 
    333.2671, 333.1133, 331.8585, 333.1306, 320.7304, 320.3724, 319.1326, 
    320.1025, 318.3373, 319.3243, 319.8932, 322.0967, 322.5826, 323.0339, 
    323.9269, 325.0765, 327.0707, 328.783, 330.3536, 330.2383, 330.2789, 
    330.6308, 329.7599, 330.7739, 330.9445, 330.4988, 333.0927, 332.3496, 
    333.11, 332.626, 320.4887, 321.0915, 320.7657, 321.3787, 320.9467, 
    322.8718, 323.451, 326.174, 325.0539, 326.8158, 325.2346, 325.5184, 
    326.8725, 325.3211, 328.6885, 326.4216, 330.6444, 328.3678, 330.7876, 
    330.3468, 331.0769, 331.7322, 332.5583, 334.0881, 333.7332, 335.0164, 
    321.992, 322.7776, 322.7082, 323.5319, 324.1424, 325.4692, 327.5592, 
    326.7806, 328.2112, 328.4992, 326.3262, 327.6589, 323.3042, 324.0125, 
    323.5905, 322.054, 326.9601, 324.4471, 329.0522, 327.7118, 331.6387, 
    329.6802, 333.538, 335.2011, 336.773, 338.6201, 323.2069, 322.6723, 
    323.63, 324.9597, 326.1965, 327.7934, 327.9572, 328.2574, 329.036, 
    329.6922, 328.3525, 329.8569, 324.1773, 327.174, 322.4705, 323.8908, 
    324.881, 324.4462, 326.6917, 327.2094, 329.3212, 328.2278, 334.79, 
    331.871, 340.0327, 337.7322, 322.4857, 323.205, 325.7202, 324.5211, 
    327.9002, 328.7234, 329.394, 330.2533, 330.3461, 330.8564, 330.0206, 
    330.8233, 327.7968, 329.1459, 325.4316, 326.3508, 325.9311, 325.4643, 
    326.8819, 328.3736, 328.4053, 328.8851, 330.2412, 327.9138, 335.169, 
    330.6704, 323.991, 325.3842, 325.5833, 325.0427, 328.6408, 327.3465, 
    330.844, 329.8951, 331.4511, 330.677, 330.5633, 329.572, 328.9563, 
    327.4058, 326.1489, 325.121, 325.3597, 326.4788, 328.465, 330.3546, 
    329.9398, 331.3326, 327.6581, 329.1942, 328.5997, 330.1519, 326.76, 
    329.6469, 326.0212, 326.342, 327.3209, 329.2988, 329.7376, 330.2072, 
    329.9173, 328.5155, 328.2863, 327.297, 327.0245, 326.2732, 325.6345, 
    326.2196, 326.8162, 328.516, 330.0553, 331.7416, 332.1555, 334.1394, 
    332.5238, 335.1943, 332.923, 336.8641, 329.8146, 332.856, 327.3654, 
    327.9526, 329.0175, 331.4722, 330.1445, 331.6976, 328.2773, 326.5166, 
    326.0587, 325.1835, 326.0787, 326.0058, 326.8408, 326.574, 328.5726, 
    327.4975, 330.5605, 331.6853, 334.8817, 336.8564, 338.8779, 339.7742, 
    340.0475, 340.1618,
  524.4308, 527.7018, 527.0638, 529.7164, 528.2429, 529.9828, 525.0918, 
    527.8323, 526.0807, 524.7241, 534.9113, 529.8351, 540.246, 536.9622, 
    545.2583, 539.7336, 546.3807, 545.0975, 548.97, 547.8571, 552.8487, 
    549.4846, 555.4581, 552.0427, 552.5754, 549.3741, 530.8516, 534.2762, 
    530.6496, 531.136, 530.9177, 528.2734, 526.9471, 524.1816, 524.6823, 
    526.714, 531.355, 529.7738, 533.7692, 533.6785, 538.1694, 536.1389, 
    543.7567, 541.5779, 547.9035, 546.3041, 547.8283, 547.3655, 547.8344, 
    545.491, 546.4935, 544.437, 536.5185, 538.8309, 531.9703, 527.897, 
    525.2117, 523.3092, 523.5839, 524.0942, 526.7259, 529.2146, 531.1209, 
    532.4008, 533.6655, 537.5172, 539.5689, 544.1988, 543.3593, 544.7821, 
    546.1453, 548.444, 548.0648, 549.0805, 544.7443, 547.6215, 542.8819, 
    544.1732, 534.0112, 530.1997, 528.5908, 527.1865, 523.7896, 526.1326, 
    525.2075, 527.4114, 528.8178, 528.1216, 532.4359, 530.7535, 539.6909, 
    535.8187, 545.9861, 543.5314, 546.5764, 545.0199, 547.6904, 545.2863, 
    549.459, 550.3731, 549.7483, 552.1529, 545.1534, 547.8284, 528.1022, 
    528.2156, 528.7445, 526.4244, 526.2828, 524.1679, 526.0492, 526.8529, 
    528.8994, 530.1146, 531.2729, 533.8306, 536.7051, 540.7564, 543.6901, 
    545.6678, 544.454, 545.5255, 544.3279, 543.7676, 550.0305, 546.5029, 
    551.8062, 551.511, 549.1047, 551.5443, 528.2953, 527.6426, 525.3846, 
    527.1508, 523.9382, 525.7336, 526.7695, 530.7889, 531.6767, 532.502, 
    534.1361, 536.2426, 539.9626, 543.2252, 546.2247, 546.0042, 546.0818, 
    546.7546, 545.0901, 547.0285, 547.3547, 546.5023, 551.4716, 550.0461, 
    551.5048, 550.576, 527.8547, 528.9539, 528.3596, 529.4779, 528.6898, 
    532.2053, 533.2649, 538.2571, 536.201, 539.4775, 536.5327, 537.0531, 
    539.5853, 536.6912, 543.0449, 538.7277, 546.7808, 542.4333, 547.0547, 
    546.2117, 547.6082, 548.8629, 550.4462, 553.3832, 552.7014, 555.1686, 
    530.5977, 532.0331, 531.9063, 533.413, 534.5308, 536.9629, 540.8926, 
    539.4106, 542.1349, 542.684, 538.5464, 541.0824, 532.9963, 534.2928, 
    533.5203, 530.7109, 539.752, 535.0887, 543.7388, 541.1832, 548.6838, 
    544.9378, 552.3265, 555.5241, 558.5367, 561.9857, 532.8183, 531.8407, 
    533.5925, 536.0283, 538.2999, 541.3387, 541.6507, 542.2228, 543.708, 
    544.9608, 542.4041, 545.2753, 534.5945, 540.1591, 531.4719, 534.0699, 
    535.8842, 535.0872, 539.2415, 540.2265, 544.2523, 542.1664, 554.733, 
    549.1287, 564.6298, 560.3266, 531.4997, 532.8148, 537.4235, 535.2245, 
    541.5422, 543.1115, 544.3912, 546.0329, 546.2103, 547.1863, 545.5881, 
    547.123, 541.3452, 543.9177, 536.8939, 538.5933, 537.8106, 536.9539, 
    539.6034, 542.4443, 542.5048, 543.4199, 546.0095, 541.568, 555.4623, 
    546.8303, 534.2535, 536.8068, 537.1723, 536.1807, 542.9539, 540.4876, 
    547.1624, 545.3483, 548.3245, 546.8431, 546.6256, 544.7311, 543.5558, 
    540.6005, 538.2104, 536.3243, 536.7621, 538.8365, 542.6186, 546.2266, 
    545.4337, 548.0977, 541.0811, 544.0098, 542.8756, 545.839, 539.3714, 
    544.874, 537.9761, 538.5765, 540.4388, 544.2094, 545.0474, 545.9447, 
    545.3907, 542.715, 542.278, 540.3934, 539.8746, 538.4456, 537.2663, 
    538.3438, 539.4783, 542.7159, 545.6545, 548.8809, 549.6739, 553.4818, 
    550.38, 555.5109, 551.1457, 558.7064, 545.1945, 551.0172, 540.5236, 
    541.642, 543.6725, 548.3649, 545.825, 548.7966, 542.2609, 538.9085, 
    538.0449, 536.4388, 538.0816, 537.9478, 539.5251, 539.0176, 542.8239, 
    540.7751, 546.6202, 548.7729, 554.9095, 558.6921, 562.4678, 564.1457, 
    564.6577, 564.8719,
  947.2746, 954.1471, 952.8041, 958.3976, 955.2874, 958.9606, 948.6606, 
    954.422, 950.7369, 947.8893, 969.2756, 958.6484, 980.3149, 973.5083, 
    990.7758, 979.2504, 993.1304, 990.439, 998.5795, 996.2345, 1006.787, 
    999.6654, 1012.341, 1005.077, 1006.207, 999.4322, 960.7985, 967.9678, 
    960.371, 961.4009, 960.9384, 955.3517, 952.5585, 946.7524, 947.8018, 
    952.0681, 961.8646, 958.5188, 966.9247, 966.7383, 976.0063, 971.8074, 
    987.6327, 983.0861, 996.3322, 992.9696, 996.1739, 995.2001, 996.1866, 
    991.2636, 993.3673, 989.0557, 972.5914, 977.3772, 963.1688, 954.5585, 
    948.9122, 944.9412, 945.5009, 946.5695, 952.0931, 957.3376, 961.3687, 
    964.0821, 966.7115, 974.6561, 978.9084, 988.5572, 986.8021, 989.7783, 
    992.6362, 997.4706, 996.6717, 998.8126, 989.699, 995.7386, 985.8052, 
    988.5037, 967.4224, 959.4193, 956.0211, 953.0621, 945.9316, 950.8459, 
    948.9034, 953.5356, 956.5001, 955.0318, 964.1565, 960.5909, 979.1615, 
    971.1466, 992.3021, 987.1618, 993.5416, 990.2764, 995.8837, 990.8345, 
    999.6115, 1001.542, 1000.222, 1005.311, 990.556, 996.1741, 954.9908, 
    955.23, 956.3455, 951.4593, 951.1616, 946.7238, 950.6706, 952.3602, 
    956.6722, 959.2393, 961.6908, 967.0511, 972.977, 981.3761, 987.4935, 
    991.6344, 989.0912, 991.3359, 988.8274, 987.6556, 1000.818, 993.3871, 
    1004.576, 1003.951, 998.8638, 1004.021, 955.3979, 954.0226, 949.2751, 
    952.9869, 946.2427, 950.0078, 952.1848, 960.6658, 962.5463, 964.2968, 
    967.6796, 972.0215, 979.726, 986.5219, 992.8029, 992.3401, 992.503, 
    993.9158, 990.4233, 994.4914, 995.1775, 993.3859, 1003.867, 1000.851, 
    1003.937, 1001.971, 954.4692, 956.7872, 955.5335, 957.8937, 956.23, 
    963.6674, 965.8881, 976.1879, 971.9358, 978.7186, 972.6207, 973.6962, 
    978.9424, 972.9482, 986.1454, 977.1631, 993.9708, 984.869, 994.5465, 
    992.7756, 995.7107, 998.3536, 1001.697, 1007.923, 1006.475, 1011.723, 
    960.2611, 963.3021, 963.0332, 966.1925, 968.4918, 973.5097, 981.6594, 
    978.5798, 984.2468, 985.392, 976.7875, 982.0543, 965.3362, 968.0021, 
    966.4129, 960.5007, 979.2885, 969.6414, 987.5953, 982.2642, 997.9761, 
    990.1043, 1005.679, 1012.481, 1018.962, 1026.64, 964.9684, 962.894, 
    966.5614, 971.5791, 976.2766, 982.588, 983.2377, 984.4302, 987.5309, 
    990.1523, 984.8082, 990.8115, 968.6232, 980.1341, 962.1122, 967.5433, 
    971.2818, 969.6381, 978.2289, 980.2744, 988.6692, 984.3126, 1010.795, 
    998.9143, 1032.446, 1022.94, 962.1712, 964.9611, 974.4622, 969.9213, 
    983.0117, 986.2846, 988.9598, 992.4003, 992.7728, 994.8232, 991.4673, 
    994.6901, 982.6015, 987.9694, 973.3672, 976.8845, 975.2633, 973.4911, 
    978.98, 984.892, 985.0183, 986.9288, 992.3512, 983.0654, 1012.349, 
    994.0748, 967.9211, 973.1871, 973.9426, 971.8937, 985.9556, 980.8171, 
    994.773, 990.9645, 997.2189, 994.1018, 993.6448, 989.6713, 987.2128, 
    981.0518, 976.0913, 972.1903, 973.0947, 977.3889, 985.2557, 992.8068, 
    991.1436, 996.741, 982.0516, 988.1618, 985.7921, 991.9934, 978.4984, 
    989.9706, 975.6059, 976.8497, 980.7156, 988.5793, 990.3339, 992.2152, 
    991.0534, 985.4568, 984.5452, 980.6212, 979.5432, 976.5786, 974.137, 
    976.3675, 978.7203, 985.4588, 991.6065, 998.3915, 1000.065, 1008.132, 
    1001.557, 1012.453, 1003.177, 1019.338, 990.642, 1002.905, 980.892, 
    983.2196, 987.4568, 997.3038, 991.9641, 998.2139, 984.5094, 977.538, 
    975.7482, 972.4268, 975.8245, 975.5472, 978.8174, 977.7643, 985.684, 
    981.415, 993.6335, 998.164, 1011.171, 1019.307, 1027.717, 1031.395, 
    1032.507, 1032.972,
  1829.892, 1849.354, 1845.526, 1861.551, 1852.614, 1863.175, 1833.792, 
    1850.139, 1839.657, 1831.62, 1893.773, 1862.274, 1928.095, 1906.815, 
    1960.691, 1924.742, 1968.122, 1959.632, 1985.507, 1977.993, 2012.213, 
    1989.004, 2030.648, 2006.596, 2010.304, 1988.252, 1868.495, 1889.772, 
    1867.256, 1870.244, 1868.901, 1852.798, 1844.827, 1828.426, 1831.374, 
    1843.433, 1871.592, 1861.9, 1886.59, 1886.023, 1914.58, 1901.557, 
    1950.848, 1936.76, 1978.305, 1967.613, 1977.799, 1974.694, 1977.839, 
    1962.227, 1968.872, 1955.294, 1903.977, 1918.864, 1875.391, 1850.529, 
    1834.501, 1823.355, 1824.92, 1827.913, 1843.505, 1858.497, 1870.15, 
    1878.058, 1885.941, 1910.377, 1923.666, 1953.735, 1948.261, 1957.558, 
    1966.558, 1981.947, 1979.39, 1986.257, 1957.31, 1976.41, 1945.164, 
    1953.567, 1888.107, 1864.501, 1854.716, 1846.26, 1826.125, 1839.966, 
    1834.476, 1847.61, 1856.09, 1851.882, 1878.276, 1867.893, 1924.462, 
    1899.52, 1965.502, 1949.381, 1969.424, 1959.122, 1976.873, 1960.876, 
    1988.83, 1995.074, 1990.801, 2007.362, 1960, 1977.8, 1851.765, 1852.45, 
    1855.647, 1841.705, 1840.861, 1828.346, 1839.47, 1844.264, 1856.585, 
    1863.981, 1871.086, 1886.975, 1905.17, 1931.448, 1950.414, 1963.395, 
    1955.405, 1962.454, 1954.58, 1950.92, 1992.729, 1968.935, 2004.955, 
    2002.911, 1986.422, 2003.141, 1852.931, 1848.999, 1835.525, 1846.047, 
    1826.997, 1837.594, 1843.765, 1868.11, 1873.576, 1878.687, 1888.892, 
    1902.217, 1926.239, 1947.39, 1967.085, 1965.622, 1966.137, 1970.611, 
    1959.583, 1972.439, 1974.622, 1968.931, 2002.637, 1992.835, 2002.867, 
    1996.467, 1850.274, 1856.915, 1853.319, 1860.098, 1855.315, 1876.846, 
    1883.437, 1915.147, 1901.953, 1923.07, 1904.068, 1907.397, 1923.773, 
    1905.081, 1946.22, 1918.194, 1970.786, 1942.264, 1972.614, 1966.999, 
    1976.321, 1984.781, 1995.576, 2015.958, 2011.183, 2028.584, 1866.937, 
    1875.78, 1874.995, 1884.362, 1891.373, 1906.819, 1932.345, 1922.634, 
    1940.34, 1943.883, 1917.019, 1933.586, 1881.762, 1889.876, 1885.032, 
    1867.631, 1924.862, 1894.894, 1950.732, 1934.231, 1983.569, 1958.581, 
    2008.57, 2031.12, 2053.035, 2079.24, 1880.653, 1874.589, 1885.484, 
    1900.853, 1915.423, 1935.226, 1937.226, 1940.906, 1950.531, 1958.732, 
    1942.075, 1960.804, 1891.775, 1927.525, 1872.312, 1888.476, 1899.937, 
    1894.884, 1921.532, 1927.967, 1954.085, 1940.543, 2025.486, 1986.584, 
    2099.509, 2066.706, 1872.484, 1880.632, 1909.774, 1895.753, 1936.53, 
    1946.653, 1954.994, 1965.813, 1966.99, 1973.494, 1962.869, 1973.071, 
    1935.268, 1951.898, 1906.378, 1917.322, 1912.265, 1906.762, 1923.891, 
    1942.335, 1942.726, 1948.656, 1965.657, 1936.696, 2030.678, 1971.116, 
    1889.629, 1905.82, 1908.161, 1901.823, 1945.631, 1929.681, 1973.334, 
    1961.285, 1981.141, 1971.202, 1969.752, 1957.223, 1949.54, 1930.422, 
    1914.845, 1902.738, 1905.534, 1918.9, 1943.461, 1967.098, 1961.849, 
    1979.611, 1933.578, 1952.499, 1945.124, 1964.528, 1922.378, 1958.162, 
    1913.332, 1917.213, 1929.36, 1953.804, 1959.302, 1965.228, 1961.565, 
    1944.084, 1941.262, 1929.062, 1925.663, 1916.366, 1908.765, 1915.707, 
    1923.075, 1944.09, 1963.307, 1984.903, 1990.294, 2016.65, 1995.122, 
    2031.025, 2000.387, 2054.321, 1960.271, 1999.501, 1929.917, 1937.171, 
    1950.3, 1981.413, 1964.435, 1984.332, 1941.151, 1919.367, 1913.776, 
    1903.469, 1914.013, 1913.149, 1923.38, 1920.076, 1944.788, 1931.571, 
    1969.716, 1984.172, 2026.741, 2054.213, 2082.9, 2095.761, 2099.725, 
    2101.389,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.536417, 4.554907, 4.551308, 4.566253, 4.557958, 4.56775, 4.540161, 
    4.555644, 4.545755, 4.538078, 4.595354, 4.56692, 4.625009, 4.606782, 
    4.652659, 4.622171, 4.658822, 4.651775, 4.673001, 4.666914, 4.694138, 
    4.675813, 4.708288, 4.689756, 4.692653, 4.675209, 4.57263, 4.591808, 
    4.571496, 4.574227, 4.573001, 4.55813, 4.55065, 4.535005, 4.537842, 
    4.549333, 4.575456, 4.566575, 4.588974, 4.588468, 4.613493, 4.602198, 
    4.644397, 4.632376, 4.667168, 4.658402, 4.666756, 4.664221, 4.666789, 
    4.653937, 4.659441, 4.648142, 4.604312, 4.617165, 4.578906, 4.556009, 
    4.54084, 4.530098, 4.531615, 4.53451, 4.5494, 4.56343, 4.574142, 
    4.581318, 4.588395, 4.609869, 4.621258, 4.646831, 4.642207, 4.650041, 
    4.65753, 4.670125, 4.66805, 4.673605, 4.649833, 4.665624, 4.639575, 
    4.64669, 4.590327, 4.568969, 4.559918, 4.552001, 4.532783, 4.546048, 
    4.540816, 4.55327, 4.561196, 4.557274, 4.581514, 4.57208, 4.621933, 
    4.600415, 4.656656, 4.643156, 4.659896, 4.651349, 4.666001, 4.652812, 
    4.675673, 4.680662, 4.677252, 4.690355, 4.652082, 4.666757, 4.557165, 
    4.557805, 4.560784, 4.547698, 4.546897, 4.534927, 4.545577, 4.550117, 
    4.561656, 4.568491, 4.574996, 4.589318, 4.605351, 4.627834, 4.64403, 
    4.654909, 4.648236, 4.654127, 4.647542, 4.644457, 4.678792, 4.659492, 
    4.688469, 4.686862, 4.673738, 4.687043, 4.558253, 4.554574, 4.541818, 
    4.551799, 4.533625, 4.543792, 4.549646, 4.572278, 4.57726, 4.581884, 
    4.591025, 4.602776, 4.623439, 4.641468, 4.657966, 4.656756, 4.657182, 
    4.660873, 4.651734, 4.662374, 4.664163, 4.65949, 4.686647, 4.678878, 
    4.686828, 4.681768, 4.55577, 4.561963, 4.558616, 4.564911, 4.560476, 
    4.580223, 4.586155, 4.61398, 4.602545, 4.620751, 4.604392, 4.607288, 
    4.621349, 4.605274, 4.640474, 4.616592, 4.661016, 4.6371, 4.662519, 
    4.657895, 4.665551, 4.672416, 4.68106, 4.697041, 4.693337, 4.706721, 
    4.571205, 4.579258, 4.578547, 4.586983, 4.593229, 4.606786, 4.628587, 
    4.62038, 4.635453, 4.638483, 4.615587, 4.629637, 4.584652, 4.591901, 
    4.587583, 4.571841, 4.622272, 4.596344, 4.644299, 4.630195, 4.671437, 
    4.650897, 4.691299, 4.708645, 4.725002, 4.744172, 4.583656, 4.578179, 
    4.587987, 4.601583, 4.614218, 4.631054, 4.632779, 4.635939, 4.644129, 
    4.651023, 4.636939, 4.652752, 4.593586, 4.624527, 4.576111, 4.590655, 
    4.60078, 4.596335, 4.619443, 4.624901, 4.647126, 4.635627, 4.704361, 
    4.673869, 4.758796, 4.734963, 4.576267, 4.583636, 4.609348, 4.597102, 
    4.632179, 4.640841, 4.64789, 4.656913, 4.657887, 4.663239, 4.654471, 
    4.662892, 4.63109, 4.645284, 4.606402, 4.615846, 4.6115, 4.606736, 
    4.621449, 4.637161, 4.637495, 4.642541, 4.656785, 4.632321, 4.70831, 
    4.661288, 4.591681, 4.605917, 4.607951, 4.602431, 4.639973, 4.626347, 
    4.663109, 4.653153, 4.669472, 4.661358, 4.660166, 4.64976, 4.64329, 
    4.626971, 4.613721, 4.603231, 4.605669, 4.617197, 4.638123, 4.657977, 
    4.653623, 4.668231, 4.62963, 4.645791, 4.639541, 4.655849, 4.620163, 
    4.650546, 4.612419, 4.615753, 4.626076, 4.64689, 4.6515, 4.656429, 
    4.653387, 4.638654, 4.636243, 4.625824, 4.622952, 4.615027, 4.608474, 
    4.614461, 4.620756, 4.63866, 4.654836, 4.672514, 4.676846, 4.697576, 
    4.680699, 4.708573, 4.684873, 4.725947, 4.652308, 4.684173, 4.626545, 
    4.63273, 4.643933, 4.669693, 4.655772, 4.672053, 4.636148, 4.617596, 
    4.612801, 4.603869, 4.613005, 4.612262, 4.621015, 4.618201, 4.639255, 
    4.627937, 4.660136, 4.671924, 4.705318, 4.725868, 4.746843, 4.756123, 
    4.75895, 4.760132,
  5.625772, 5.649026, 5.644499, 5.663298, 5.652863, 5.665181, 5.630479, 
    5.649951, 5.637515, 5.627861, 5.699914, 5.664137, 5.737241, 5.714297, 
    5.772058, 5.733668, 5.77982, 5.770945, 5.797681, 5.790012, 5.824312, 
    5.801223, 5.842145, 5.818791, 5.822441, 5.800463, 5.671321, 5.695451, 
    5.669894, 5.67333, 5.671788, 5.653079, 5.643671, 5.623995, 5.627563, 
    5.642015, 5.674875, 5.663703, 5.691885, 5.691248, 5.722744, 5.708528, 
    5.761653, 5.746517, 5.790332, 5.779291, 5.789814, 5.786621, 5.789855, 
    5.773668, 5.7806, 5.76637, 5.711188, 5.727366, 5.679216, 5.650411, 
    5.631332, 5.617825, 5.619733, 5.623373, 5.642099, 5.659746, 5.673223, 
    5.682251, 5.691156, 5.718182, 5.732519, 5.764719, 5.758895, 5.768761, 
    5.778193, 5.794058, 5.791444, 5.798442, 5.768498, 5.788387, 5.755581, 
    5.764541, 5.693588, 5.666715, 5.655329, 5.64537, 5.621201, 5.637883, 
    5.631303, 5.646966, 5.656937, 5.652003, 5.682498, 5.670628, 5.733369, 
    5.706283, 5.777092, 5.76009, 5.781173, 5.770408, 5.788863, 5.772251, 
    5.801047, 5.807332, 5.803037, 5.819546, 5.771332, 5.789814, 5.651865, 
    5.65267, 5.656417, 5.639957, 5.638951, 5.623898, 5.63729, 5.643001, 
    5.657514, 5.666113, 5.674296, 5.692318, 5.712496, 5.740798, 5.761191, 
    5.774891, 5.766487, 5.773907, 5.765614, 5.761729, 5.804977, 5.780665, 
    5.817169, 5.815145, 5.798609, 5.815373, 5.653234, 5.648607, 5.632564, 
    5.645116, 5.62226, 5.635046, 5.642408, 5.670878, 5.677145, 5.682964, 
    5.694466, 5.709254, 5.735265, 5.757965, 5.778742, 5.777218, 5.777754, 
    5.782404, 5.770894, 5.784295, 5.786547, 5.780661, 5.814874, 5.805085, 
    5.815102, 5.808726, 5.650111, 5.6579, 5.65369, 5.66161, 5.65603, 
    5.680873, 5.688337, 5.723357, 5.708963, 5.731881, 5.711288, 5.714933, 
    5.732633, 5.712399, 5.756713, 5.726645, 5.782585, 5.752465, 5.784476, 
    5.778652, 5.788296, 5.796944, 5.807835, 5.827971, 5.823303, 5.84017, 
    5.669528, 5.679659, 5.678765, 5.68938, 5.69724, 5.714302, 5.741746, 
    5.731414, 5.750391, 5.754206, 5.725379, 5.743068, 5.686446, 5.695568, 
    5.690135, 5.670327, 5.733796, 5.70116, 5.761529, 5.74377, 5.795711, 
    5.769839, 5.820735, 5.842595, 5.863214, 5.887383, 5.685193, 5.678302, 
    5.690643, 5.707752, 5.723656, 5.744852, 5.747023, 5.751002, 5.761315, 
    5.769998, 5.752262, 5.772176, 5.697689, 5.736634, 5.6757, 5.694001, 
    5.706742, 5.701149, 5.730234, 5.737105, 5.76509, 5.75061, 5.837196, 
    5.798774, 5.905828, 5.875772, 5.675896, 5.685168, 5.717526, 5.702113, 
    5.746268, 5.757176, 5.766052, 5.777416, 5.778643, 5.785385, 5.77434, 
    5.784947, 5.744897, 5.76277, 5.713819, 5.725706, 5.720235, 5.714239, 
    5.732759, 5.752541, 5.752962, 5.759316, 5.777255, 5.746448, 5.842174, 
    5.782926, 5.695291, 5.713209, 5.715768, 5.708821, 5.756082, 5.738925, 
    5.78522, 5.772681, 5.793235, 5.783015, 5.781513, 5.768407, 5.76026, 
    5.739711, 5.723031, 5.709827, 5.712895, 5.727406, 5.753752, 5.778755, 
    5.773272, 5.791671, 5.743058, 5.763408, 5.755538, 5.776075, 5.73114, 
    5.769397, 5.721392, 5.725589, 5.738585, 5.764792, 5.770598, 5.776806, 
    5.772974, 5.754422, 5.751385, 5.738268, 5.734651, 5.724675, 5.716426, 
    5.723963, 5.731886, 5.754428, 5.774799, 5.797067, 5.802525, 5.828645, 
    5.80738, 5.842505, 5.812638, 5.864406, 5.771616, 5.811756, 5.739176, 
    5.746963, 5.761069, 5.793513, 5.775979, 5.796487, 5.751266, 5.727908, 
    5.721873, 5.71063, 5.72213, 5.721194, 5.732213, 5.72867, 5.755178, 
    5.740928, 5.781476, 5.796324, 5.838402, 5.864305, 5.890752, 5.902456, 
    5.906021, 5.907512,
  8.093964, 8.128147, 8.121491, 8.149132, 8.133788, 8.151902, 8.100883, 
    8.129508, 8.111224, 8.097034, 8.202996, 8.150367, 8.257939, 8.224163, 
    8.309218, 8.252678, 8.320656, 8.307579, 8.346976, 8.335674, 8.386237, 
    8.352197, 8.412537, 8.378096, 8.383477, 8.351077, 8.160933, 8.196429, 
    8.158834, 8.163887, 8.161618, 8.134107, 8.120274, 8.091353, 8.096597, 
    8.117839, 8.16616, 8.149729, 8.191184, 8.190246, 8.236597, 8.215672, 
    8.293891, 8.271598, 8.336146, 8.319876, 8.335382, 8.330677, 8.335443, 
    8.311591, 8.321804, 8.300838, 8.219588, 8.243402, 8.172545, 8.130183, 
    8.102137, 8.082286, 8.08509, 8.090438, 8.117964, 8.14391, 8.16373, 
    8.17701, 8.190111, 8.229882, 8.250986, 8.298407, 8.289829, 8.304361, 
    8.318258, 8.341637, 8.337785, 8.348098, 8.303975, 8.33328, 8.284947, 
    8.298145, 8.193688, 8.154159, 8.137414, 8.122771, 8.087246, 8.111766, 
    8.102093, 8.125118, 8.139778, 8.132524, 8.177373, 8.159914, 8.252239, 
    8.212368, 8.316636, 8.291589, 8.322648, 8.306787, 8.333981, 8.309504, 
    8.351938, 8.361202, 8.354871, 8.37921, 8.308148, 8.335382, 8.132322, 
    8.133505, 8.139015, 8.114815, 8.113336, 8.09121, 8.110894, 8.119289, 
    8.140628, 8.153274, 8.165308, 8.19182, 8.221513, 8.263176, 8.293211, 
    8.313394, 8.301012, 8.311942, 8.299725, 8.294003, 8.357731, 8.3219, 
    8.375705, 8.37272, 8.348344, 8.373056, 8.134336, 8.127531, 8.103946, 
    8.122398, 8.088803, 8.107595, 8.118419, 8.160281, 8.169498, 8.178058, 
    8.194981, 8.216742, 8.25503, 8.288458, 8.319067, 8.316821, 8.317612, 
    8.324462, 8.307503, 8.327249, 8.330567, 8.321894, 8.37232, 8.357889, 
    8.372657, 8.363257, 8.129742, 8.141195, 8.135005, 8.14665, 8.138446, 
    8.174983, 8.185964, 8.237499, 8.216313, 8.250048, 8.219734, 8.2251, 
    8.251155, 8.22137, 8.286614, 8.24234, 8.324728, 8.280357, 8.327516, 
    8.318934, 8.333144, 8.34589, 8.361943, 8.391632, 8.384749, 8.409624, 
    8.158295, 8.173197, 8.171882, 8.187497, 8.199061, 8.22417, 8.264573, 
    8.24936, 8.277303, 8.282923, 8.240476, 8.266519, 8.183181, 8.196602, 
    8.188607, 8.159471, 8.252867, 8.204829, 8.293709, 8.267552, 8.344071, 
    8.305949, 8.380963, 8.413201, 8.44362, 8.479292, 8.181337, 8.171201, 
    8.189355, 8.214531, 8.237939, 8.269147, 8.272344, 8.278203, 8.293393, 
    8.306184, 8.280059, 8.309392, 8.199721, 8.257047, 8.167374, 8.194296, 
    8.213044, 8.204813, 8.247622, 8.257739, 8.298953, 8.277626, 8.405237, 
    8.348587, 8.506523, 8.462153, 8.167662, 8.181301, 8.228916, 8.206232, 
    8.271232, 8.287296, 8.300371, 8.317113, 8.31892, 8.328855, 8.312581, 
    8.32821, 8.269214, 8.295536, 8.223459, 8.240957, 8.232903, 8.224077, 
    8.251341, 8.28047, 8.28109, 8.290449, 8.316875, 8.271496, 8.412579, 
    8.325232, 8.196195, 8.222561, 8.226328, 8.216104, 8.285685, 8.260419, 
    8.328611, 8.310137, 8.340424, 8.325363, 8.323149, 8.303841, 8.291838, 
    8.261577, 8.237019, 8.217586, 8.2221, 8.24346, 8.282254, 8.319086, 
    8.311007, 8.338119, 8.266505, 8.296476, 8.284883, 8.315138, 8.248957, 
    8.305299, 8.234607, 8.240785, 8.259918, 8.298514, 8.307068, 8.316215, 
    8.310569, 8.28324, 8.278768, 8.259451, 8.254127, 8.239439, 8.227297, 
    8.238391, 8.250055, 8.28325, 8.313257, 8.346072, 8.354116, 8.392627, 
    8.361272, 8.413068, 8.369024, 8.445378, 8.308567, 8.367723, 8.260788, 
    8.272255, 8.293031, 8.340833, 8.314995, 8.345217, 8.278592, 8.244199, 
    8.235314, 8.218766, 8.235693, 8.234315, 8.250536, 8.24532, 8.284353, 
    8.263369, 8.323094, 8.344976, 8.407016, 8.44523, 8.484264, 8.501545, 
    8.506809, 8.509011,
  12.66567, 12.72113, 12.71033, 12.7552, 12.73029, 12.7597, 12.67689, 
    12.72334, 12.69367, 12.67065, 12.8427, 12.7572, 12.93205, 12.87711, 
    13.01552, 12.92349, 13.03415, 13.01285, 13.07704, 13.05862, 13.14106, 
    13.08555, 13.18397, 13.12778, 13.13656, 13.08372, 12.77436, 12.83203, 
    12.77095, 12.77916, 12.77547, 12.73081, 12.70835, 12.66144, 12.66994, 
    12.7044, 12.78285, 12.75617, 12.8235, 12.82198, 12.89733, 12.8633, 
    12.99056, 12.95427, 13.05939, 13.03288, 13.05815, 13.05048, 13.05825, 
    13.01939, 13.03602, 13.00188, 12.86967, 12.9084, 12.79322, 12.72444, 
    12.67893, 12.64673, 12.65128, 12.65995, 12.70461, 12.74672, 12.7789, 
    12.80047, 12.82176, 12.88641, 12.92074, 12.99791, 12.98395, 13.00761, 
    13.03025, 13.06834, 13.06206, 13.07887, 13.00698, 13.05472, 12.976, 
    12.99749, 12.82757, 12.76336, 12.73617, 12.71241, 12.65478, 12.69455, 
    12.67886, 12.71622, 12.74001, 12.72824, 12.80106, 12.77271, 12.92277, 
    12.85793, 13.02761, 12.98681, 13.0374, 13.01156, 13.05586, 13.01599, 
    13.08513, 13.10023, 13.08991, 13.12959, 13.01378, 13.05815, 12.72791, 
    12.72983, 12.73877, 12.6995, 12.6971, 12.66121, 12.69314, 12.70676, 
    12.74139, 12.76192, 12.78147, 12.82454, 12.8728, 12.94057, 12.98946, 
    13.02232, 13.00216, 13.01996, 13.00006, 12.99074, 13.09457, 13.03618, 
    13.12388, 13.11901, 13.07927, 13.11956, 12.73118, 12.72013, 12.68186, 
    12.7118, 12.6573, 12.68779, 12.70535, 12.7733, 12.78827, 12.80218, 
    12.82967, 12.86504, 12.92731, 12.98172, 13.03156, 13.02791, 13.02919, 
    13.04035, 13.01273, 13.04489, 13.0503, 13.03617, 13.11836, 13.09483, 
    13.11891, 13.10358, 12.72372, 12.74231, 12.73226, 12.75117, 12.73785, 
    12.79718, 12.81502, 12.8988, 12.86435, 12.91921, 12.86991, 12.87863, 
    12.92101, 12.87257, 12.97872, 12.90667, 13.04079, 12.96853, 13.04533, 
    13.03135, 13.0545, 13.07527, 13.10144, 13.14986, 13.13863, 13.17922, 
    12.77008, 12.79428, 12.79214, 12.81751, 12.8363, 12.87712, 12.94284, 
    12.91809, 12.96356, 12.97271, 12.90364, 12.94601, 12.8105, 12.83231, 
    12.81932, 12.77199, 12.92379, 12.84568, 12.99026, 12.94769, 13.07231, 
    13.0102, 13.13246, 13.18505, 13.23472, 13.29299, 12.8075, 12.79104, 
    12.82053, 12.86145, 12.89951, 12.95028, 12.95549, 12.96502, 12.98975, 
    13.01058, 12.96804, 13.01581, 12.83738, 12.93059, 12.78482, 12.82856, 
    12.85903, 12.84565, 12.91526, 12.93172, 12.99881, 12.96408, 13.17206, 
    13.07967, 13.33751, 13.26499, 12.78529, 12.80744, 12.88484, 12.84796, 
    12.95368, 12.97983, 13.00111, 13.02838, 13.03133, 13.04751, 13.021, 
    13.04646, 12.95039, 12.99324, 12.87597, 12.90442, 12.89132, 12.87697, 
    12.92131, 12.96871, 12.96972, 12.98496, 13.02799, 12.95411, 13.18404, 
    13.04161, 12.83165, 12.87451, 12.88063, 12.86401, 12.9772, 12.93608, 
    13.04711, 13.01702, 13.06636, 13.04182, 13.03821, 13.00676, 12.98722, 
    12.93797, 12.89802, 12.86641, 12.87376, 12.90849, 12.97162, 13.0316, 
    13.01844, 13.06261, 12.94598, 12.99477, 12.9759, 13.02516, 12.91743, 
    13.00914, 12.89409, 12.90414, 12.93527, 12.99809, 13.01202, 13.02692, 
    13.01772, 12.97322, 12.96594, 12.93451, 12.92584, 12.90195, 12.8822, 
    12.90025, 12.91922, 12.97324, 13.0221, 13.07557, 13.08868, 13.15148, 
    13.10035, 13.18484, 13.11298, 13.23759, 13.01446, 13.11086, 12.93668, 
    12.95534, 12.98916, 13.06703, 13.02493, 13.07417, 12.96566, 12.90969, 
    12.89524, 12.86833, 12.89586, 12.89362, 12.92, 12.91152, 12.97504, 
    12.94088, 13.03813, 13.07378, 13.17496, 13.23735, 13.30112, 13.32937, 
    13.33798, 13.34158,
  20.60038, 20.69644, 20.67772, 20.7555, 20.71231, 20.7633, 20.61981, 
    20.70027, 20.64886, 20.609, 20.9074, 20.75898, 21.0628, 20.96721, 
    21.20826, 21.0479, 21.24076, 21.20361, 21.31564, 21.28347, 21.42753, 
    21.3305, 21.50263, 21.40431, 21.41966, 21.32731, 20.78874, 20.88885, 
    20.78283, 20.79706, 20.79067, 20.71321, 20.6743, 20.59305, 20.60777, 
    20.66746, 20.80347, 20.75718, 20.87405, 20.8714, 21.00238, 20.94321, 
    21.16474, 21.1015, 21.28481, 21.23855, 21.28264, 21.26926, 21.28282, 
    21.215, 21.24403, 21.18446, 20.95428, 21.02163, 20.82147, 20.70217, 
    20.62333, 20.5676, 20.57547, 20.59048, 20.6678, 20.7408, 20.79662, 
    20.83406, 20.87102, 20.98338, 21.04311, 21.17756, 21.15321, 21.19447, 
    21.23395, 21.30044, 21.28948, 21.31883, 21.19337, 21.27666, 21.13936, 
    21.17682, 20.88112, 20.76966, 20.72251, 20.68132, 20.58152, 20.65038, 
    20.62321, 20.68792, 20.72917, 20.70876, 20.83508, 20.78587, 21.04665, 
    20.93387, 21.22934, 21.15821, 21.24643, 21.20136, 21.27865, 21.20907, 
    21.32977, 21.35615, 21.33812, 21.40748, 21.20522, 21.28264, 20.70819, 
    20.71151, 20.72702, 20.65895, 20.6548, 20.59265, 20.64794, 20.67153, 
    20.73156, 20.76716, 20.80107, 20.87584, 20.95972, 21.07763, 21.16281, 
    21.22012, 21.18496, 21.216, 21.1813, 21.16506, 21.34626, 21.2443, 
    21.39749, 21.38898, 21.31953, 21.38994, 20.71385, 20.69471, 20.62841, 
    20.68027, 20.58589, 20.63867, 20.66908, 20.7869, 20.81288, 20.83702, 
    20.88477, 20.94623, 21.05456, 21.14932, 21.23625, 21.22986, 21.23211, 
    21.25159, 21.20339, 21.25951, 21.26895, 21.24428, 21.38784, 21.34671, 
    21.3888, 21.36201, 20.70093, 20.73316, 20.71573, 20.74851, 20.72542, 
    20.82834, 20.85932, 21.00493, 20.94502, 21.04045, 20.95469, 20.96986, 
    21.04358, 20.95931, 21.14409, 21.01863, 21.25234, 21.12634, 21.26027, 
    21.23587, 21.27628, 21.31254, 21.35826, 21.44293, 21.42329, 21.4943, 
    20.78131, 20.82331, 20.8196, 20.86364, 20.89629, 20.96723, 21.08159, 
    21.0385, 21.11768, 21.13362, 21.01335, 21.08711, 20.85147, 20.88934, 
    20.86678, 20.78462, 21.04843, 20.91257, 21.16422, 21.09004, 21.30737, 
    21.19898, 21.41249, 21.50453, 21.59153, 21.69375, 20.84626, 20.81768, 
    20.86889, 20.93998, 21.00618, 21.09455, 21.10362, 21.12023, 21.16333, 
    21.19964, 21.12549, 21.20876, 20.89815, 21.06027, 20.80689, 20.88283, 
    20.93578, 20.91253, 21.03358, 21.06223, 21.17911, 21.11859, 21.48177, 
    21.32022, 21.77194, 21.64461, 20.8077, 20.84616, 20.98065, 20.91654, 
    21.10047, 21.14602, 21.18314, 21.23069, 21.23583, 21.26407, 21.21782, 
    21.26224, 21.09474, 21.16941, 20.96522, 21.01472, 20.99193, 20.96697, 
    21.04411, 21.12666, 21.12842, 21.15497, 21.23002, 21.10122, 21.50275, 
    21.25377, 20.88819, 20.96268, 20.97333, 20.94443, 21.14145, 21.06982, 
    21.26338, 21.21087, 21.29699, 21.25414, 21.24785, 21.19299, 21.15891, 
    21.0731, 21.00357, 20.94861, 20.96138, 21.0218, 21.13172, 21.2363, 
    21.21334, 21.29043, 21.08707, 21.17208, 21.13918, 21.22508, 21.03736, 
    21.19713, 20.99675, 21.01423, 21.0684, 21.17786, 21.20215, 21.22814, 
    21.2121, 21.13452, 21.12183, 21.06708, 21.052, 21.01042, 20.97607, 
    21.00745, 21.04047, 21.13454, 21.21974, 21.31306, 21.33597, 21.44576, 
    21.35635, 21.50415, 21.37844, 21.59656, 21.20641, 21.37474, 21.07087, 
    21.10336, 21.1623, 21.29815, 21.22467, 21.31063, 21.12133, 21.02389, 
    20.99875, 20.95195, 20.99982, 20.99592, 21.04183, 21.02707, 21.13768, 
    21.07818, 21.2477, 21.30995, 21.48685, 21.59614, 21.70802, 21.75763, 
    21.77276, 21.77909,
  34.64215, 34.82292, 34.78766, 34.93425, 34.85282, 34.94897, 34.67868, 
    34.83013, 34.73333, 34.65836, 35.22134, 34.94081, 35.51616, 35.33468, 
    35.79315, 35.48784, 35.85518, 35.78427, 35.99827, 35.93677, 36.21262, 
    36.02671, 36.35683, 36.16808, 36.19752, 36.02061, 34.99699, 35.18624, 
    34.98582, 35.01271, 35.00064, 34.85451, 34.78121, 34.62838, 34.65605, 
    34.76833, 35.02481, 34.93742, 35.15822, 35.15321, 35.4014, 35.28918, 
    35.71017, 35.58976, 35.93933, 35.85094, 35.93518, 35.9096, 35.93551, 
    35.80601, 35.86141, 35.74776, 35.31016, 35.43795, 35.05881, 34.83371, 
    34.68531, 34.58057, 34.59535, 34.62355, 34.76899, 34.90652, 35.01187, 
    35.0826, 35.15249, 35.36535, 35.47874, 35.7346, 35.68821, 35.76683, 
    35.84217, 35.9692, 35.94825, 36.00438, 35.76474, 35.92375, 35.66182, 
    35.73318, 35.1716, 34.96096, 34.87205, 34.79444, 34.60672, 34.7362, 
    34.68507, 34.80687, 34.88459, 34.84612, 35.08454, 34.99157, 35.48547, 
    35.27149, 35.83337, 35.69772, 35.866, 35.77998, 35.92756, 35.7947, 
    36.0253, 36.07581, 36.04128, 36.17417, 35.78735, 35.93518, 34.84504, 
    34.85131, 34.88054, 34.75233, 34.7445, 34.62762, 34.73159, 34.776, 
    34.8891, 34.95626, 35.02027, 35.16162, 35.32047, 35.54436, 35.70649, 
    35.81578, 35.7487, 35.80791, 35.74173, 35.71077, 36.05688, 35.86193, 
    36.15501, 36.1387, 36.00572, 36.14054, 34.85572, 34.81965, 34.69486, 
    34.79247, 34.61493, 34.71415, 34.77139, 34.99352, 35.04259, 35.08819, 
    35.1785, 35.29491, 35.50049, 35.68079, 35.84656, 35.83437, 35.83866, 
    35.87584, 35.78386, 35.89098, 35.90901, 35.8619, 36.13652, 36.05774, 
    36.13835, 36.08703, 34.83137, 34.89211, 34.85927, 34.92107, 34.87752, 
    35.0718, 35.13036, 35.40624, 35.29262, 35.47369, 35.31094, 35.3397, 
    35.47964, 35.31971, 35.67083, 35.43225, 35.87729, 35.63703, 35.89243, 
    35.84584, 35.92302, 35.99236, 36.07986, 36.24216, 36.20448, 36.34083, 
    34.98296, 35.06228, 35.05527, 35.13854, 35.20031, 35.33472, 35.55189, 
    35.46999, 35.62054, 35.65088, 35.42223, 35.56237, 35.11551, 35.18716, 
    35.14447, 34.98921, 35.48885, 35.23115, 35.70918, 35.56795, 35.98246, 
    35.77544, 36.18376, 36.36047, 36.5279, 36.72512, 35.10567, 35.05165, 
    35.14846, 35.28307, 35.40861, 35.57654, 35.59378, 35.6254, 35.70748, 
    35.77671, 35.63542, 35.79409, 35.20383, 35.51135, 35.03127, 35.17484, 
    35.27511, 35.23106, 35.46064, 35.51508, 35.73756, 35.62228, 36.31675, 
    36.00704, 36.87632, 36.63025, 35.0328, 35.10548, 35.36017, 35.23865, 
    35.58779, 35.67451, 35.74523, 35.83596, 35.84576, 35.8997, 35.81138, 
    35.8962, 35.5769, 35.71907, 35.33091, 35.42482, 35.38157, 35.33422, 
    35.48064, 35.63764, 35.64098, 35.69156, 35.83466, 35.58921, 36.35706, 
    35.88002, 35.18499, 35.32609, 35.34629, 35.29149, 35.66581, 35.52951, 
    35.89838, 35.79813, 35.9626, 35.88073, 35.86871, 35.76402, 35.69907, 
    35.53574, 35.40366, 35.29943, 35.32362, 35.43826, 35.64727, 35.84666, 
    35.80285, 35.95006, 35.5623, 35.72415, 35.66148, 35.82524, 35.46782, 
    35.77191, 35.39071, 35.42389, 35.52681, 35.73518, 35.7815, 35.83108, 
    35.80047, 35.6526, 35.62845, 35.5243, 35.49563, 35.41666, 35.35149, 
    35.41103, 35.47373, 35.65265, 35.81505, 35.99335, 36.03717, 36.24761, 
    36.07619, 36.35974, 36.11851, 36.53761, 35.78962, 36.1114, 35.5315, 
    35.5933, 35.70552, 35.96483, 35.82447, 35.98869, 35.6275, 35.44224, 
    35.39451, 35.30576, 35.39654, 35.38914, 35.47631, 35.44827, 35.65862, 
    35.54539, 35.86842, 35.98738, 36.32651, 36.53679, 36.75269, 36.84863, 
    36.8779, 36.89016,
  60.67875, 61.07146, 60.99472, 61.31435, 61.13662, 61.34652, 60.75795, 
    61.08717, 60.87659, 60.71387, 61.94424, 61.32869, 62.59662, 62.19437, 
    63.21482, 62.53371, 63.35397, 63.19492, 63.67599, 63.53741, 64.16105, 
    63.74016, 64.48923, 64.05999, 64.12677, 63.72638, 61.45155, 61.86695, 
    61.42712, 61.48597, 61.45954, 61.1403, 60.98068, 60.64891, 60.70887, 
    60.95266, 61.51246, 61.32128, 61.8053, 61.79429, 62.342, 62.09385, 
    63.02907, 62.76039, 63.54318, 63.34447, 63.53383, 63.47628, 63.53458, 
    63.24365, 63.36797, 63.11317, 62.14018, 62.42301, 61.58699, 61.09497, 
    60.77232, 60.54541, 60.57739, 60.63845, 60.95409, 61.25378, 61.48413, 
    61.63918, 61.79271, 62.2622, 62.5135, 63.08371, 62.97999, 63.15587, 
    63.32476, 63.61046, 63.56325, 63.68977, 63.15118, 63.50811, 62.92107, 
    63.08054, 61.83472, 61.37273, 61.17855, 61.00946, 60.602, 60.88282, 
    60.77182, 61.03652, 61.20592, 61.12202, 61.64343, 61.43968, 62.52845, 
    62.05481, 63.30502, 63.00125, 63.37827, 63.1853, 63.51668, 63.21828, 
    63.73698, 63.85109, 63.77307, 64.0738, 63.20183, 63.53384, 61.11967, 
    61.13334, 61.19708, 60.91787, 60.90086, 60.64727, 60.8728, 60.96935, 
    61.21576, 61.36245, 61.50253, 61.81277, 62.16297, 62.65933, 63.02085, 
    63.26556, 63.11527, 63.24792, 63.09967, 63.03043, 63.80829, 63.36914, 
    64.03036, 63.9934, 63.69279, 63.99757, 61.14294, 61.06435, 60.79306, 
    61.00517, 60.61978, 60.83493, 60.95933, 61.44396, 61.55142, 61.65145, 
    61.84991, 62.10651, 62.56181, 62.96343, 63.33461, 63.30726, 63.31689, 
    63.40039, 63.19399, 63.4344, 63.47495, 63.36907, 63.98846, 63.81024, 
    63.99262, 63.87645, 61.08987, 61.22233, 61.15069, 61.28555, 61.19049, 
    61.61548, 61.74404, 62.35273, 62.10144, 62.50229, 62.14191, 62.20547, 
    62.51551, 62.16127, 62.94118, 62.41036, 63.40364, 62.86575, 63.43766, 
    63.333, 63.50645, 63.66264, 63.86023, 64.22816, 64.14257, 64.45275, 
    61.42084, 61.59461, 61.57924, 61.76203, 61.89791, 62.19445, 62.67607, 
    62.49408, 62.82898, 62.89666, 62.38816, 62.69941, 61.71143, 61.86897, 
    61.77505, 61.43452, 62.53596, 61.96585, 63.02687, 62.71181, 63.64033, 
    63.17514, 64.09556, 64.49754, 64.88052, 65.33427, 61.68983, 61.57129, 
    61.78383, 62.08036, 62.35797, 62.73095, 62.76934, 62.83981, 63.02306, 
    63.17798, 62.86216, 63.21693, 61.90568, 62.58593, 61.52662, 61.84186, 
    62.06279, 61.96566, 62.47334, 62.59422, 63.09032, 62.83287, 64.39787, 
    63.69578, 65.68413, 65.11563, 61.52999, 61.68941, 62.25074, 61.98239, 
    62.75599, 62.94941, 63.10751, 63.31082, 63.33283, 63.45401, 63.25569, 
    63.44614, 62.73175, 63.04897, 62.18603, 62.39389, 62.29808, 62.19336, 
    62.51773, 62.86711, 62.87457, 62.98747, 63.30792, 62.75916, 64.48975, 
    63.40977, 61.86419, 62.17539, 62.22004, 62.09895, 62.92996, 62.6263, 
    63.45104, 63.22597, 63.59559, 63.41138, 63.38437, 63.14955, 63.00426, 
    62.64016, 62.34702, 62.11648, 62.16993, 62.4237, 62.8886, 63.33485, 
    63.23655, 63.56734, 62.69925, 63.06034, 62.9203, 63.28678, 62.48927, 
    63.16724, 62.31833, 62.39183, 62.6203, 63.08502, 63.18871, 63.29988, 
    63.23122, 62.90048, 62.84661, 62.61472, 62.55101, 62.37581, 62.23153, 
    62.36334, 62.50238, 62.9006, 63.26391, 63.66488, 63.76378, 64.24053, 
    63.85195, 64.49587, 63.94768, 64.90276, 63.20691, 63.9316, 62.63072, 
    62.76827, 63.01868, 63.6006, 63.28504, 63.65438, 62.8445, 62.43251, 
    62.32674, 62.13046, 62.33125, 62.31487, 62.50812, 62.44588, 62.91391, 
    62.66163, 63.3837, 63.65144, 64.42011, 64.90089, 65.39793, 65.61993, 
    65.68781, 65.71623,
  116.3177, 117.5457, 117.3041, 118.3152, 117.7513, 118.4177, 116.5638, 
    117.5952, 116.9339, 116.4268, 120.3482, 118.3608, 122.5137, 121.1711, 
    124.6258, 122.3021, 125.1096, 124.5568, 126.2418, 125.7524, 127.9808, 
    126.4695, 129.1813, 127.6151, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9487, 118.3372, 119.895, 119.8592, 121.661, 120.8393, 
    123.9848, 123.0674, 125.7727, 125.0765, 125.7398, 125.5376, 125.7425, 
    124.7258, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9053, 116.004, 116.1928, 117.1766, 118.1225, 118.8578, 
    119.3567, 119.854, 121.3958, 122.2343, 124.1728, 123.8164, 124.4218, 
    125.0078, 126.01, 125.8434, 126.2906, 124.4056, 125.6494, 123.6147, 
    124.1619, 119.9907, 118.5013, 117.884, 117.3505, 116.0801, 116.9533, 
    116.607, 117.4356, 117.9707, 117.7052, 119.3704, 118.7153, 122.2845, 
    120.7108, 124.9391, 123.8893, 125.1945, 124.5236, 125.6795, 124.6378, 
    126.4582, 126.8648, 126.5865, 127.6649, 124.5808, 125.7399, 117.6978, 
    117.741, 117.9427, 117.063, 117.0098, 116.2202, 116.922, 117.2245, 
    118.0019, 118.4685, 118.9168, 119.9193, 121.0673, 122.7252, 123.9566, 
    124.8019, 124.2816, 124.7406, 124.2278, 123.9895, 126.712, 125.1626, 
    127.5082, 127.3751, 126.3013, 127.3901, 117.7713, 117.5232, 116.6731, 
    117.337, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.881, 122.3966, 123.7596, 125.0422, 124.9469, 124.9804, 
    125.2718, 124.5536, 125.3908, 125.5329, 125.1623, 127.3573, 126.719, 
    127.3723, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9218, 
    119.2802, 119.696, 121.6967, 120.8643, 122.1966, 120.9977, 121.2078, 
    122.241, 121.0616, 123.6834, 121.889, 125.2831, 123.4258, 125.4022, 
    125.0365, 125.6436, 126.1945, 126.8974, 128.2247, 127.9138, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1968, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8149, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3097, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4884, 127.7436, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7949, 121.7142, 122.9675, 123.0978, 123.3374, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9942, 120.014, 
    120.7371, 120.4183, 122.0996, 122.5056, 124.1956, 123.3137, 128.8452, 
    126.3119, 133.7281, 131.5293, 119.005, 119.5191, 121.3578, 120.4731, 
    123.0524, 123.7116, 124.2548, 124.9593, 125.0359, 125.4595, 124.7676, 
    125.4319, 122.9702, 124.0532, 121.1435, 121.834, 121.5149, 121.1677, 
    122.2485, 123.4304, 123.4559, 123.842, 124.9492, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1083, 121.256, 120.8561, 123.6451, 122.6137, 
    125.4491, 124.6645, 125.9575, 125.3102, 125.2158, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.043, 
    124.7012, 125.8578, 122.8602, 124.0923, 123.612, 124.8756, 122.153, 
    124.4611, 121.5822, 121.8271, 122.5935, 124.1773, 124.5353, 124.9212, 
    124.6827, 123.5443, 123.3605, 122.5747, 122.3603, 121.7737, 121.2941, 
    121.7321, 122.197, 123.5447, 124.7961, 126.2024, 126.5535, 128.2698, 
    126.8679, 129.2059, 127.2107, 130.7229, 124.5984, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9752, 124.8696, 126.1653, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5902, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6129, 133.4765, 
    133.7426, 133.8544,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02029295, -0.01996183, -0.02002575, -0.01976198, -0.01990785, 
    -0.0197358, -0.02022536, -0.01994879, -0.02012488, -0.02026292, 
    -0.01926068, -0.01975031, -0.01876604, -0.01906815, -0.01831904, 
    -0.01881269, -0.01822122, -0.01833312, -0.01799864, -0.01809378, 
    -0.01767309, -0.01795491, -0.01745925, -0.01773997, -0.01769572, 
    -0.01796428, -0.01965074, -0.01932091, -0.01967046, -0.01962301, 
    -0.01964429, -0.01990481, -0.02003748, -0.02031853, -0.0202672, 
    -0.02006094, -0.01960171, -0.01975634, -0.0193692, -0.01937785, 
    -0.01895622, -0.01914509, -0.0184512, -0.01864562, -0.0180898, 
    -0.01822787, -0.01809626, -0.01813606, -0.01809574, -0.01829869, 
    -0.01821144, -0.01839115, -0.01910955, -0.01889531, -0.01954204, 
    -0.01994232, -0.02021314, -0.02040769, -0.02038006, -0.0203275, 
    -0.02005974, -0.01981147, -0.01962449, -0.01950047, -0.0193791, 
    -0.01901656, -0.01882772, -0.01841214, -0.01848643, -0.01836079, 
    -0.01824167, -0.01804351, -0.01807597, -0.01798923, -0.01836412, 
    -0.01811402, -0.01852888, -0.0184144, -0.01934612, -0.0197145, 
    -0.01987326, -0.02001344, -0.02035885, -0.02011963, -0.02021357, 
    -0.01999088, -0.01985074, -0.01991993, -0.01949709, -0.01966031, 
    -0.01881659, -0.01917513, -0.01825552, -0.01847116, -0.01820424, 
    -0.01833992, -0.0181081, -0.0183166, -0.01795707, -0.01787979, 
    -0.01793256, -0.01773081, -0.01832823, -0.01809624, -0.01992186, 
    -0.01991056, -0.01985801, -0.02009014, -0.02010444, -0.02031993, 
    -0.02012808, -0.02004696, -0.01984266, -0.01972285, -0.01960969, 
    -0.01936334, -0.01909212, -0.01871975, -0.0184571, -0.01828326, 
    -0.01838965, -0.01829568, -0.01840076, -0.01845023, -0.0179087, 
    -0.01821062, -0.01775967, -0.01778431, -0.01798717, -0.01778153, 
    -0.01990263, -0.01996774, -0.02019553, -0.02001702, -0.02034355, 
    -0.02016006, -0.02005536, -0.01965686, -0.01957048, -0.01949072, 
    -0.01933423, -0.01913537, -0.01879182, -0.01849834, -0.01823477, 
    -0.01825394, -0.01824719, -0.01818881, -0.01833377, -0.01816513, 
    -0.01813698, -0.01821067, -0.01778761, -0.01790738, -0.01778484, 
    -0.01786271, -0.01994655, -0.01983726, -0.01989624, -0.01978549, 
    -0.01986343, -0.01951933, -0.01941741, -0.01894813, -0.01913926, 
    -0.01883608, -0.01910823, -0.01905969, -0.01882622, -0.01909342, 
    -0.01851437, -0.0189048, -0.01818655, -0.01856891, -0.01816287, 
    -0.0182359, -0.01811517, -0.01800776, -0.01787363, -0.01762895, 
    -0.01768529, -0.01748277, -0.01967554, -0.01953597, -0.01954823, 
    -0.01940323, -0.01929673, -0.01906809, -0.01870743, -0.01884219, 
    -0.01859562, -0.01854653, -0.01892147, -0.01869028, -0.01944317, 
    -0.01931933, -0.01939298, -0.01966448, -0.01881102, -0.0192439, 
    -0.01845278, -0.01868118, -0.01802303, -0.01834713, -0.01771638, 
    -0.0174539, -0.0172108, -0.01693126, -0.01946027, -0.01955459, 
    -0.01938607, -0.01915545, -0.01894418, -0.01866716, -0.01863907, 
    -0.01858774, -0.01845551, -0.01834511, -0.01857152, -0.01831755, 
    -0.01929068, -0.01877395, -0.01959036, -0.01934053, -0.01916897, 
    -0.01924405, -0.01885767, -0.01876782, -0.01840742, -0.01859279, 
    -0.01751827, -0.01798513, -0.01672178, -0.01706482, -0.01958765, 
    -0.0194606, -0.01902526, -0.01923108, -0.01864883, -0.01850844, 
    -0.01839518, -0.01825145, -0.01823602, -0.01815151, -0.01829021, 
    -0.01815697, -0.01866657, -0.01843696, -0.01907451, -0.01891716, 
    -0.01898938, -0.01906893, -0.01882458, -0.01856793, -0.01856252, 
    -0.01848105, -0.01825348, -0.01864651, -0.01745891, -0.01818226, 
    -0.01932307, -0.01908264, -0.0190486, -0.01914117, -0.01852247, 
    -0.01874411, -0.01815357, -0.01831117, -0.01805372, -0.01818115, 
    -0.01819998, -0.01836528, -0.018469, -0.01873388, -0.01895243, 
    -0.01912772, -0.01908681, -0.0188948, -0.01855236, -0.0182346, 
    -0.0183037, -0.01807315, -0.0186904, -0.01842883, -0.01852944, 
    -0.01826833, -0.01884578, -0.01835272, -0.01897408, -0.01891871, 
    -0.01874854, -0.0184112, -0.01833752, -0.01825912, -0.01830746, 
    -0.01854376, -0.01858281, -0.01875266, -0.01879984, -0.01893075, 
    -0.01903987, -0.01894014, -0.018836, -0.01854368, -0.01828442, 
    -0.01800623, -0.01793887, -0.01762083, -0.01787921, -0.01745497, 
    -0.01781488, -0.01719688, -0.01832463, -0.01782565, -0.01874084, 
    -0.01863986, -0.01845865, -0.01805028, -0.01826955, -0.01801341, 
    -0.01858434, -0.01888819, -0.01896773, -0.019117, -0.01896433, 
    -0.0189767, -0.01883173, -0.01887819, -0.01853406, -0.01871806, 
    -0.01820045, -0.01801542, -0.01750387, -0.01719805, -0.01689275, 
    -0.01675983, -0.0167196, -0.01670282,
  -0.05425788, -0.0532087, -0.053411, -0.05257698, -0.05303796, -0.05249428, 
    -0.05404347, -0.05316745, -0.05372497, -0.05416261, -0.05099726, 
    -0.0525401, -0.04944564, -0.05039249, -0.04804965, -0.04959168, 
    -0.04774494, -0.04809352, -0.04705269, -0.04734841, -0.04604295, 
    -0.04691686, -0.04538146, -0.04625013, -0.04611304, -0.04694597, 
    -0.05222581, -0.05118667, -0.05228804, -0.05213833, -0.05220548, 
    -0.05302836, -0.05344814, -0.05433904, -0.05417616, -0.05352242, 
    -0.05207116, -0.05255916, -0.05133863, -0.05136586, -0.05004137, 
    -0.05063403, -0.04846177, -0.04906898, -0.04733603, -0.04776564, 
    -0.0473561, -0.04747991, -0.04735449, -0.04798624, -0.04771448, 
    -0.04827442, -0.05052245, -0.04985047, -0.05188303, -0.05314698, 
    -0.05400471, -0.05462212, -0.05453438, -0.05436752, -0.05351862, 
    -0.05273332, -0.05214299, -0.05175199, -0.05136978, -0.05023062, 
    -0.04963875, -0.04833991, -0.04857171, -0.04817978, -0.04780861, 
    -0.04719213, -0.04729303, -0.04702347, -0.04819015, -0.04741137, 
    -0.04870425, -0.04834696, -0.05126601, -0.05242705, -0.05292859, 
    -0.05337204, -0.05446702, -0.05370833, -0.05400606, -0.05330065, 
    -0.05285741, -0.05307616, -0.05174135, -0.05225601, -0.0496039, 
    -0.0507284, -0.04785175, -0.04852404, -0.04769209, -0.04811473, 
    -0.04739293, -0.04804203, -0.04692359, -0.04668369, -0.04684748, 
    -0.04622173, -0.04807827, -0.04735607, -0.05308228, -0.05304654, 
    -0.05288037, -0.05361489, -0.0536602, -0.05434349, -0.05373508, 
    -0.05347815, -0.05283187, -0.05245341, -0.05209631, -0.05132018, 
    -0.05046773, -0.04930081, -0.04848016, -0.04793815, -0.04826976, 
    -0.04797687, -0.0483044, -0.04845874, -0.0467734, -0.04771193, 
    -0.04631118, -0.04638755, -0.04701707, -0.04637894, -0.05302146, 
    -0.0532274, -0.05394887, -0.05338339, -0.05441846, -0.05383644, 
    -0.05350474, -0.05224512, -0.05197268, -0.05172127, -0.05122859, 
    -0.05060351, -0.04952634, -0.0486089, -0.04778713, -0.04784684, 
    -0.04782581, -0.04764406, -0.04809556, -0.04757036, -0.04748278, 
    -0.04771208, -0.04639779, -0.04676931, -0.04638917, -0.04663068, 
    -0.05316037, -0.0528148, -0.05300124, -0.05265121, -0.05289752, 
    -0.05181142, -0.0514904, -0.050016, -0.05061572, -0.0496649, -0.05051829, 
    -0.05036593, -0.04963405, -0.05047181, -0.04865894, -0.0498802, 
    -0.047637, -0.04882928, -0.04756332, -0.04779065, -0.04741492, 
    -0.04708103, -0.04666458, -0.04590628, -0.04608072, -0.04545414, 
    -0.05230406, -0.05186387, -0.05190254, -0.05144575, -0.05111064, 
    -0.05039229, -0.04926227, -0.04968406, -0.04891271, -0.04875937, 
    -0.04993243, -0.04920863, -0.05157151, -0.0511817, -0.05141347, 
    -0.05226915, -0.04958643, -0.05094451, -0.0484667, -0.04918016, 
    -0.04712848, -0.04813718, -0.04617703, -0.04536491, -0.04461471, 
    -0.04375433, -0.05162536, -0.05192257, -0.05139173, -0.05066659, 
    -0.05000363, -0.04913632, -0.04904852, -0.0488881, -0.04847522, 
    -0.04813091, -0.04883743, -0.04804501, -0.0510916, -0.04947039, 
    -0.05203534, -0.05124842, -0.05070907, -0.050945, -0.04973252, 
    -0.04945119, -0.04832518, -0.04890388, -0.04556387, -0.04701073, 
    -0.04311126, -0.04416511, -0.05202682, -0.05162641, -0.05025791, 
    -0.05090421, -0.04907903, -0.04864043, -0.048287, -0.04783906, 
    -0.04779101, -0.04752797, -0.0479598, -0.04754497, -0.04913449, 
    -0.04841733, -0.05041245, -0.04991894, -0.05014536, -0.05039492, 
    -0.04962889, -0.0488262, -0.04880931, -0.04855492, -0.04784539, 
    -0.04907178, -0.04538041, -0.04762368, -0.05119348, -0.05043795, 
    -0.05033113, -0.05062172, -0.04868421, -0.04937701, -0.04753438, 
    -0.04802511, -0.04722387, -0.04762022, -0.04767883, -0.04819376, 
    -0.0485173, -0.04934499, -0.0500295, -0.05057948, -0.05045104, 
    -0.04984885, -0.04877758, -0.04778661, -0.04800183, -0.04728426, 
    -0.04920901, -0.04839196, -0.048706, -0.04789165, -0.04969529, 
    -0.04815463, -0.05009736, -0.04992379, -0.04939087, -0.04833699, 
    -0.04810722, -0.04786297, -0.04801355, -0.04875072, -0.04887268, 
    -0.04940378, -0.04955143, -0.04996153, -0.05030372, -0.04999095, 
    -0.04966468, -0.04875045, -0.04794176, -0.04707628, -0.04686705, 
    -0.04588116, -0.04668189, -0.04536822, -0.04648232, -0.0445718, 
    -0.04806707, -0.04651573, -0.0493668, -0.04905097, -0.04848502, 
    -0.04721316, -0.04789545, -0.04709858, -0.04887747, -0.04982816, 
    -0.05007744, -0.05054584, -0.05006679, -0.05010558, -0.04965129, 
    -0.0497968, -0.0487204, -0.04929551, -0.04768027, -0.04710485, 
    -0.04551935, -0.0445754, -0.04363602, -0.04322796, -0.04310458, -0.0430531,
  -0.07889416, -0.07723925, -0.07755817, -0.07624393, -0.07697016, 
    -0.07611369, -0.07855578, -0.07717424, -0.0780533, -0.07874379, 
    -0.07375871, -0.07618586, -0.07132304, -0.07280873, -0.06913635, 
    -0.07155206, -0.06865965, -0.06920501, -0.06757747, -0.06803963, 
    -0.06600105, -0.06736527, -0.06496966, -0.06632429, -0.06611039, 
    -0.06741075, -0.075691, -0.07405642, -0.07578897, -0.07555331, 
    -0.07565899, -0.07695502, -0.07761673, -0.07902227, -0.07876518, 
    -0.07773386, -0.07544759, -0.07621587, -0.0742953, -0.07433811, 
    -0.07225756, -0.07318804, -0.06978144, -0.0707326, -0.06802028, 
    -0.06869203, -0.06805165, -0.06824519, -0.06804913, -0.06903714, 
    -0.068612, -0.06948813, -0.07301281, -0.07195801, -0.07515153, 
    -0.07714198, -0.07849462, -0.07946923, -0.07933069, -0.07906725, 
    -0.07772787, -0.07649017, -0.07556064, -0.07494538, -0.07434427, 
    -0.0725546, -0.07162589, -0.06959065, -0.06995358, -0.06934, -0.06875924, 
    -0.06779537, -0.06795307, -0.06753182, -0.06935622, -0.06813804, 
    -0.07016116, -0.06960168, -0.07418114, -0.07600784, -0.07679782, 
    -0.07749674, -0.07922433, -0.07802705, -0.07849675, -0.07738419, 
    -0.07668567, -0.07703035, -0.07492863, -0.07573855, -0.07157123, 
    -0.07333627, -0.06882672, -0.06987894, -0.06857699, -0.06923819, 
    -0.06810923, -0.06912442, -0.06737579, -0.0670011, -0.06725691, 
    -0.06627998, -0.06918114, -0.06805161, -0.07704, -0.07698367, 
    -0.07672185, -0.07787968, -0.07795113, -0.0790293, -0.07806925, 
    -0.07766405, -0.07664543, -0.07604934, -0.07548718, -0.07426629, 
    -0.07292687, -0.07109598, -0.06981023, -0.06896189, -0.06948084, 
    -0.06902246, -0.06953505, -0.06977669, -0.06714121, -0.06860802, 
    -0.06641957, -0.06653877, -0.06752182, -0.06652533, -0.07694415, 
    -0.07726873, -0.07840652, -0.07751463, -0.07914765, -0.07822914, 
    -0.07770597, -0.0757214, -0.0752926, -0.07489706, -0.0741223, 
    -0.07314011, -0.0714496, -0.07001182, -0.06872563, -0.06881905, 
    -0.06878614, -0.06850187, -0.06920819, -0.06838664, -0.0682497, 
    -0.06860826, -0.06655475, -0.06713482, -0.06654131, -0.06691833, 
    -0.07716308, -0.07661854, -0.07691228, -0.07636084, -0.07674886, 
    -0.07503888, -0.07453393, -0.07221775, -0.07315929, -0.0716669, 
    -0.07300627, -0.07276703, -0.07161853, -0.07293327, -0.0700902, 
    -0.07200465, -0.06849084, -0.07035702, -0.06837562, -0.06873114, 
    -0.0681436, -0.06762176, -0.06697126, -0.06578787, -0.06605998, 
    -0.06508294, -0.07581419, -0.0751214, -0.07518224, -0.07446373, 
    -0.07393691, -0.07280842, -0.07103556, -0.07169694, -0.07048772, 
    -0.0702475, -0.07208661, -0.07095148, -0.07466149, -0.0740486, 
    -0.07441296, -0.07575923, -0.07154383, -0.07367583, -0.06978916, 
    -0.07090686, -0.06769589, -0.06927332, -0.06621024, -0.06494386, 
    -0.0637755, -0.0624373, -0.07474618, -0.07521376, -0.07437879, 
    -0.07323919, -0.07219834, -0.07083814, -0.07070053, -0.07044917, 
    -0.0698025, -0.06926351, -0.07036978, -0.06912909, -0.07390699, 
    -0.07136186, -0.07539122, -0.07415348, -0.07330591, -0.07367658, 
    -0.07177297, -0.07133176, -0.06956759, -0.07047389, -0.06525397, 
    -0.06751193, -0.06143834, -0.06307599, -0.07537781, -0.07474785, 
    -0.07259744, -0.0736125, -0.07074834, -0.07006121, -0.06950782, 
    -0.06880687, -0.06873171, -0.06832035, -0.06899577, -0.06834694, 
    -0.07083527, -0.06971186, -0.07284008, -0.07206544, -0.07242078, 
    -0.07281255, -0.07161043, -0.0703522, -0.07032574, -0.06992729, 
    -0.06881678, -0.07073698, -0.06496803, -0.06847001, -0.07406711, 
    -0.07288011, -0.0727124, -0.07316872, -0.07012978, -0.07121544, 
    -0.06833037, -0.06909794, -0.06784497, -0.0684646, -0.06855625, 
    -0.06936188, -0.06986838, -0.07116525, -0.07223893, -0.07310237, 
    -0.07290066, -0.07195548, -0.07027602, -0.06872483, -0.06906153, 
    -0.06793936, -0.07095207, -0.06967213, -0.07016391, -0.06888915, 
    -0.07171457, -0.06930064, -0.07234544, -0.07207304, -0.07123716, 
    -0.06958608, -0.06922644, -0.06884428, -0.06907987, -0.07023396, 
    -0.070425, -0.0712574, -0.07148894, -0.07213227, -0.07266936, 
    -0.07217844, -0.07166655, -0.07023353, -0.06896754, -0.06761434, 
    -0.06728747, -0.06574869, -0.06699829, -0.06494903, -0.06668671, 
    -0.06370872, -0.06916361, -0.06673887, -0.07119942, -0.07070437, 
    -0.06981783, -0.06782823, -0.06889509, -0.06764919, -0.07043251, 
    -0.07192301, -0.07231417, -0.07304954, -0.07229745, -0.07235833, 
    -0.07164555, -0.07187381, -0.07018647, -0.07108767, -0.06855851, 
    -0.06765898, -0.06518456, -0.06371434, -0.06225343, -0.06161955, 
    -0.06142796, -0.06134805,
  -0.08614223, -0.08423331, -0.08460107, -0.08308587, -0.08392303, 
    -0.08293578, -0.08575179, -0.08415834, -0.08517212, -0.08596871, 
    -0.08022315, -0.08301895, -0.07742072, -0.07912973, -0.07490762, 
    -0.07768407, -0.07436012, -0.07498647, -0.07311773, -0.07364822, 
    -0.07130922, -0.0728742, -0.07012681, -0.07167993, -0.07143461, 
    -0.07292639, -0.08244867, -0.0805659, -0.08256157, -0.08229002, 
    -0.0824118, -0.08390559, -0.0846686, -0.08629005, -0.08599339, 
    -0.08480369, -0.08216821, -0.08305354, -0.08084095, -0.08089026, 
    -0.07849555, -0.07956625, -0.0756487, -0.07674187, -0.073626, -0.0743973, 
    -0.07366203, -0.07388422, -0.07365914, -0.07479364, -0.0743054, 
    -0.07531171, -0.07936457, -0.07815098, -0.08182714, -0.08412115, 
    -0.08568123, -0.08680588, -0.08664598, -0.08634195, -0.08479677, 
    -0.0833697, -0.08229847, -0.08158967, -0.08089735, -0.07883731, 
    -0.07776898, -0.07542949, -0.07584651, -0.07514154, -0.07447448, 
    -0.07336783, -0.07354885, -0.07306535, -0.07516017, -0.0737612, 
    -0.07608505, -0.07544216, -0.08070951, -0.08281378, -0.08372435, 
    -0.08453023, -0.08652323, -0.08514185, -0.0856837, -0.08440043, 
    -0.08359506, -0.08399244, -0.08157037, -0.08250346, -0.07770612, 
    -0.07973686, -0.07455198, -0.07576074, -0.07426519, -0.07502459, 
    -0.07372813, -0.0748939, -0.07288627, -0.07245633, -0.07274985, 
    -0.07162909, -0.07495905, -0.07366197, -0.08400357, -0.08393861, 
    -0.08363676, -0.08497187, -0.08505428, -0.08629817, -0.08519053, 
    -0.08472317, -0.08354867, -0.0828616, -0.08221383, -0.08080755, 
    -0.07926568, -0.07715963, -0.07568178, -0.07470722, -0.07530333, 
    -0.07477679, -0.07536562, -0.07564325, -0.07261708, -0.07430083, 
    -0.07178921, -0.07192593, -0.07305387, -0.07191051, -0.08389305, 
    -0.08426729, -0.08557959, -0.08455085, -0.08643474, -0.08537497, 
    -0.08477152, -0.0824837, -0.08198965, -0.081534, -0.08064176, 
    -0.07951109, -0.07756625, -0.07591343, -0.07443589, -0.07454316, 
    -0.07450537, -0.07417893, -0.07499012, -0.07404662, -0.07388939, 
    -0.0743011, -0.07194426, -0.07260975, -0.07192884, -0.07236136, 
    -0.08414547, -0.08351768, -0.08385631, -0.08322064, -0.08366791, 
    -0.08169737, -0.08111577, -0.07844976, -0.07953315, -0.07781616, 
    -0.07935705, -0.07908174, -0.07776052, -0.07927304, -0.07600351, 
    -0.07820463, -0.07416628, -0.07631016, -0.07403397, -0.07444222, 
    -0.07376758, -0.07316857, -0.07242209, -0.07106477, -0.07137679, 
    -0.07025664, -0.08259062, -0.08179242, -0.0818625, -0.08103491, 
    -0.08042829, -0.07912937, -0.07709017, -0.07785071, -0.07646038, 
    -0.07618427, -0.0782989, -0.0769935, -0.08126269, -0.08055689, 
    -0.08097646, -0.0825273, -0.07767461, -0.08012772, -0.07565758, 
    -0.0769422, -0.07325365, -0.07506495, -0.07154912, -0.07009725, 
    -0.06875864, -0.06722657, -0.08136022, -0.08189882, -0.0809371, 
    -0.07962512, -0.07842743, -0.07686319, -0.076705, -0.07641607, 
    -0.0756729, -0.07505367, -0.07632482, -0.07489926, -0.08039385, 
    -0.07746536, -0.08210327, -0.08067767, -0.07970191, -0.08012859, 
    -0.07793815, -0.07743074, -0.075403, -0.07644448, -0.07045268, 
    -0.07304251, -0.06608365, -0.06795764, -0.08208782, -0.08136214, 
    -0.0788866, -0.08005481, -0.07675996, -0.07597019, -0.07533433, 
    -0.07452919, -0.07444286, -0.07397051, -0.07474613, -0.07400104, 
    -0.07685989, -0.07556875, -0.0791658, -0.07827456, -0.07868333, 
    -0.07913411, -0.0777512, -0.07630461, -0.07627419, -0.0758163, 
    -0.07454057, -0.0767469, -0.07012495, -0.07414236, -0.0805782, 
    -0.07921187, -0.07901887, -0.079544, -0.07604899, -0.07729698, 
    -0.07398202, -0.07486349, -0.07342476, -0.07413614, -0.07424138, 
    -0.07516667, -0.0757486, -0.07723927, -0.07847413, -0.07946765, 
    -0.07923551, -0.07814807, -0.07621706, -0.07443497, -0.07482167, 
    -0.07353312, -0.07699417, -0.07552311, -0.0760882, -0.07462367, 
    -0.07787098, -0.07509632, -0.07859666, -0.0782833, -0.07732197, 
    -0.07542424, -0.07501109, -0.07457215, -0.07484273, -0.07616871, 
    -0.07638829, -0.07734524, -0.07761148, -0.07835143, -0.07896934, 
    -0.07840454, -0.07781575, -0.07616822, -0.07471371, -0.07316004, 
    -0.07278492, -0.07101984, -0.0724531, -0.07010317, -0.07209565, 
    -0.06868217, -0.07493892, -0.07215548, -0.07727857, -0.07670941, 
    -0.07569052, -0.07340556, -0.0746305, -0.07320005, -0.07639692, 
    -0.07811072, -0.07856069, -0.07940684, -0.07854145, -0.07861149, 
    -0.0777916, -0.07805413, -0.07611413, -0.07715007, -0.07424398, 
    -0.07321128, -0.07037313, -0.06868859, -0.06701615, -0.06629092, 
    -0.06607177, -0.06598037,
  -0.06724078, -0.06569531, -0.06599306, -0.06476631, -0.0654441, 
    -0.06464478, -0.06692469, -0.06563461, -0.06645539, -0.06710031, 
    -0.06244846, -0.06471212, -0.06017934, -0.06156312, -0.05814446, 
    -0.06039258, -0.05770115, -0.05820831, -0.05669519, -0.05712473, 
    -0.05523086, -0.05649801, -0.05427349, -0.05553101, -0.05533239, 
    -0.05654026, -0.06425039, -0.06272598, -0.0643418, -0.06412194, 
    -0.06422054, -0.06542998, -0.06604773, -0.06736046, -0.06712029, 
    -0.0661571, -0.06402332, -0.06474012, -0.06294868, -0.0629886, 
    -0.06104964, -0.06191657, -0.05874452, -0.05962967, -0.05710674, 
    -0.05773126, -0.0571359, -0.05731582, -0.05713356, -0.05805218, 
    -0.05765685, -0.05847166, -0.06175327, -0.06077063, -0.06374717, 
    -0.0656045, -0.06686757, -0.06777807, -0.06764861, -0.06740247, 
    -0.0661515, -0.06499611, -0.06412879, -0.06355489, -0.06299434, 
    -0.06132636, -0.06046133, -0.05856703, -0.05890469, -0.05833387, 
    -0.05779376, -0.05689769, -0.05704426, -0.05665277, -0.05834896, 
    -0.05721621, -0.05909785, -0.05857729, -0.06284226, -0.064546, 
    -0.06528325, -0.0659357, -0.06754924, -0.06643087, -0.06686956, 
    -0.06583062, -0.06517857, -0.06550029, -0.06353927, -0.06429476, 
    -0.06041044, -0.06205472, -0.0578565, -0.05883524, -0.05762429, 
    -0.05823918, -0.05718943, -0.05813336, -0.05650778, -0.05615966, 
    -0.05639732, -0.05548985, -0.05818611, -0.05713586, -0.0655093, 
    -0.06545672, -0.06521232, -0.06629327, -0.06635998, -0.06736703, 
    -0.06647029, -0.06609192, -0.065141, -0.06458472, -0.06406025, 
    -0.06292164, -0.0616732, -0.05996794, -0.05877131, -0.0579822, 
    -0.05846487, -0.05803853, -0.05851531, -0.05874011, -0.05628982, 
    -0.05765314, -0.05561949, -0.05573019, -0.05664347, -0.05571771, 
    -0.06541982, -0.06572282, -0.06678528, -0.0659524, -0.0674776, 
    -0.06661961, -0.06613106, -0.06427876, -0.06387874, -0.06350981, 
    -0.06278739, -0.06187191, -0.06029718, -0.05895888, -0.0577625, 
    -0.05784936, -0.05781876, -0.05755444, -0.05821127, -0.05744731, 
    -0.05732, -0.05765336, -0.05574504, -0.05628388, -0.05573255, 
    -0.05608276, -0.06562419, -0.06511591, -0.06539008, -0.06487542, 
    -0.06523754, -0.06364209, -0.06317119, -0.06101256, -0.06188978, 
    -0.06049953, -0.06174719, -0.06152427, -0.06045448, -0.06167916, 
    -0.05903181, -0.06081408, -0.05754419, -0.05928012, -0.05743706, 
    -0.05776763, -0.05722137, -0.05673635, -0.05613193, -0.05503293, 
    -0.05528557, -0.05437861, -0.06436533, -0.06371906, -0.0637758, 
    -0.06310572, -0.06261455, -0.06156283, -0.05991169, -0.0605275, 
    -0.05940175, -0.05917818, -0.06089041, -0.05983341, -0.06329014, 
    -0.06271868, -0.06305839, -0.06431406, -0.06038492, -0.06237119, 
    -0.05875171, -0.05979188, -0.05680525, -0.05827186, -0.05542509, 
    -0.05424956, -0.05316576, -0.05192537, -0.06336912, -0.0638052, 
    -0.06302653, -0.06196424, -0.06099447, -0.0597279, -0.05959982, 
    -0.05936586, -0.05876412, -0.05826272, -0.05929198, -0.0581377, 
    -0.06258667, -0.06021548, -0.06397074, -0.06281647, -0.06202642, 
    -0.06237189, -0.0605983, -0.06018745, -0.05854558, -0.05938887, 
    -0.05453734, -0.05663428, -0.05100009, -0.05251725, -0.06395823, 
    -0.06337066, -0.06136626, -0.06231216, -0.05964432, -0.05900484, 
    -0.05848998, -0.05783805, -0.05776815, -0.05738568, -0.05801371, 
    -0.0574104, -0.05972524, -0.05867979, -0.06159233, -0.06087069, 
    -0.06120168, -0.06156668, -0.06044693, -0.05927562, -0.05925099, 
    -0.05888022, -0.05784727, -0.05963375, -0.05427199, -0.05752483, 
    -0.06273594, -0.06162963, -0.06147336, -0.06189856, -0.05906864, 
    -0.06007915, -0.057395, -0.05810873, -0.0569438, -0.05751979, 
    -0.05760501, -0.05835423, -0.05882541, -0.06003242, -0.06103228, 
    -0.06183673, -0.06164877, -0.06076828, -0.05920473, -0.05776176, 
    -0.05807487, -0.05703153, -0.05983396, -0.05864283, -0.0591004, 
    -0.05791456, -0.06054392, -0.05829727, -0.0611315, -0.06087777, 
    -0.06009938, -0.05856278, -0.05822825, -0.05787283, -0.05809192, 
    -0.05916558, -0.05934338, -0.06011822, -0.0603338, -0.06093294, 
    -0.06143326, -0.06097594, -0.0604992, -0.05916519, -0.05798746, 
    -0.05672945, -0.05642571, -0.05499656, -0.05615705, -0.05425436, 
    -0.05586762, -0.05310385, -0.05816982, -0.05591606, -0.06006424, 
    -0.05960339, -0.05877839, -0.05692824, -0.05792008, -0.05676184, 
    -0.05935036, -0.06073804, -0.06110238, -0.0617875, -0.0610868, 
    -0.06114351, -0.06047964, -0.06069221, -0.05912139, -0.05996019, 
    -0.05760711, -0.05677094, -0.05447293, -0.05310905, -0.05175501, 
    -0.05116788, -0.05099047, -0.05091648,
  -0.06388431, -0.06219237, -0.06251808, -0.06117686, -0.06191765, 
    -0.0610441, -0.063538, -0.06212598, -0.06302408, -0.06373039, 
    -0.05864837, -0.06111766, -0.05618052, -0.05768459, -0.05397406, 
    -0.05641212, -0.05349423, -0.05404319, -0.05240658, -0.0528708, 
    -0.05082632, -0.05219357, -0.04979515, -0.05114995, -0.05093577, 
    -0.05223922, -0.0606134, -0.05895071, -0.06071321, -0.06047317, 
    -0.06058081, -0.06190221, -0.06257791, -0.06401546, -0.06375229, 
    -0.06269759, -0.06036553, -0.06114825, -0.0591934, -0.05923691, 
    -0.05712614, -0.05806922, -0.05462405, -0.05558387, -0.05285135, 
    -0.05352681, -0.05288288, -0.05307741, -0.05288035, -0.05387415, 
    -0.05344629, -0.05432842, -0.05789149, -0.05682287, -0.06006417, 
    -0.06209305, -0.06347543, -0.06447324, -0.06433131, -0.06406151, 
    -0.06269147, -0.06142794, -0.06048064, -0.05985441, -0.05924317, 
    -0.05742705, -0.0564868, -0.05443173, -0.05479764, -0.05417917, 
    -0.05359444, -0.05262539, -0.05278381, -0.05236075, -0.0541955, 
    -0.05296971, -0.05500703, -0.05444284, -0.05907742, -0.06093621, 
    -0.06174179, -0.06245533, -0.06422237, -0.06299725, -0.06347762, 
    -0.06234037, -0.06162736, -0.06197909, -0.05983737, -0.06066184, 
    -0.05643151, -0.0582196, -0.05366234, -0.05472236, -0.05341107, 
    -0.05407662, -0.05294074, -0.05396203, -0.05220413, -0.05182824, 
    -0.05208483, -0.05110556, -0.05401915, -0.05288283, -0.06198895, 
    -0.06193144, -0.06166426, -0.06284662, -0.06291965, -0.06402266, 
    -0.0630404, -0.06262626, -0.0615863, -0.0609785, -0.06040584, 
    -0.05916393, -0.05780436, -0.055951, -0.05465307, -0.0537984, 
    -0.05432106, -0.05385938, -0.0543757, -0.05461926, -0.05196876, 
    -0.05344229, -0.05124538, -0.05136479, -0.05235071, -0.05135132, 
    -0.06189111, -0.06222245, -0.06338531, -0.0624736, -0.06414384, 
    -0.06320389, -0.0626691, -0.06064438, -0.06020774, -0.05980524, 
    -0.05901763, -0.0580206, -0.05630849, -0.05485638, -0.05356061, 
    -0.05365461, -0.0536215, -0.05333551, -0.0540464, -0.05321962, 
    -0.05308194, -0.05344253, -0.05138079, -0.05196235, -0.05136733, 
    -0.05174523, -0.06211459, -0.06155888, -0.06185858, -0.06129606, 
    -0.06169183, -0.05994954, -0.05943597, -0.05708583, -0.05804005, 
    -0.05652829, -0.05788487, -0.05764232, -0.05647935, -0.05781085, 
    -0.05493544, -0.05687008, -0.05332442, -0.05520468, -0.05320854, 
    -0.05356616, -0.05297528, -0.05245105, -0.05179831, -0.05061301, 
    -0.0508853, -0.04990829, -0.0607389, -0.0600335, -0.06009541, 
    -0.05936459, -0.0588293, -0.05768428, -0.05588993, -0.05655868, 
    -0.0553366, -0.05509414, -0.05695304, -0.05580498, -0.05956567, 
    -0.05894276, -0.059313, -0.06068292, -0.05640379, -0.05856421, 
    -0.05463184, -0.0557599, -0.05252549, -0.05411201, -0.05103573, 
    -0.04976939, -0.04860402, -0.04727286, -0.05965179, -0.06012749, 
    -0.05927826, -0.0581211, -0.05706616, -0.05569047, -0.05555148, 
    -0.05529768, -0.05464528, -0.05410212, -0.05521756, -0.05396673, 
    -0.05879893, -0.05621977, -0.06030814, -0.05904931, -0.05818879, 
    -0.05856497, -0.0566356, -0.05618933, -0.05440849, -0.05532264, 
    -0.05007919, -0.05234078, -0.04628174, -0.0479077, -0.06029448, 
    -0.05965347, -0.05747045, -0.05849991, -0.05559977, -0.0549062, 
    -0.05434826, -0.05364237, -0.05356673, -0.05315297, -0.0538325, 
    -0.0531797, -0.05568757, -0.0545539, -0.05771637, -0.05693161, 
    -0.05729145, -0.05768846, -0.05647115, -0.05519981, -0.0551731, 
    -0.05477112, -0.05365236, -0.05558829, -0.04979353, -0.05330348, 
    -0.05896156, -0.05775695, -0.05758694, -0.05804961, -0.05497537, 
    -0.05607173, -0.05316304, -0.05393538, -0.05267522, -0.05329802, 
    -0.05339021, -0.05420121, -0.05471171, -0.056021, -0.05710727, 
    -0.05798232, -0.05777778, -0.0568203, -0.05512293, -0.05355981, 
    -0.05389871, -0.05277004, -0.05580557, -0.05451385, -0.0550098, 
    -0.05372518, -0.05657651, -0.05413953, -0.05721514, -0.05693931, 
    -0.0560937, -0.05442712, -0.05406478, -0.05368001, -0.05391718, 
    -0.05508048, -0.05527329, -0.05611416, -0.05634827, -0.05699927, 
    -0.05754332, -0.05704601, -0.05652793, -0.05508005, -0.05380409, 
    -0.0524436, -0.0521155, -0.05057382, -0.05182542, -0.04977455, 
    -0.05151306, -0.04853751, -0.05400151, -0.05156532, -0.05605555, 
    -0.05555535, -0.05466075, -0.05265841, -0.05373115, -0.0524786, 
    -0.05528087, -0.05678744, -0.05718347, -0.05792874, -0.05716654, 
    -0.0572282, -0.05650668, -0.05673765, -0.05503256, -0.05594259, 
    -0.05339248, -0.05248842, -0.05000983, -0.04854309, -0.04709026, 
    -0.04646135, -0.04627145, -0.04619226,
  -0.04034989, -0.03907157, -0.03931751, -0.03830527, -0.0388642, 
    -0.03820515, -0.04008809, -0.03902146, -0.03969972, -0.04023352, 
    -0.03640055, -0.03826062, -0.03454635, -0.03567582, -0.032893, 
    -0.03472014, -0.03253405, -0.03294473, -0.03172122, -0.032068, 
    -0.03054241, -0.03156218, -0.02977462, -0.0307836, -0.03062397, 
    -0.03159625, -0.03788041, -0.03662804, -0.03795565, -0.0377747, 
    -0.03785584, -0.03885255, -0.0393627, -0.04044905, -0.04025007, 
    -0.03945309, -0.03769357, -0.03828369, -0.03681071, -0.03684347, 
    -0.03525623, -0.03596495, -0.03337959, -0.03409883, -0.03205347, 
    -0.03255841, -0.03207703, -0.03222241, -0.03207513, -0.03281824, 
    -0.0324982, -0.03315822, -0.03583134, -0.03502848, -0.03746649, 
    -0.0389966, -0.04004079, -0.04079528, -0.04068792, -0.04048387, 
    -0.03944846, -0.03849467, -0.03778033, -0.03730846, -0.03684818, 
    -0.03548229, -0.03477619, -0.03323557, -0.03350961, -0.0330465, 
    -0.03260899, -0.03188465, -0.032003, -0.031687, -0.03305873, -0.03214191, 
    -0.03366648, -0.03324389, -0.03672341, -0.03812378, -0.03873148, 
    -0.03927013, -0.04060553, -0.03967945, -0.04004245, -0.03918332, 
    -0.03864513, -0.03891058, -0.03729562, -0.03791692, -0.03473469, 
    -0.03607803, -0.03265978, -0.03345322, -0.03247185, -0.03296974, 
    -0.03212027, -0.032884, -0.03157006, -0.0312895, -0.031481, -0.03075052, 
    -0.03292674, -0.03207699, -0.03891801, -0.03887461, -0.03867298, 
    -0.03956565, -0.03962082, -0.0404545, -0.03971205, -0.03939921, 
    -0.03861415, -0.03815567, -0.03772395, -0.03678852, -0.03576584, 
    -0.03437416, -0.03340133, -0.03276156, -0.03315272, -0.03280719, 
    -0.03319362, -0.033376, -0.03139437, -0.0324952, -0.03085475, 
    -0.03094379, -0.0316795, -0.03093375, -0.03884417, -0.03909429, 
    -0.03997268, -0.03928392, -0.04054614, -0.03983558, -0.03943156, 
    -0.03790376, -0.03757466, -0.03727143, -0.03667841, -0.0359284, 
    -0.03464237, -0.03355361, -0.03258369, -0.032654, -0.03262923, 
    -0.03241536, -0.03294713, -0.03232871, -0.03222579, -0.03249538, 
    -0.03095573, -0.03138958, -0.03094568, -0.03122756, -0.03901286, 
    -0.03859346, -0.03881962, -0.03839519, -0.03869378, -0.03738012, 
    -0.03699333, -0.03522596, -0.03594302, -0.03480733, -0.03582636, 
    -0.03564405, -0.0347706, -0.03577072, -0.03361284, -0.03506393, 
    -0.03240706, -0.03381459, -0.03232043, -0.03258784, -0.03214608, 
    -0.03175443, -0.03126716, -0.03038348, -0.03058635, -0.02985881, 
    -0.03797501, -0.03744338, -0.03749002, -0.03693959, -0.03653668, 
    -0.03567558, -0.03432836, -0.03483014, -0.03391346, -0.03373175, 
    -0.03512623, -0.03426464, -0.03709099, -0.03662206, -0.03690074, 
    -0.03793281, -0.03471389, -0.03633723, -0.03338542, -0.03423082, 
    -0.03181003, -0.03299623, -0.03069847, -0.02975546, -0.02888924, 
    -0.02790177, -0.03715585, -0.03751419, -0.03687459, -0.03600397, 
    -0.03521119, -0.03417876, -0.03407455, -0.03388429, -0.03339549, 
    -0.03298883, -0.03382424, -0.03288751, -0.03651382, -0.0345758, 
    -0.03765032, -0.03670225, -0.03605486, -0.0363378, -0.03488788, 
    -0.03455296, -0.03321818, -0.033903, -0.02998599, -0.03167209, 
    -0.02716798, -0.02837243, -0.03764003, -0.03715712, -0.03551489, 
    -0.03628886, -0.03411075, -0.03359093, -0.03317308, -0.03264484, 
    -0.03258827, -0.03227889, -0.03278708, -0.03229887, -0.03417659, 
    -0.03332706, -0.0356997, -0.03511014, -0.03538041, -0.03567873, 
    -0.03476444, -0.03381094, -0.03379092, -0.03348975, -0.03265231, 
    -0.03410215, -0.02977343, -0.03239141, -0.0366362, -0.03573021, 
    -0.03560244, -0.03595021, -0.03364275, -0.03446473, -0.03228642, 
    -0.03286405, -0.03192187, -0.03238733, -0.03245626, -0.033063, 
    -0.03344524, -0.03442667, -0.03524206, -0.03589962, -0.03574586, 
    -0.03502655, -0.03375332, -0.03258309, -0.03283662, -0.03199272, 
    -0.03426508, -0.03329707, -0.03366855, -0.03270678, -0.03484353, 
    -0.03301683, -0.03532309, -0.03511592, -0.03448121, -0.03323212, 
    -0.03296089, -0.032673, -0.03285043, -0.03372151, -0.03386601, 
    -0.03449655, -0.03467222, -0.03516095, -0.03556966, -0.03519605, 
    -0.03480706, -0.03372119, -0.03276582, -0.03174886, -0.03150389, 
    -0.03035429, -0.03128739, -0.0297593, -0.03105436, -0.02883985, 
    -0.03291354, -0.03109335, -0.03445259, -0.03407745, -0.03340707, 
    -0.03190931, -0.03271126, -0.03177501, -0.03387169, -0.03500188, 
    -0.0352993, -0.03585934, -0.03528658, -0.03533289, -0.03479112, 
    -0.03496449, -0.03368561, -0.03436785, -0.03245796, -0.03178234, 
    -0.02993437, -0.028844, -0.02776648, -0.02730087, -0.02716037, -0.0271018,
  -0.01970494, -0.0187005, -0.01889312, -0.01810233, -0.01853833, -0.0180244, 
    -0.01949858, -0.01866129, -0.01919306, -0.01961317, -0.0166292, 
    -0.01806757, -0.01521542, -0.01607412, -0.01397334, -0.01534703, 
    -0.01370616, -0.01401192, -0.01310461, -0.01336065, -0.01224113, 
    -0.01298748, -0.01168475, -0.01241691, -0.01230052, -0.01301256, 
    -0.01777201, -0.01680408, -0.01783044, -0.01768998, -0.01775294, 
    -0.01852922, -0.01892854, -0.0197832, -0.01962622, -0.01899943, 
    -0.01762706, -0.01808553, -0.01694472, -0.01696995, -0.0157542, 
    -0.01629521, -0.01433697, -0.01487742, -0.0133499, -0.01372426, 
    -0.01336733, -0.01347495, -0.01336593, -0.01391762, -0.01367953, 
    -0.01417134, -0.01619298, -0.015581, -0.01745114, -0.01864185, 
    -0.01946134, -0.02005677, -0.01997188, -0.01981068, -0.0189958, 
    -0.01824989, -0.01769435, -0.01732888, -0.01697358, -0.01592643, 
    -0.01538951, -0.01422917, -0.01443441, -0.01408787, -0.01376186, 
    -0.01322516, -0.01331259, -0.01307939, -0.014097, -0.01341534, 
    -0.01455212, -0.0142354, -0.01687748, -0.01796111, -0.01843465, 
    -0.01885598, -0.01990677, -0.01917714, -0.01946264, -0.01878798, 
    -0.01836725, -0.01857458, -0.01731896, -0.01780036, -0.01535805, 
    -0.0163818, -0.01379964, -0.01439214, -0.01365996, -0.01403058, 
    -0.01339932, -0.01396663, -0.01299328, -0.01278711, -0.01292777, 
    -0.01239277, -0.0139985, -0.0133673, -0.01858039, -0.01854647, 
    -0.01838898, -0.01908777, -0.01913109, -0.01978749, -0.01920275, 
    -0.01895717, -0.01834307, -0.01798592, -0.01765062, -0.01692762, 
    -0.0161429, -0.01508521, -0.01435325, -0.0138754, -0.01416722, 
    -0.01390938, -0.0141978, -0.01433428, -0.0128641, -0.0136773, 
    -0.01246885, -0.01253391, -0.01307386, -0.01252657, -0.01852267, 
    -0.01871828, -0.01940771, -0.0188668, -0.01985985, -0.01929986, 
    -0.01898255, -0.01779014, -0.01753491, -0.01730025, -0.01684284, 
    -0.01626723, -0.01528811, -0.01446741, -0.01374306, -0.01379534, 
    -0.01377692, -0.01361802, -0.01401371, -0.01355374, -0.01347746, 
    -0.01367743, -0.01254264, -0.01286058, -0.0125353, -0.01274168, 
    -0.01865456, -0.01832693, -0.0185035, -0.01817236, -0.01840522, 
    -0.01738431, -0.0170855, -0.01573116, -0.01627842, -0.01541313, 
    -0.01618917, -0.01604987, -0.01538528, -0.01614663, -0.01451186, 
    -0.01560794, -0.01361186, -0.01466342, -0.0135476, -0.01374614, 
    -0.01341843, -0.01312909, -0.01277072, -0.01212556, -0.01227312, 
    -0.01174551, -0.01784548, -0.01743325, -0.01746936, -0.01704405, 
    -0.01673382, -0.01607395, -0.01505061, -0.01543043, -0.0147378, 
    -0.01460115, -0.0156553, -0.01500249, -0.01716087, -0.01679948, 
    -0.0170141, -0.0178127, -0.01534229, -0.01658059, -0.01434134, 
    -0.01497698, -0.01317009, -0.01405035, -0.01235481, -0.01167093, 
    -0.01104941, -0.0103492, -0.01721095, -0.01748807, -0.01699394, 
    -0.01632507, -0.01571992, -0.01493769, -0.01485912, -0.01471585, 
    -0.01434888, -0.01404482, -0.01467067, -0.01396925, -0.01671625, 
    -0.01523771, -0.01759353, -0.01686119, -0.01636405, -0.01658102, 
    -0.01547424, -0.01522042, -0.01421616, -0.01472992, -0.01183743, 
    -0.0130684, -0.009834951, -0.0106818, -0.01758556, -0.01721193, 
    -0.0159513, -0.01654346, -0.01488641, -0.01449541, -0.01418244, 
    -0.01378853, -0.01374646, -0.0135168, -0.0138944, -0.01353161, 
    -0.01493606, -0.01429763, -0.01609237, -0.01564306, -0.01584877, 
    -0.01607634, -0.01538061, -0.01466067, -0.01464562, -0.01441951, 
    -0.01379409, -0.01487992, -0.01168388, -0.01360025, -0.01681036, 
    -0.01611567, -0.01601809, -0.01628392, -0.01453431, -0.01515368, 
    -0.01352238, -0.01395176, -0.01325265, -0.01359722, -0.01364838, 
    -0.01410019, -0.01438616, -0.0151249, -0.01574341, -0.0162452, 
    -0.01612764, -0.01557953, -0.01461736, -0.01374261, -0.01393131, 
    -0.01330499, -0.01500283, -0.01427518, -0.01455368, -0.01383462, 
    -0.01544058, -0.01406572, -0.0158051, -0.01564745, -0.01516614, 
    -0.01422659, -0.01402397, -0.01380948, -0.01394161, -0.01459346, 
    -0.01470209, -0.01517775, -0.01531072, -0.0156817, -0.01599308, 
    -0.0157084, -0.01541292, -0.01459322, -0.01387857, -0.01312498, 
    -0.0129446, -0.01210436, -0.01278557, -0.0116737, -0.0126148, 
    -0.01101418, -0.01398866, -0.01264334, -0.01514449, -0.01486131, 
    -0.01435756, -0.01324337, -0.01383795, -0.01314426, -0.01470637, 
    -0.01556079, -0.01578699, -0.01621439, -0.0157773, -0.01581257, 
    -0.01540083, -0.0155324, -0.01456649, -0.01508045, -0.01364964, 
    -0.01314967, -0.0118001, -0.01101713, -0.01025399, -0.009927679, 
    -0.009829645, -0.009788835,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  363.1486, 364.9598, 364.6072, 366.0715, 365.2586, 366.2182, 363.5153, 
    365.032, 364.0632, 363.3113, 368.9243, 366.1369, 371.821, 370.0447, 
    374.5131, 371.5448, 375.1133, 374.4269, 376.4946, 375.9015, 378.5548, 
    376.7685, 379.9343, 378.1275, 378.4099, 376.7097, 366.6964, 368.5766, 
    366.5853, 366.853, 366.7328, 365.2755, 364.5428, 363.0099, 363.2882, 
    364.4138, 366.9734, 366.103, 368.2985, 368.2488, 370.7001, 369.5951, 
    373.7084, 372.538, 375.9262, 375.0723, 375.8861, 375.6392, 375.8893, 
    374.6375, 375.1735, 374.0731, 369.8025, 371.0575, 367.3115, 365.0679, 
    363.5818, 362.5281, 362.6771, 362.9613, 364.4203, 365.7948, 366.8445, 
    367.5479, 368.2416, 370.3477, 371.4559, 373.9455, 373.4951, 374.2581, 
    374.9874, 376.2144, 376.0122, 376.5535, 374.2377, 375.7758, 373.2388, 
    373.9317, 368.4315, 366.3376, 365.4509, 364.675, 362.7917, 364.092, 
    363.5795, 364.7993, 365.5759, 365.1917, 367.5671, 366.6425, 371.5217, 
    369.4203, 374.9023, 373.5875, 375.2178, 374.3853, 375.8126, 374.5279, 
    376.7549, 377.2411, 376.9089, 378.1859, 374.4568, 375.8862, 365.1809, 
    365.2436, 365.5355, 364.2535, 364.1752, 363.0023, 364.0457, 364.4906, 
    365.6209, 366.2907, 366.9282, 368.3322, 369.9044, 372.0959, 373.6727, 
    374.732, 374.0821, 374.6559, 374.0146, 373.7142, 377.059, 375.1786, 
    378.002, 377.8454, 376.5664, 377.863, 365.2876, 364.9271, 363.6776, 
    364.6552, 362.8744, 363.871, 364.4445, 366.662, 367.1501, 367.6034, 
    368.4995, 369.6518, 371.6681, 373.4232, 375.0298, 374.9119, 374.9534, 
    375.313, 374.4229, 375.4593, 375.6335, 375.1783, 377.8244, 377.0672, 
    377.8421, 377.3489, 365.0442, 365.651, 365.3231, 365.9399, 365.5054, 
    367.4407, 368.0222, 370.7477, 369.6292, 371.4066, 369.8102, 370.0943, 
    371.4649, 369.8968, 373.3265, 371.0019, 375.327, 372.9981, 375.4733, 
    375.0229, 375.7687, 376.4376, 377.2799, 378.8377, 378.4766, 379.7815, 
    366.5567, 367.346, 367.2763, 368.1033, 368.7157, 370.045, 372.1692, 
    371.3704, 372.8375, 373.1325, 370.9038, 372.2714, 367.8748, 368.5855, 
    368.1621, 366.619, 371.5546, 369.0212, 373.6988, 372.3256, 376.3422, 
    374.3415, 378.2779, 379.9693, 381.5645, 383.4352, 367.7771, 367.2402, 
    368.2016, 369.5348, 370.7707, 372.4093, 372.5771, 372.8848, 373.6822, 
    374.3536, 372.9823, 374.522, 368.7509, 371.774, 367.0376, 368.4634, 
    369.4561, 369.0202, 371.2791, 371.8103, 373.9742, 372.8544, 379.5516, 
    376.5793, 384.8626, 382.5365, 367.0528, 367.7751, 370.2964, 369.0954, 
    372.5188, 373.3622, 374.0485, 374.9274, 375.0222, 375.5436, 374.6894, 
    375.5097, 372.4128, 373.7947, 370.0074, 370.9291, 370.5061, 370.0401, 
    371.4743, 373.0039, 373.0363, 373.5277, 374.9153, 372.5326, 379.937, 
    375.3539, 368.5638, 369.96, 370.1593, 369.618, 373.2776, 371.951, 
    375.5308, 374.5611, 376.1507, 375.3603, 375.2441, 374.2306, 373.6006, 
    372.0119, 370.7223, 369.6964, 369.9355, 371.0605, 373.0975, 375.0309, 
    374.6069, 376.0297, 372.2706, 373.8441, 373.2356, 374.8236, 371.3492, 
    374.3076, 370.5956, 370.92, 371.9247, 373.9512, 374.4, 374.8802, 
    374.5838, 373.1493, 372.9145, 371.9002, 371.6207, 370.8493, 370.2105, 
    370.7943, 371.4069, 373.1497, 374.725, 376.4471, 376.8692, 378.8901, 
    377.245, 379.9626, 377.652, 381.6571, 374.479, 377.5835, 371.9704, 
    372.5724, 373.6633, 376.1724, 374.8161, 376.4024, 372.9052, 371.0995, 
    370.6328, 369.7589, 370.6526, 370.5803, 371.4321, 371.1582, 373.2077, 
    372.1059, 375.2413, 376.3897, 379.6447, 381.6491, 383.6957, 384.6016, 
    384.8776, 384.993 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.194319e-08, 6.221824e-08, 6.216477e-08, 6.238663e-08, 6.226357e-08, 
    6.240884e-08, 6.199895e-08, 6.222916e-08, 6.20822e-08, 6.196796e-08, 
    6.281724e-08, 6.239654e-08, 6.325438e-08, 6.2986e-08, 6.366027e-08, 
    6.321261e-08, 6.375054e-08, 6.364737e-08, 6.395796e-08, 6.386897e-08, 
    6.426626e-08, 6.399903e-08, 6.447225e-08, 6.420245e-08, 6.424465e-08, 
    6.399021e-08, 6.248121e-08, 6.276485e-08, 6.24644e-08, 6.250485e-08, 
    6.24867e-08, 6.22661e-08, 6.215493e-08, 6.192218e-08, 6.196444e-08, 
    6.213539e-08, 6.252303e-08, 6.239145e-08, 6.272312e-08, 6.271563e-08, 
    6.308491e-08, 6.29184e-08, 6.35392e-08, 6.336274e-08, 6.387269e-08, 
    6.374443e-08, 6.386666e-08, 6.38296e-08, 6.386715e-08, 6.367905e-08, 
    6.375964e-08, 6.359412e-08, 6.294958e-08, 6.313898e-08, 6.257413e-08, 
    6.223455e-08, 6.200905e-08, 6.184904e-08, 6.187166e-08, 6.191478e-08, 
    6.213639e-08, 6.234479e-08, 6.250362e-08, 6.260986e-08, 6.271455e-08, 
    6.303143e-08, 6.31992e-08, 6.357487e-08, 6.350708e-08, 6.362193e-08, 
    6.373168e-08, 6.391591e-08, 6.388559e-08, 6.396677e-08, 6.361891e-08, 
    6.385008e-08, 6.346847e-08, 6.357283e-08, 6.274296e-08, 6.242695e-08, 
    6.22926e-08, 6.217505e-08, 6.188905e-08, 6.208655e-08, 6.200869e-08, 
    6.219393e-08, 6.231164e-08, 6.225343e-08, 6.261276e-08, 6.247306e-08, 
    6.320914e-08, 6.289206e-08, 6.371887e-08, 6.352099e-08, 6.37663e-08, 
    6.364113e-08, 6.385561e-08, 6.366258e-08, 6.399698e-08, 6.406979e-08, 
    6.402004e-08, 6.421121e-08, 6.365187e-08, 6.386666e-08, 6.225179e-08, 
    6.226129e-08, 6.230552e-08, 6.211108e-08, 6.209918e-08, 6.192101e-08, 
    6.207955e-08, 6.214706e-08, 6.231847e-08, 6.241986e-08, 6.251624e-08, 
    6.272818e-08, 6.296489e-08, 6.329594e-08, 6.353382e-08, 6.369329e-08, 
    6.359551e-08, 6.368183e-08, 6.358533e-08, 6.35401e-08, 6.404251e-08, 
    6.376038e-08, 6.418371e-08, 6.416029e-08, 6.39687e-08, 6.416293e-08, 
    6.226796e-08, 6.221332e-08, 6.202362e-08, 6.217208e-08, 6.190162e-08, 
    6.2053e-08, 6.214005e-08, 6.247596e-08, 6.254979e-08, 6.261823e-08, 
    6.275342e-08, 6.292692e-08, 6.323132e-08, 6.349621e-08, 6.373806e-08, 
    6.372034e-08, 6.372658e-08, 6.37806e-08, 6.364677e-08, 6.380257e-08, 
    6.382872e-08, 6.376035e-08, 6.415715e-08, 6.404378e-08, 6.415979e-08, 
    6.408597e-08, 6.223108e-08, 6.232302e-08, 6.227334e-08, 6.236676e-08, 
    6.230094e-08, 6.259361e-08, 6.268137e-08, 6.309205e-08, 6.29235e-08, 
    6.319176e-08, 6.295076e-08, 6.299346e-08, 6.32005e-08, 6.296379e-08, 
    6.348159e-08, 6.313051e-08, 6.37827e-08, 6.343204e-08, 6.380468e-08, 
    6.373701e-08, 6.384905e-08, 6.394939e-08, 6.407564e-08, 6.430859e-08, 
    6.425465e-08, 6.444949e-08, 6.246009e-08, 6.257934e-08, 6.256885e-08, 
    6.269367e-08, 6.278598e-08, 6.298608e-08, 6.330703e-08, 6.318634e-08, 
    6.340794e-08, 6.345242e-08, 6.311577e-08, 6.332245e-08, 6.265917e-08, 
    6.276631e-08, 6.270252e-08, 6.24695e-08, 6.321414e-08, 6.283195e-08, 
    6.353775e-08, 6.333067e-08, 6.393508e-08, 6.363447e-08, 6.422496e-08, 
    6.44774e-08, 6.471507e-08, 6.499279e-08, 6.264444e-08, 6.256341e-08, 
    6.270852e-08, 6.290927e-08, 6.309559e-08, 6.334329e-08, 6.336865e-08, 
    6.341506e-08, 6.353527e-08, 6.363636e-08, 6.342972e-08, 6.366169e-08, 
    6.279114e-08, 6.324732e-08, 6.253276e-08, 6.274789e-08, 6.289744e-08, 
    6.283185e-08, 6.317255e-08, 6.325285e-08, 6.35792e-08, 6.34105e-08, 
    6.441508e-08, 6.397057e-08, 6.52043e-08, 6.485946e-08, 6.253509e-08, 
    6.264417e-08, 6.302381e-08, 6.284317e-08, 6.335984e-08, 6.348703e-08, 
    6.359044e-08, 6.372262e-08, 6.37369e-08, 6.381522e-08, 6.368688e-08, 
    6.381016e-08, 6.334383e-08, 6.355221e-08, 6.298043e-08, 6.311958e-08, 
    6.305557e-08, 6.298534e-08, 6.320207e-08, 6.343297e-08, 6.343792e-08, 
    6.351196e-08, 6.372059e-08, 6.336194e-08, 6.447243e-08, 6.378654e-08, 
    6.276311e-08, 6.297321e-08, 6.300324e-08, 6.292185e-08, 6.347427e-08, 
    6.32741e-08, 6.381332e-08, 6.366758e-08, 6.390638e-08, 6.378771e-08, 
    6.377025e-08, 6.361785e-08, 6.352296e-08, 6.328327e-08, 6.308827e-08, 
    6.293366e-08, 6.296961e-08, 6.313945e-08, 6.34471e-08, 6.373818e-08, 
    6.367442e-08, 6.388823e-08, 6.332237e-08, 6.355963e-08, 6.346792e-08, 
    6.370704e-08, 6.318313e-08, 6.362922e-08, 6.306912e-08, 6.311822e-08, 
    6.327013e-08, 6.35757e-08, 6.364334e-08, 6.371553e-08, 6.367099e-08, 
    6.345491e-08, 6.341952e-08, 6.326643e-08, 6.322416e-08, 6.310753e-08, 
    6.301097e-08, 6.309919e-08, 6.319184e-08, 6.3455e-08, 6.369219e-08, 
    6.395081e-08, 6.401412e-08, 6.43163e-08, 6.407029e-08, 6.447625e-08, 
    6.413108e-08, 6.472865e-08, 6.36551e-08, 6.412095e-08, 6.327704e-08, 
    6.336795e-08, 6.353237e-08, 6.390953e-08, 6.370593e-08, 6.394406e-08, 
    6.341813e-08, 6.314531e-08, 6.307474e-08, 6.294306e-08, 6.307775e-08, 
    6.306679e-08, 6.319569e-08, 6.315427e-08, 6.346375e-08, 6.329751e-08, 
    6.376981e-08, 6.394218e-08, 6.442907e-08, 6.472758e-08, 6.503151e-08, 
    6.51657e-08, 6.520654e-08, 6.522362e-08 ;

 SOM_C_LEACHED =
  -1.182477e-20, -2.601569e-20, -2.34767e-20, -1.301268e-20, -2.518354e-21, 
    3.460844e-20, 1.612764e-20, 2.733447e-20, -1.638961e-20, 5.825766e-20, 
    1.490369e-20, -7.576481e-20, 6.217534e-20, 1.590697e-20, -2.361731e-20, 
    -6.248373e-21, 2.145471e-21, -5.304007e-20, 7.33436e-20, -2.327935e-21, 
    3.838925e-20, 3.178481e-20, 3.05175e-20, 5.769225e-20, -4.408063e-20, 
    -5.349289e-20, -6.290416e-20, 2.993178e-20, -3.71387e-20, 3.736754e-20, 
    1.017639e-20, 2.442018e-20, -3.481807e-20, -1.441853e-20, 9.422452e-23, 
    8.412555e-21, -5.94291e-20, -4.028371e-20, -4.234712e-22, 4.70995e-20, 
    -9.336059e-21, -1.444764e-20, -2.620468e-20, -5.500884e-20, -1.93967e-21, 
    -9.794889e-20, 7.481811e-21, -9.527274e-22, -7.067712e-21, 1.250601e-20, 
    1.917698e-20, -5.047199e-21, -3.459571e-20, 4.499851e-20, 5.281374e-20, 
    -2.759899e-20, -2.527514e-20, -5.273082e-20, 4.967155e-20, -2.830899e-20, 
    7.983581e-21, 9.287923e-20, -2.821194e-20, 3.606604e-20, 8.209621e-21, 
    4.295256e-20, 7.78027e-20, -2.831766e-20, -2.303145e-20, 5.721339e-21, 
    4.488034e-20, -4.826403e-21, -1.981922e-20, 1.32163e-20, -5.69521e-20, 
    -4.42445e-20, 3.474999e-20, 5.246696e-20, -4.471545e-21, 5.29968e-20, 
    -7.989225e-20, 2.339459e-20, 4.73709e-20, -1.856438e-20, -2.053759e-20, 
    1.291882e-20, -2.981316e-20, -3.08288e-20, 1.424514e-20, 2.678039e-20, 
    3.674746e-20, 5.607903e-20, -3.315467e-20, -7.672601e-20, 1.501834e-20, 
    1.395772e-20, -3.645009e-20, -4.790584e-20, 9.400588e-22, -1.426464e-20, 
    -5.126996e-21, -1.098602e-20, 1.570229e-20, 3.072212e-20, 3.917131e-20, 
    -2.425872e-20, 3.176556e-20, 3.431031e-20, -7.722487e-21, -1.060202e-20, 
    -2.330226e-20, -8.12595e-22, -3.090773e-20, 3.496715e-20, 3.548903e-20, 
    -1.846493e-20, 3.443839e-20, 4.866262e-20, -2.256752e-20, -3.48545e-21, 
    -6.618413e-20, 8.745269e-21, 3.874891e-20, 2.661325e-20, -1.1408e-20, 
    -2.62441e-20, -3.862331e-20, 8.335346e-20, -2.211887e-20, 3.953664e-20, 
    -1.622592e-20, 2.995216e-20, -1.890575e-20, -3.113574e-20, -9.344069e-21, 
    1.975482e-20, 3.218198e-20, 5.226935e-20, 8.085881e-21, -1.419353e-20, 
    6.614572e-21, 2.374299e-20, -1.361332e-20, -6.138354e-20, 9.349928e-20, 
    -2.139534e-20, 1.89192e-20, 3.963535e-20, -4.756321e-20, 7.083776e-20, 
    -2.21932e-20, -4.575047e-20, 1.047875e-20, 1.745944e-20, 1.596916e-20, 
    7.289521e-21, 5.687401e-20, 1.544226e-20, -3.249265e-20, -2.105412e-20, 
    4.729689e-20, 1.857252e-20, -7.217404e-20, 2.965507e-20, 4.603403e-20, 
    2.010353e-20, 1.450983e-20, 4.284534e-21, -1.568953e-20, -1.504156e-20, 
    1.270362e-20, -5.183202e-20, -6.866857e-20, -2.255369e-20, -1.322811e-20, 
    -2.420561e-20, -3.275507e-20, 3.792195e-20, 5.851602e-21, -3.643251e-20, 
    -8.522016e-21, -4.602616e-20, 5.509006e-20, 4.994056e-21, 3.474385e-20, 
    3.291892e-20, 2.005698e-20, -5.978786e-20, 1.238229e-20, -6.400008e-20, 
    1.922117e-21, -1.600738e-20, 3.438089e-20, -3.281182e-20, 4.28251e-20, 
    1.835345e-20, 1.039286e-19, 4.38728e-20, 1.31405e-20, 4.85855e-21, 
    -6.124373e-20, -3.782094e-20, 6.803328e-20, -7.17496e-20, 6.802254e-20, 
    -9.578936e-20, 4.326812e-20, 3.923172e-20, 1.396667e-20, 2.449321e-21, 
    5.014785e-21, -1.421239e-21, 3.261186e-20, -2.832808e-20, 2.273815e-20, 
    -4.871813e-20, -1.948595e-20, 4.135405e-21, 1.108571e-20, -4.726103e-20, 
    5.914714e-22, 1.819105e-20, 1.493503e-20, -2.938236e-20, -1.753115e-20, 
    2.028979e-20, 2.575939e-20, -7.077639e-20, 5.783837e-20, 5.337188e-20, 
    4.872807e-20, 2.818125e-20, -6.532411e-20, 4.346962e-20, -6.398523e-22, 
    1.329829e-20, 2.037737e-20, 2.927852e-20, 1.208457e-20, 2.51156e-20, 
    -3.028562e-20, -3.496377e-20, 4.191848e-20, 6.716296e-21, -3.763447e-20, 
    1.044191e-20, -4.258199e-20, -4.519518e-20, 5.075281e-20, 3.538285e-20, 
    -4.115156e-20, 1.884755e-20, -3.236108e-20, -7.541673e-20, 9.983011e-21, 
    -1.662834e-20, 9.979438e-21, -1.920103e-20, 3.041375e-20, 2.598769e-20, 
    -5.473106e-20, 6.863032e-20, -1.661637e-20, 6.644165e-21, -5.438327e-21, 
    -5.823017e-20, -1.907265e-20, 2.06156e-20, -8.471532e-20, 9.478473e-21, 
    3.459108e-20, 3.37488e-20, -6.707497e-20, -2.125255e-21, -2.090387e-20, 
    -8.948279e-22, -4.813302e-20, 3.070399e-20, 7.800716e-20, -3.371756e-20, 
    2.026862e-20, 4.375029e-20, -2.627965e-20, 1.607427e-20, -1.318952e-20, 
    6.366713e-20, -1.876828e-20, 1.986714e-20, -1.190291e-20, -1.020442e-20, 
    -4.188722e-21, 5.419983e-21, -4.736524e-20, -2.97326e-20, -1.636561e-20, 
    -3.984328e-20, -6.559126e-21, -8.737105e-22, 4.92214e-20, -7.263649e-21, 
    2.088488e-20, 2.109619e-20, -4.973516e-21, -5.441853e-20, 2.924216e-20, 
    -4.49288e-21, -3.982829e-21, -6.376841e-20, 3.353464e-20, 2.542208e-20, 
    -1.456299e-20, -4.546707e-21, 1.893524e-20, 6.70968e-20, 5.223148e-20, 
    1.09807e-20, 1.900437e-20, -5.602667e-20, 2.789057e-20, 4.279362e-20, 
    1.122005e-20, -2.303763e-20, 3.611915e-20, 3.570133e-20, -4.533734e-21, 
    -2.241725e-20, -5.639212e-20, 3.112817e-20, 9.418056e-21, -1.95021e-20, 
    -4.756255e-20, 1.957267e-20, 5.742362e-20, -1.150679e-19, -4.631152e-20, 
    3.693092e-20, -2.974299e-20, 1.794585e-21 ;

 SR =
  6.194416e-08, 6.221921e-08, 6.216575e-08, 6.238761e-08, 6.226454e-08, 
    6.240981e-08, 6.199993e-08, 6.223013e-08, 6.208317e-08, 6.196893e-08, 
    6.281821e-08, 6.239751e-08, 6.325536e-08, 6.298698e-08, 6.366125e-08, 
    6.321359e-08, 6.375153e-08, 6.364835e-08, 6.395895e-08, 6.386996e-08, 
    6.426725e-08, 6.400002e-08, 6.447324e-08, 6.420344e-08, 6.424563e-08, 
    6.39912e-08, 6.248218e-08, 6.276583e-08, 6.246538e-08, 6.250582e-08, 
    6.248767e-08, 6.226708e-08, 6.215591e-08, 6.192315e-08, 6.19654e-08, 
    6.213637e-08, 6.2524e-08, 6.239242e-08, 6.272409e-08, 6.27166e-08, 
    6.308589e-08, 6.291938e-08, 6.354018e-08, 6.336372e-08, 6.387368e-08, 
    6.374542e-08, 6.386765e-08, 6.383059e-08, 6.386814e-08, 6.368003e-08, 
    6.376062e-08, 6.359511e-08, 6.295056e-08, 6.313996e-08, 6.25751e-08, 
    6.223551e-08, 6.201002e-08, 6.185e-08, 6.187263e-08, 6.191575e-08, 
    6.213737e-08, 6.234576e-08, 6.250459e-08, 6.261083e-08, 6.271553e-08, 
    6.303241e-08, 6.320018e-08, 6.357585e-08, 6.350807e-08, 6.362291e-08, 
    6.373266e-08, 6.39169e-08, 6.388658e-08, 6.396775e-08, 6.361989e-08, 
    6.385107e-08, 6.346945e-08, 6.357381e-08, 6.274394e-08, 6.242792e-08, 
    6.229357e-08, 6.217602e-08, 6.189002e-08, 6.208752e-08, 6.200966e-08, 
    6.219491e-08, 6.231262e-08, 6.22544e-08, 6.261374e-08, 6.247403e-08, 
    6.321012e-08, 6.289304e-08, 6.371985e-08, 6.352198e-08, 6.376729e-08, 
    6.364211e-08, 6.38566e-08, 6.366356e-08, 6.399797e-08, 6.407078e-08, 
    6.402102e-08, 6.421219e-08, 6.365286e-08, 6.386765e-08, 6.225277e-08, 
    6.226226e-08, 6.23065e-08, 6.211204e-08, 6.210015e-08, 6.192198e-08, 
    6.208052e-08, 6.214803e-08, 6.231944e-08, 6.242083e-08, 6.251722e-08, 
    6.272915e-08, 6.296587e-08, 6.329692e-08, 6.353481e-08, 6.369427e-08, 
    6.359649e-08, 6.368282e-08, 6.358631e-08, 6.354109e-08, 6.40435e-08, 
    6.376137e-08, 6.41847e-08, 6.416128e-08, 6.396969e-08, 6.416391e-08, 
    6.226892e-08, 6.221429e-08, 6.202459e-08, 6.217304e-08, 6.190258e-08, 
    6.205396e-08, 6.214101e-08, 6.247694e-08, 6.255076e-08, 6.26192e-08, 
    6.27544e-08, 6.29279e-08, 6.32323e-08, 6.349719e-08, 6.373904e-08, 
    6.372132e-08, 6.372756e-08, 6.378159e-08, 6.364776e-08, 6.380356e-08, 
    6.38297e-08, 6.376134e-08, 6.415814e-08, 6.404477e-08, 6.416078e-08, 
    6.408697e-08, 6.223205e-08, 6.232399e-08, 6.227431e-08, 6.236773e-08, 
    6.230191e-08, 6.259458e-08, 6.268234e-08, 6.309303e-08, 6.292449e-08, 
    6.319274e-08, 6.295173e-08, 6.299444e-08, 6.320148e-08, 6.296477e-08, 
    6.348257e-08, 6.313149e-08, 6.378369e-08, 6.343302e-08, 6.380566e-08, 
    6.3738e-08, 6.385004e-08, 6.395038e-08, 6.407663e-08, 6.430958e-08, 
    6.425564e-08, 6.445048e-08, 6.246106e-08, 6.258032e-08, 6.256982e-08, 
    6.269464e-08, 6.278695e-08, 6.298706e-08, 6.330801e-08, 6.318732e-08, 
    6.340892e-08, 6.345341e-08, 6.311675e-08, 6.332343e-08, 6.266014e-08, 
    6.276728e-08, 6.27035e-08, 6.247047e-08, 6.321512e-08, 6.283292e-08, 
    6.353874e-08, 6.333165e-08, 6.393607e-08, 6.363545e-08, 6.422594e-08, 
    6.447839e-08, 6.471606e-08, 6.499378e-08, 6.264541e-08, 6.256438e-08, 
    6.270949e-08, 6.291025e-08, 6.309657e-08, 6.334428e-08, 6.336963e-08, 
    6.341604e-08, 6.353626e-08, 6.363734e-08, 6.34307e-08, 6.366268e-08, 
    6.279212e-08, 6.32483e-08, 6.253374e-08, 6.274887e-08, 6.289842e-08, 
    6.283283e-08, 6.317353e-08, 6.325383e-08, 6.358018e-08, 6.341148e-08, 
    6.441608e-08, 6.397156e-08, 6.52053e-08, 6.486045e-08, 6.253607e-08, 
    6.264514e-08, 6.302479e-08, 6.284415e-08, 6.336082e-08, 6.348802e-08, 
    6.359143e-08, 6.372361e-08, 6.373789e-08, 6.381621e-08, 6.368786e-08, 
    6.381114e-08, 6.334481e-08, 6.355319e-08, 6.298141e-08, 6.312055e-08, 
    6.305654e-08, 6.298632e-08, 6.320305e-08, 6.343395e-08, 6.34389e-08, 
    6.351294e-08, 6.372157e-08, 6.336292e-08, 6.447343e-08, 6.378752e-08, 
    6.276409e-08, 6.297419e-08, 6.300422e-08, 6.292283e-08, 6.347526e-08, 
    6.327508e-08, 6.38143e-08, 6.366856e-08, 6.390736e-08, 6.37887e-08, 
    6.377123e-08, 6.361883e-08, 6.352395e-08, 6.328425e-08, 6.308925e-08, 
    6.293464e-08, 6.297059e-08, 6.314043e-08, 6.344808e-08, 6.373917e-08, 
    6.367541e-08, 6.388921e-08, 6.332336e-08, 6.356061e-08, 6.34689e-08, 
    6.370803e-08, 6.318411e-08, 6.36302e-08, 6.307009e-08, 6.31192e-08, 
    6.327111e-08, 6.357669e-08, 6.364433e-08, 6.371651e-08, 6.367197e-08, 
    6.34559e-08, 6.34205e-08, 6.326741e-08, 6.322514e-08, 6.310851e-08, 
    6.301195e-08, 6.310017e-08, 6.319282e-08, 6.345599e-08, 6.369318e-08, 
    6.39518e-08, 6.401511e-08, 6.431729e-08, 6.407128e-08, 6.447725e-08, 
    6.413207e-08, 6.472964e-08, 6.365608e-08, 6.412193e-08, 6.327802e-08, 
    6.336893e-08, 6.353335e-08, 6.391052e-08, 6.370691e-08, 6.394504e-08, 
    6.341912e-08, 6.314629e-08, 6.307572e-08, 6.294403e-08, 6.307872e-08, 
    6.306777e-08, 6.319667e-08, 6.315525e-08, 6.346473e-08, 6.329849e-08, 
    6.377079e-08, 6.394317e-08, 6.443005e-08, 6.472857e-08, 6.503251e-08, 
    6.51667e-08, 6.520754e-08, 6.522462e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3407592, -0.3407649, -0.3407638, -0.3407683, -0.3407659, -0.3407688, 
    -0.3407604, -0.3407651, -0.3407621, -0.3407598, -0.3407897, -0.3407685, 
    -0.3408154, -0.3407935, -0.3408239, -0.3407981, -0.3408258, -0.3408237, 
    -0.3408302, -0.3408284, -0.3408365, -0.3408311, -0.3408408, -0.3408352, 
    -0.3408361, -0.3408309, -0.3407704, -0.3407886, -0.34077, -0.3407708, 
    -0.3407705, -0.3407659, -0.3407635, -0.3407589, -0.3407597, -0.3407632, 
    -0.3407712, -0.3407685, -0.340788, -0.3407879, -0.3407956, -0.3407921, 
    -0.3408215, -0.3408178, -0.3408284, -0.3408258, -0.3408283, -0.3408276, 
    -0.3408283, -0.3408244, -0.3408261, -0.3408226, -0.3407927, -0.3407967, 
    -0.3407723, -0.3407651, -0.3407606, -0.3407573, -0.3407578, -0.3407587, 
    -0.3407632, -0.3407676, -0.3407709, -0.3407857, -0.3407879, -0.3407943, 
    -0.3407979, -0.3408222, -0.3408208, -0.3408231, -0.3408255, -0.3408293, 
    -0.3408287, -0.3408304, -0.3408231, -0.3408279, -0.34082, -0.3408222, 
    -0.3407881, -0.3407692, -0.3407663, -0.340764, -0.3407581, -0.3407622, 
    -0.3407606, -0.3407645, -0.3407669, -0.3407657, -0.3407857, -0.3407702, 
    -0.3407981, -0.3407915, -0.3408252, -0.3408211, -0.3408262, -0.3408236, 
    -0.3408281, -0.3408241, -0.340831, -0.3408325, -0.3408315, -0.3408355, 
    -0.3408238, -0.3408283, -0.3407657, -0.3407658, -0.3407668, -0.3407627, 
    -0.3407625, -0.3407588, -0.3407621, -0.3407634, -0.3407671, -0.3407691, 
    -0.3407711, -0.3407881, -0.340793, -0.3408163, -0.3408214, -0.3408247, 
    -0.3408227, -0.3408245, -0.3408225, -0.3408215, -0.3408319, -0.3408261, 
    -0.3408349, -0.3408344, -0.3408304, -0.3408345, -0.340766, -0.3407649, 
    -0.3407609, -0.340764, -0.3407584, -0.3407615, -0.3407633, -0.3407702, 
    -0.3407718, -0.3407858, -0.3407887, -0.3407923, -0.3408149, -0.3408205, 
    -0.3408256, -0.3408253, -0.3408254, -0.3408265, -0.3408237, -0.340827, 
    -0.3408275, -0.3408261, -0.3408344, -0.340832, -0.3408344, -0.3408329, 
    -0.3407652, -0.3407671, -0.3407661, -0.340768, -0.3407666, -0.3407852, 
    -0.340787, -0.3407956, -0.3407922, -0.3407978, -0.3407928, -0.3407936, 
    -0.3407978, -0.3407931, -0.3408202, -0.3407964, -0.3408266, -0.340819, 
    -0.340827, -0.3408256, -0.340828, -0.34083, -0.3408327, -0.3408374, 
    -0.3408364, -0.3408404, -0.3407699, -0.3407724, -0.3407722, -0.3407874, 
    -0.3407893, -0.3407936, -0.3408166, -0.3407977, -0.3408187, -0.3408197, 
    -0.3407963, -0.3408169, -0.3407866, -0.3407888, -0.3407876, -0.3407701, 
    -0.3407982, -0.3407902, -0.3408214, -0.3408171, -0.3408297, -0.3408234, 
    -0.3408358, -0.3408408, -0.340846, -0.3408516, -0.3407863, -0.3407721, 
    -0.3407877, -0.3407918, -0.3407958, -0.3408174, -0.3408179, -0.3408189, 
    -0.3408214, -0.3408235, -0.3408191, -0.3408241, -0.3407892, -0.3408153, 
    -0.3407714, -0.3407884, -0.3407916, -0.3407903, -0.3407975, -0.3408155, 
    -0.3408222, -0.3408188, -0.3408395, -0.3408304, -0.340856, -0.3408488, 
    -0.3407715, -0.3407864, -0.3407943, -0.3407905, -0.3408177, -0.3408204, 
    -0.3408226, -0.3408253, -0.3408256, -0.3408272, -0.3408246, -0.3408271, 
    -0.3408174, -0.3408217, -0.3407934, -0.3407963, -0.340795, -0.3407936, 
    -0.3407981, -0.3408192, -0.3408194, -0.3408209, -0.3408249, -0.3408178, 
    -0.3408405, -0.3408263, -0.3407889, -0.3407931, -0.3407939, -0.3407922, 
    -0.3408201, -0.3408159, -0.3408272, -0.3408242, -0.3408292, -0.3408267, 
    -0.3408263, -0.3408231, -0.3408211, -0.3408161, -0.3407956, -0.3407925, 
    -0.3407932, -0.3407967, -0.3408195, -0.3408256, -0.3408242, -0.3408288, 
    -0.3408169, -0.3408219, -0.3408199, -0.340825, -0.3407976, -0.340823, 
    -0.3407953, -0.3407963, -0.3408158, -0.3408221, -0.3408237, -0.3408251, 
    -0.3408242, -0.3408197, -0.3408189, -0.3408158, -0.3407985, -0.3407961, 
    -0.3407941, -0.3407959, -0.3407978, -0.3408197, -0.3408246, -0.34083, 
    -0.3408314, -0.3408374, -0.3408324, -0.3408406, -0.3408334, -0.3408459, 
    -0.3408237, -0.3408334, -0.340816, -0.3408179, -0.3408212, -0.3408291, 
    -0.340825, -0.3408298, -0.3408189, -0.3407968, -0.3407954, -0.3407926, 
    -0.3407955, -0.3407952, -0.3407979, -0.3407971, -0.3408199, -0.3408164, 
    -0.3408263, -0.3408298, -0.34084, -0.3408461, -0.3408525, -0.3408553, 
    -0.3408562, -0.3408565 ;

 TAUY =
  -0.3407592, -0.3407649, -0.3407638, -0.3407683, -0.3407659, -0.3407688, 
    -0.3407604, -0.3407651, -0.3407621, -0.3407598, -0.3407897, -0.3407685, 
    -0.3408154, -0.3407935, -0.3408239, -0.3407981, -0.3408258, -0.3408237, 
    -0.3408302, -0.3408284, -0.3408365, -0.3408311, -0.3408408, -0.3408352, 
    -0.3408361, -0.3408309, -0.3407704, -0.3407886, -0.34077, -0.3407708, 
    -0.3407705, -0.3407659, -0.3407635, -0.3407589, -0.3407597, -0.3407632, 
    -0.3407712, -0.3407685, -0.340788, -0.3407879, -0.3407956, -0.3407921, 
    -0.3408215, -0.3408178, -0.3408284, -0.3408258, -0.3408283, -0.3408276, 
    -0.3408283, -0.3408244, -0.3408261, -0.3408226, -0.3407927, -0.3407967, 
    -0.3407723, -0.3407651, -0.3407606, -0.3407573, -0.3407578, -0.3407587, 
    -0.3407632, -0.3407676, -0.3407709, -0.3407857, -0.3407879, -0.3407943, 
    -0.3407979, -0.3408222, -0.3408208, -0.3408231, -0.3408255, -0.3408293, 
    -0.3408287, -0.3408304, -0.3408231, -0.3408279, -0.34082, -0.3408222, 
    -0.3407881, -0.3407692, -0.3407663, -0.340764, -0.3407581, -0.3407622, 
    -0.3407606, -0.3407645, -0.3407669, -0.3407657, -0.3407857, -0.3407702, 
    -0.3407981, -0.3407915, -0.3408252, -0.3408211, -0.3408262, -0.3408236, 
    -0.3408281, -0.3408241, -0.340831, -0.3408325, -0.3408315, -0.3408355, 
    -0.3408238, -0.3408283, -0.3407657, -0.3407658, -0.3407668, -0.3407627, 
    -0.3407625, -0.3407588, -0.3407621, -0.3407634, -0.3407671, -0.3407691, 
    -0.3407711, -0.3407881, -0.340793, -0.3408163, -0.3408214, -0.3408247, 
    -0.3408227, -0.3408245, -0.3408225, -0.3408215, -0.3408319, -0.3408261, 
    -0.3408349, -0.3408344, -0.3408304, -0.3408345, -0.340766, -0.3407649, 
    -0.3407609, -0.340764, -0.3407584, -0.3407615, -0.3407633, -0.3407702, 
    -0.3407718, -0.3407858, -0.3407887, -0.3407923, -0.3408149, -0.3408205, 
    -0.3408256, -0.3408253, -0.3408254, -0.3408265, -0.3408237, -0.340827, 
    -0.3408275, -0.3408261, -0.3408344, -0.340832, -0.3408344, -0.3408329, 
    -0.3407652, -0.3407671, -0.3407661, -0.340768, -0.3407666, -0.3407852, 
    -0.340787, -0.3407956, -0.3407922, -0.3407978, -0.3407928, -0.3407936, 
    -0.3407978, -0.3407931, -0.3408202, -0.3407964, -0.3408266, -0.340819, 
    -0.340827, -0.3408256, -0.340828, -0.34083, -0.3408327, -0.3408374, 
    -0.3408364, -0.3408404, -0.3407699, -0.3407724, -0.3407722, -0.3407874, 
    -0.3407893, -0.3407936, -0.3408166, -0.3407977, -0.3408187, -0.3408197, 
    -0.3407963, -0.3408169, -0.3407866, -0.3407888, -0.3407876, -0.3407701, 
    -0.3407982, -0.3407902, -0.3408214, -0.3408171, -0.3408297, -0.3408234, 
    -0.3408358, -0.3408408, -0.340846, -0.3408516, -0.3407863, -0.3407721, 
    -0.3407877, -0.3407918, -0.3407958, -0.3408174, -0.3408179, -0.3408189, 
    -0.3408214, -0.3408235, -0.3408191, -0.3408241, -0.3407892, -0.3408153, 
    -0.3407714, -0.3407884, -0.3407916, -0.3407903, -0.3407975, -0.3408155, 
    -0.3408222, -0.3408188, -0.3408395, -0.3408304, -0.340856, -0.3408488, 
    -0.3407715, -0.3407864, -0.3407943, -0.3407905, -0.3408177, -0.3408204, 
    -0.3408226, -0.3408253, -0.3408256, -0.3408272, -0.3408246, -0.3408271, 
    -0.3408174, -0.3408217, -0.3407934, -0.3407963, -0.340795, -0.3407936, 
    -0.3407981, -0.3408192, -0.3408194, -0.3408209, -0.3408249, -0.3408178, 
    -0.3408405, -0.3408263, -0.3407889, -0.3407931, -0.3407939, -0.3407922, 
    -0.3408201, -0.3408159, -0.3408272, -0.3408242, -0.3408292, -0.3408267, 
    -0.3408263, -0.3408231, -0.3408211, -0.3408161, -0.3407956, -0.3407925, 
    -0.3407932, -0.3407967, -0.3408195, -0.3408256, -0.3408242, -0.3408288, 
    -0.3408169, -0.3408219, -0.3408199, -0.340825, -0.3407976, -0.340823, 
    -0.3407953, -0.3407963, -0.3408158, -0.3408221, -0.3408237, -0.3408251, 
    -0.3408242, -0.3408197, -0.3408189, -0.3408158, -0.3407985, -0.3407961, 
    -0.3407941, -0.3407959, -0.3407978, -0.3408197, -0.3408246, -0.34083, 
    -0.3408314, -0.3408374, -0.3408324, -0.3408406, -0.3408334, -0.3408459, 
    -0.3408237, -0.3408334, -0.340816, -0.3408179, -0.3408212, -0.3408291, 
    -0.340825, -0.3408298, -0.3408189, -0.3407968, -0.3407954, -0.3407926, 
    -0.3407955, -0.3407952, -0.3407979, -0.3407971, -0.3408199, -0.3408164, 
    -0.3408263, -0.3408298, -0.34084, -0.3408461, -0.3408525, -0.3408553, 
    -0.3408562, -0.3408565 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.4583, 261.4795, 261.4754, 261.4925, 261.483, 261.4942, 261.4626, 
    261.4803, 261.469, 261.4602, 261.5255, 261.4932, 261.559, 261.5385, 
    261.5902, 261.5559, 261.5971, 261.5892, 261.6131, 261.6062, 261.6367, 
    261.6162, 261.6525, 261.6318, 261.635, 261.6155, 261.4997, 261.5214, 
    261.4984, 261.5016, 261.5002, 261.4832, 261.4746, 261.4567, 261.46, 
    261.4731, 261.503, 261.4928, 261.5182, 261.5177, 261.5461, 261.5333, 
    261.5809, 261.5674, 261.6065, 261.5966, 261.606, 261.6032, 261.6061, 
    261.5916, 261.5978, 261.5851, 261.5357, 261.5502, 261.5069, 261.4807, 
    261.4634, 261.4511, 261.4528, 261.4561, 261.4732, 261.4892, 261.5015, 
    261.5096, 261.5176, 261.5419, 261.5548, 261.5836, 261.5784, 261.5872, 
    261.5957, 261.6098, 261.6075, 261.6137, 261.587, 261.6048, 261.5755, 
    261.5835, 261.5197, 261.4956, 261.4852, 261.4762, 261.4541, 261.4694, 
    261.4633, 261.4776, 261.4867, 261.4822, 261.5098, 261.4991, 261.5556, 
    261.5312, 261.5947, 261.5795, 261.5984, 261.5887, 261.6052, 261.5904, 
    261.6161, 261.6216, 261.6178, 261.6325, 261.5896, 261.606, 261.4821, 
    261.4828, 261.4862, 261.4713, 261.4703, 261.4566, 261.4688, 261.474, 
    261.4872, 261.495, 261.5024, 261.5186, 261.5368, 261.5622, 261.5805, 
    261.5927, 261.5852, 261.5919, 261.5844, 261.581, 261.6195, 261.5979, 
    261.6304, 261.6286, 261.6139, 261.6288, 261.4833, 261.4791, 261.4645, 
    261.476, 261.4551, 261.4668, 261.4735, 261.4993, 261.505, 261.5102, 
    261.5206, 261.5339, 261.5573, 261.5776, 261.5962, 261.5948, 261.5953, 
    261.5994, 261.5892, 261.6011, 261.6031, 261.5979, 261.6283, 261.6196, 
    261.6285, 261.6229, 261.4805, 261.4875, 261.4837, 261.4909, 261.4859, 
    261.5083, 261.515, 261.5466, 261.5337, 261.5543, 261.5358, 261.539, 
    261.5549, 261.5368, 261.5765, 261.5496, 261.5996, 261.5727, 261.6013, 
    261.5961, 261.6047, 261.6124, 261.6221, 261.64, 261.6358, 261.6508, 
    261.4981, 261.5073, 261.5065, 261.516, 261.5231, 261.5385, 261.5631, 
    261.5539, 261.5708, 261.5742, 261.5485, 261.5642, 261.5133, 261.5216, 
    261.5167, 261.4988, 261.556, 261.5266, 261.5808, 261.5649, 261.6113, 
    261.5882, 261.6335, 261.6529, 261.6711, 261.6924, 261.5122, 261.5061, 
    261.5172, 261.5326, 261.5469, 261.5659, 261.5678, 261.5714, 261.5806, 
    261.5884, 261.5725, 261.5903, 261.5235, 261.5585, 261.5037, 261.5201, 
    261.5316, 261.5266, 261.5528, 261.5589, 261.584, 261.571, 261.6481, 
    261.614, 261.7086, 261.6822, 261.5039, 261.5122, 261.5414, 261.5275, 
    261.5671, 261.5769, 261.5848, 261.595, 261.5961, 261.6021, 261.5923, 
    261.6017, 261.5659, 261.5819, 261.5381, 261.5487, 261.5438, 261.5384, 
    261.5551, 261.5727, 261.5731, 261.5788, 261.5948, 261.5673, 261.6525, 
    261.5999, 261.5213, 261.5375, 261.5398, 261.5335, 261.5759, 261.5605, 
    261.602, 261.5908, 261.6091, 261.6, 261.5986, 261.5869, 261.5797, 
    261.5612, 261.5463, 261.5345, 261.5372, 261.5503, 261.5738, 261.5962, 
    261.5913, 261.6077, 261.5642, 261.5825, 261.5754, 261.5938, 261.5536, 
    261.5878, 261.5449, 261.5486, 261.5602, 261.5837, 261.5889, 261.5945, 
    261.591, 261.5744, 261.5717, 261.56, 261.5568, 261.5478, 261.5404, 
    261.5472, 261.5543, 261.5744, 261.5927, 261.6125, 261.6174, 261.6405, 
    261.6216, 261.6527, 261.6263, 261.6721, 261.5898, 261.6255, 261.5608, 
    261.5677, 261.5804, 261.6093, 261.5937, 261.612, 261.5716, 261.5507, 
    261.5453, 261.5352, 261.5455, 261.5447, 261.5546, 261.5514, 261.5751, 
    261.5623, 261.5986, 261.6118, 261.6492, 261.6721, 261.6953, 261.7056, 
    261.7087, 261.7101 ;

 TG_R =
  261.4583, 261.4795, 261.4754, 261.4925, 261.483, 261.4942, 261.4626, 
    261.4803, 261.469, 261.4602, 261.5255, 261.4932, 261.559, 261.5385, 
    261.5902, 261.5559, 261.5971, 261.5892, 261.6131, 261.6062, 261.6367, 
    261.6162, 261.6525, 261.6318, 261.635, 261.6155, 261.4997, 261.5214, 
    261.4984, 261.5016, 261.5002, 261.4832, 261.4746, 261.4567, 261.46, 
    261.4731, 261.503, 261.4928, 261.5182, 261.5177, 261.5461, 261.5333, 
    261.5809, 261.5674, 261.6065, 261.5966, 261.606, 261.6032, 261.6061, 
    261.5916, 261.5978, 261.5851, 261.5357, 261.5502, 261.5069, 261.4807, 
    261.4634, 261.4511, 261.4528, 261.4561, 261.4732, 261.4892, 261.5015, 
    261.5096, 261.5176, 261.5419, 261.5548, 261.5836, 261.5784, 261.5872, 
    261.5957, 261.6098, 261.6075, 261.6137, 261.587, 261.6048, 261.5755, 
    261.5835, 261.5197, 261.4956, 261.4852, 261.4762, 261.4541, 261.4694, 
    261.4633, 261.4776, 261.4867, 261.4822, 261.5098, 261.4991, 261.5556, 
    261.5312, 261.5947, 261.5795, 261.5984, 261.5887, 261.6052, 261.5904, 
    261.6161, 261.6216, 261.6178, 261.6325, 261.5896, 261.606, 261.4821, 
    261.4828, 261.4862, 261.4713, 261.4703, 261.4566, 261.4688, 261.474, 
    261.4872, 261.495, 261.5024, 261.5186, 261.5368, 261.5622, 261.5805, 
    261.5927, 261.5852, 261.5919, 261.5844, 261.581, 261.6195, 261.5979, 
    261.6304, 261.6286, 261.6139, 261.6288, 261.4833, 261.4791, 261.4645, 
    261.476, 261.4551, 261.4668, 261.4735, 261.4993, 261.505, 261.5102, 
    261.5206, 261.5339, 261.5573, 261.5776, 261.5962, 261.5948, 261.5953, 
    261.5994, 261.5892, 261.6011, 261.6031, 261.5979, 261.6283, 261.6196, 
    261.6285, 261.6229, 261.4805, 261.4875, 261.4837, 261.4909, 261.4859, 
    261.5083, 261.515, 261.5466, 261.5337, 261.5543, 261.5358, 261.539, 
    261.5549, 261.5368, 261.5765, 261.5496, 261.5996, 261.5727, 261.6013, 
    261.5961, 261.6047, 261.6124, 261.6221, 261.64, 261.6358, 261.6508, 
    261.4981, 261.5073, 261.5065, 261.516, 261.5231, 261.5385, 261.5631, 
    261.5539, 261.5708, 261.5742, 261.5485, 261.5642, 261.5133, 261.5216, 
    261.5167, 261.4988, 261.556, 261.5266, 261.5808, 261.5649, 261.6113, 
    261.5882, 261.6335, 261.6529, 261.6711, 261.6924, 261.5122, 261.5061, 
    261.5172, 261.5326, 261.5469, 261.5659, 261.5678, 261.5714, 261.5806, 
    261.5884, 261.5725, 261.5903, 261.5235, 261.5585, 261.5037, 261.5201, 
    261.5316, 261.5266, 261.5528, 261.5589, 261.584, 261.571, 261.6481, 
    261.614, 261.7086, 261.6822, 261.5039, 261.5122, 261.5414, 261.5275, 
    261.5671, 261.5769, 261.5848, 261.595, 261.5961, 261.6021, 261.5923, 
    261.6017, 261.5659, 261.5819, 261.5381, 261.5487, 261.5438, 261.5384, 
    261.5551, 261.5727, 261.5731, 261.5788, 261.5948, 261.5673, 261.6525, 
    261.5999, 261.5213, 261.5375, 261.5398, 261.5335, 261.5759, 261.5605, 
    261.602, 261.5908, 261.6091, 261.6, 261.5986, 261.5869, 261.5797, 
    261.5612, 261.5463, 261.5345, 261.5372, 261.5503, 261.5738, 261.5962, 
    261.5913, 261.6077, 261.5642, 261.5825, 261.5754, 261.5938, 261.5536, 
    261.5878, 261.5449, 261.5486, 261.5602, 261.5837, 261.5889, 261.5945, 
    261.591, 261.5744, 261.5717, 261.56, 261.5568, 261.5478, 261.5404, 
    261.5472, 261.5543, 261.5744, 261.5927, 261.6125, 261.6174, 261.6405, 
    261.6216, 261.6527, 261.6263, 261.6721, 261.5898, 261.6255, 261.5608, 
    261.5677, 261.5804, 261.6093, 261.5937, 261.612, 261.5716, 261.5507, 
    261.5453, 261.5352, 261.5455, 261.5447, 261.5546, 261.5514, 261.5751, 
    261.5623, 261.5986, 261.6118, 261.6492, 261.6721, 261.6953, 261.7056, 
    261.7087, 261.7101 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.593, 254.5947, 254.5944, 254.5957, 254.595, 254.5959, 254.5933, 
    254.5948, 254.5939, 254.5932, 254.5984, 254.5958, 254.6012, 254.5995, 
    254.6037, 254.6009, 254.6043, 254.6036, 254.6056, 254.605, 254.6075, 
    254.6059, 254.6088, 254.6071, 254.6074, 254.6058, 254.5963, 254.5981, 
    254.5962, 254.5965, 254.5964, 254.595, 254.5943, 254.5929, 254.5931, 
    254.5942, 254.5966, 254.5958, 254.5979, 254.5978, 254.6001, 254.5991, 
    254.603, 254.6019, 254.6051, 254.6042, 254.605, 254.6048, 254.605, 
    254.6038, 254.6043, 254.6033, 254.5993, 254.6004, 254.5969, 254.5948, 
    254.5934, 254.5924, 254.5925, 254.5928, 254.5942, 254.5955, 254.5965, 
    254.5971, 254.5978, 254.5997, 254.6008, 254.6032, 254.6028, 254.6035, 
    254.6042, 254.6053, 254.6051, 254.6056, 254.6035, 254.6049, 254.6025, 
    254.6032, 254.5979, 254.596, 254.5951, 254.5944, 254.5927, 254.5939, 
    254.5934, 254.5946, 254.5953, 254.5949, 254.5972, 254.5963, 254.6009, 
    254.5989, 254.6041, 254.6028, 254.6044, 254.6036, 254.6049, 254.6037, 
    254.6058, 254.6063, 254.606, 254.6072, 254.6037, 254.605, 254.5949, 
    254.595, 254.5952, 254.594, 254.5939, 254.5928, 254.5938, 254.5943, 
    254.5953, 254.5959, 254.5966, 254.5979, 254.5993, 254.6014, 254.6029, 
    254.6039, 254.6033, 254.6039, 254.6032, 254.603, 254.6061, 254.6043, 
    254.607, 254.6069, 254.6057, 254.6069, 254.595, 254.5947, 254.5935, 
    254.5944, 254.5927, 254.5937, 254.5942, 254.5963, 254.5968, 254.5972, 
    254.598, 254.5991, 254.601, 254.6027, 254.6042, 254.6041, 254.6041, 
    254.6045, 254.6036, 254.6046, 254.6048, 254.6043, 254.6068, 254.6061, 
    254.6069, 254.6064, 254.5948, 254.5954, 254.595, 254.5956, 254.5952, 
    254.597, 254.5976, 254.6001, 254.5991, 254.6008, 254.5993, 254.5995, 
    254.6008, 254.5993, 254.6026, 254.6004, 254.6045, 254.6022, 254.6046, 
    254.6042, 254.6049, 254.6055, 254.6063, 254.6078, 254.6075, 254.6087, 
    254.5962, 254.5969, 254.5969, 254.5977, 254.5982, 254.5995, 254.6015, 
    254.6007, 254.6021, 254.6024, 254.6003, 254.6016, 254.5974, 254.5981, 
    254.5977, 254.5963, 254.6009, 254.5985, 254.6029, 254.6016, 254.6054, 
    254.6035, 254.6073, 254.6088, 254.6104, 254.6121, 254.5974, 254.5968, 
    254.5978, 254.599, 254.6002, 254.6017, 254.6019, 254.6022, 254.6029, 
    254.6036, 254.6022, 254.6037, 254.5982, 254.6011, 254.5966, 254.598, 
    254.5989, 254.5985, 254.6007, 254.6012, 254.6032, 254.6021, 254.6084, 
    254.6057, 254.6135, 254.6113, 254.5967, 254.5974, 254.5997, 254.5986, 
    254.6018, 254.6026, 254.6033, 254.6041, 254.6042, 254.6047, 254.6039, 
    254.6047, 254.6017, 254.603, 254.5995, 254.6003, 254.5999, 254.5995, 
    254.6008, 254.6023, 254.6023, 254.6028, 254.604, 254.6018, 254.6088, 
    254.6044, 254.5981, 254.5994, 254.5996, 254.5991, 254.6025, 254.6013, 
    254.6047, 254.6038, 254.6053, 254.6045, 254.6044, 254.6035, 254.6028, 
    254.6013, 254.6001, 254.5992, 254.5994, 254.6004, 254.6024, 254.6042, 
    254.6038, 254.6051, 254.6016, 254.6031, 254.6025, 254.604, 254.6007, 
    254.6035, 254.6, 254.6003, 254.6013, 254.6032, 254.6036, 254.604, 
    254.6038, 254.6024, 254.6022, 254.6012, 254.601, 254.6003, 254.5997, 
    254.6002, 254.6008, 254.6024, 254.6039, 254.6055, 254.6059, 254.6078, 
    254.6063, 254.6088, 254.6066, 254.6104, 254.6037, 254.6066, 254.6013, 
    254.6019, 254.6029, 254.6053, 254.604, 254.6055, 254.6022, 254.6005, 
    254.6001, 254.5992, 254.6001, 254.6, 254.6008, 254.6005, 254.6025, 
    254.6014, 254.6044, 254.6055, 254.6086, 254.6104, 254.6124, 254.6132, 
    254.6135, 254.6136 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24018, 18.24017, 18.24017, 18.24016, 18.24017, 18.24016, 18.24018, 
    18.24017, 18.24018, 18.24018, 18.24014, 18.24016, 18.24012, 18.24013, 
    18.2401, 18.24012, 18.2401, 18.2401, 18.24009, 18.24009, 18.24007, 
    18.24009, 18.24006, 18.24008, 18.24007, 18.24009, 18.24016, 18.24014, 
    18.24016, 18.24016, 18.24016, 18.24017, 18.24017, 18.24018, 18.24018, 
    18.24018, 18.24016, 18.24016, 18.24015, 18.24015, 18.24013, 18.24014, 
    18.24011, 18.24012, 18.24009, 18.2401, 18.24009, 18.24009, 18.24009, 
    18.2401, 18.2401, 18.2401, 18.24014, 18.24013, 18.24015, 18.24017, 
    18.24018, 18.24019, 18.24019, 18.24018, 18.24018, 18.24017, 18.24016, 
    18.24015, 18.24015, 18.24013, 18.24012, 18.24011, 18.24011, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24009, 18.2401, 18.24009, 18.24011, 
    18.24011, 18.24015, 18.24016, 18.24017, 18.24017, 18.24019, 18.24018, 
    18.24018, 18.24017, 18.24017, 18.24017, 18.24015, 18.24016, 18.24012, 
    18.24014, 18.2401, 18.24011, 18.2401, 18.2401, 18.24009, 18.2401, 
    18.24009, 18.24008, 18.24008, 18.24008, 18.2401, 18.24009, 18.24017, 
    18.24017, 18.24017, 18.24018, 18.24018, 18.24018, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24016, 18.24015, 18.24014, 18.24012, 18.24011, 
    18.2401, 18.2401, 18.2401, 18.2401, 18.24011, 18.24008, 18.2401, 
    18.24008, 18.24008, 18.24009, 18.24008, 18.24017, 18.24017, 18.24018, 
    18.24017, 18.24019, 18.24018, 18.24018, 18.24016, 18.24015, 18.24015, 
    18.24014, 18.24014, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.2401, 18.24008, 18.24008, 
    18.24008, 18.24008, 18.24017, 18.24017, 18.24017, 18.24016, 18.24017, 
    18.24015, 18.24015, 18.24013, 18.24014, 18.24012, 18.24014, 18.24013, 
    18.24012, 18.24014, 18.24011, 18.24013, 18.2401, 18.24011, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24008, 18.24007, 18.24007, 18.24006, 
    18.24016, 18.24015, 18.24015, 18.24015, 18.24014, 18.24013, 18.24012, 
    18.24012, 18.24011, 18.24011, 18.24013, 18.24012, 18.24015, 18.24014, 
    18.24015, 18.24016, 18.24012, 18.24014, 18.24011, 18.24012, 18.24009, 
    18.2401, 18.24007, 18.24006, 18.24005, 18.24004, 18.24015, 18.24015, 
    18.24015, 18.24014, 18.24013, 18.24012, 18.24012, 18.24011, 18.24011, 
    18.2401, 18.24011, 18.2401, 18.24014, 18.24012, 18.24016, 18.24014, 
    18.24014, 18.24014, 18.24013, 18.24012, 18.24011, 18.24011, 18.24007, 
    18.24009, 18.24003, 18.24004, 18.24016, 18.24015, 18.24013, 18.24014, 
    18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24012, 18.24011, 18.24014, 18.24013, 18.24013, 18.24013, 18.24012, 
    18.24011, 18.24011, 18.24011, 18.2401, 18.24012, 18.24006, 18.2401, 
    18.24014, 18.24014, 18.24013, 18.24014, 18.24011, 18.24012, 18.2401, 
    18.2401, 18.24009, 18.2401, 18.2401, 18.2401, 18.24011, 18.24012, 
    18.24013, 18.24014, 18.24014, 18.24013, 18.24011, 18.2401, 18.2401, 
    18.24009, 18.24012, 18.24011, 18.24011, 18.2401, 18.24012, 18.2401, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.24011, 18.24012, 18.24012, 18.24013, 18.24013, 18.24013, 
    18.24012, 18.24011, 18.2401, 18.24009, 18.24009, 18.24007, 18.24008, 
    18.24006, 18.24008, 18.24005, 18.2401, 18.24008, 18.24012, 18.24012, 
    18.24011, 18.24009, 18.2401, 18.24009, 18.24011, 18.24013, 18.24013, 
    18.24014, 18.24013, 18.24013, 18.24012, 18.24013, 18.24011, 18.24012, 
    18.2401, 18.24009, 18.24006, 18.24005, 18.24004, 18.24003, 18.24003, 
    18.24003 ;

 TOTCOLCH4 =
  1.442902e-05, 1.421366e-05, 1.425548e-05, 1.408212e-05, 1.417825e-05, 
    1.40648e-05, 1.438532e-05, 1.420511e-05, 1.432011e-05, 1.440963e-05, 
    1.374688e-05, 1.40744e-05, 1.340851e-05, 1.361611e-05, 1.309597e-05, 
    1.344075e-05, 1.302669e-05, 1.310592e-05, 1.286787e-05, 1.293597e-05, 
    1.263252e-05, 1.283647e-05, 1.247594e-05, 1.268118e-05, 1.264901e-05, 
    1.284321e-05, 1.400839e-05, 1.378756e-05, 1.402149e-05, 1.398996e-05, 
    1.400411e-05, 1.417625e-05, 1.426314e-05, 1.444553e-05, 1.441239e-05, 
    1.427845e-05, 1.397578e-05, 1.40784e-05, 1.382012e-05, 1.382595e-05, 
    1.353953e-05, 1.366852e-05, 1.318906e-05, 1.332496e-05, 1.293313e-05, 
    1.303142e-05, 1.293774e-05, 1.296613e-05, 1.293737e-05, 1.308159e-05, 
    1.301975e-05, 1.314683e-05, 1.364434e-05, 1.34977e-05, 1.393599e-05, 
    1.420086e-05, 1.43774e-05, 1.450292e-05, 1.448516e-05, 1.445131e-05, 
    1.427767e-05, 1.411481e-05, 1.399094e-05, 1.39082e-05, 1.382678e-05, 
    1.358085e-05, 1.345113e-05, 1.316161e-05, 1.321378e-05, 1.312544e-05, 
    1.304121e-05, 1.290003e-05, 1.292324e-05, 1.286112e-05, 1.312779e-05, 
    1.295042e-05, 1.324351e-05, 1.31632e-05, 1.380456e-05, 1.40507e-05, 
    1.41555e-05, 1.424744e-05, 1.447151e-05, 1.431669e-05, 1.437768e-05, 
    1.423269e-05, 1.414069e-05, 1.418618e-05, 1.390594e-05, 1.401475e-05, 
    1.344345e-05, 1.368892e-05, 1.305103e-05, 1.320307e-05, 1.301465e-05, 
    1.311072e-05, 1.294619e-05, 1.309425e-05, 1.283803e-05, 1.278238e-05, 
    1.28204e-05, 1.267453e-05, 1.310246e-05, 1.293773e-05, 1.418745e-05, 
    1.418003e-05, 1.414548e-05, 1.429749e-05, 1.43068e-05, 1.444643e-05, 
    1.432219e-05, 1.426933e-05, 1.413537e-05, 1.405623e-05, 1.398109e-05, 
    1.381618e-05, 1.363245e-05, 1.337645e-05, 1.31932e-05, 1.307067e-05, 
    1.314578e-05, 1.307947e-05, 1.31536e-05, 1.318839e-05, 1.280322e-05, 
    1.301917e-05, 1.269548e-05, 1.271335e-05, 1.285964e-05, 1.271134e-05, 
    1.417482e-05, 1.421753e-05, 1.436599e-05, 1.424978e-05, 1.446166e-05, 
    1.434297e-05, 1.427481e-05, 1.401246e-05, 1.395497e-05, 1.390168e-05, 
    1.379657e-05, 1.366191e-05, 1.342635e-05, 1.322213e-05, 1.303632e-05, 
    1.304991e-05, 1.304512e-05, 1.300368e-05, 1.310638e-05, 1.298684e-05, 
    1.296679e-05, 1.301921e-05, 1.271574e-05, 1.280227e-05, 1.271373e-05, 
    1.277006e-05, 1.420365e-05, 1.413181e-05, 1.417062e-05, 1.409766e-05, 
    1.414904e-05, 1.392081e-05, 1.385253e-05, 1.353398e-05, 1.366455e-05, 
    1.34569e-05, 1.364343e-05, 1.361034e-05, 1.345009e-05, 1.363335e-05, 
    1.323335e-05, 1.350422e-05, 1.300207e-05, 1.327148e-05, 1.298523e-05, 
    1.303712e-05, 1.295124e-05, 1.287442e-05, 1.277794e-05, 1.260034e-05, 
    1.264142e-05, 1.249324e-05, 1.402486e-05, 1.393193e-05, 1.394013e-05, 
    1.384301e-05, 1.377127e-05, 1.361607e-05, 1.336791e-05, 1.346112e-05, 
    1.329013e-05, 1.325585e-05, 1.351568e-05, 1.3356e-05, 1.386982e-05, 
    1.378651e-05, 1.383612e-05, 1.401752e-05, 1.34396e-05, 1.373555e-05, 
    1.319017e-05, 1.334969e-05, 1.288536e-05, 1.31158e-05, 1.266404e-05, 
    1.247199e-05, 1.229197e-05, 1.208229e-05, 1.388129e-05, 1.394437e-05, 
    1.383148e-05, 1.367556e-05, 1.353128e-05, 1.333994e-05, 1.332041e-05, 
    1.328463e-05, 1.319209e-05, 1.311439e-05, 1.327331e-05, 1.309493e-05, 
    1.376717e-05, 1.341399e-05, 1.396822e-05, 1.380081e-05, 1.368475e-05, 
    1.373565e-05, 1.347179e-05, 1.340975e-05, 1.315829e-05, 1.328816e-05, 
    1.251931e-05, 1.285818e-05, 1.19233e-05, 1.218283e-05, 1.396642e-05, 
    1.388151e-05, 1.358681e-05, 1.372687e-05, 1.33272e-05, 1.32292e-05, 
    1.314968e-05, 1.304814e-05, 1.30372e-05, 1.297714e-05, 1.307559e-05, 
    1.298103e-05, 1.333953e-05, 1.317906e-05, 1.362046e-05, 1.351272e-05, 
    1.356227e-05, 1.361664e-05, 1.344897e-05, 1.32708e-05, 1.326703e-05, 
    1.321e-05, 1.304955e-05, 1.332559e-05, 1.247567e-05, 1.2999e-05, 
    1.378904e-05, 1.362598e-05, 1.360277e-05, 1.366585e-05, 1.323902e-05, 
    1.339334e-05, 1.29786e-05, 1.309041e-05, 1.290734e-05, 1.299824e-05, 
    1.301162e-05, 1.312861e-05, 1.320155e-05, 1.338625e-05, 1.353694e-05, 
    1.36567e-05, 1.362884e-05, 1.349735e-05, 1.325992e-05, 1.30362e-05, 
    1.308513e-05, 1.292123e-05, 1.335609e-05, 1.317334e-05, 1.32439e-05, 
    1.30601e-05, 1.346359e-05, 1.311973e-05, 1.355178e-05, 1.351379e-05, 
    1.33964e-05, 1.316094e-05, 1.310902e-05, 1.305358e-05, 1.308779e-05, 
    1.325391e-05, 1.328119e-05, 1.339926e-05, 1.343189e-05, 1.352206e-05, 
    1.35968e-05, 1.35285e-05, 1.345685e-05, 1.325386e-05, 1.307149e-05, 
    1.287332e-05, 1.282494e-05, 1.25944e-05, 1.278195e-05, 1.247276e-05, 
    1.273545e-05, 1.228157e-05, 1.309991e-05, 1.274326e-05, 1.339108e-05, 
    1.332095e-05, 1.319429e-05, 1.290486e-05, 1.306097e-05, 1.287846e-05, 
    1.328226e-05, 1.34928e-05, 1.354743e-05, 1.364941e-05, 1.35451e-05, 
    1.355358e-05, 1.345391e-05, 1.348592e-05, 1.324713e-05, 1.337528e-05, 
    1.301195e-05, 1.287991e-05, 1.250874e-05, 1.228246e-05, 1.205319e-05, 
    1.19523e-05, 1.192164e-05, 1.190882e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24018, 18.24017, 18.24017, 18.24016, 18.24017, 18.24016, 18.24018, 
    18.24017, 18.24018, 18.24018, 18.24014, 18.24016, 18.24012, 18.24013, 
    18.2401, 18.24012, 18.2401, 18.2401, 18.24009, 18.24009, 18.24007, 
    18.24009, 18.24006, 18.24008, 18.24007, 18.24009, 18.24016, 18.24014, 
    18.24016, 18.24016, 18.24016, 18.24017, 18.24017, 18.24018, 18.24018, 
    18.24018, 18.24016, 18.24016, 18.24015, 18.24015, 18.24013, 18.24014, 
    18.24011, 18.24012, 18.24009, 18.2401, 18.24009, 18.24009, 18.24009, 
    18.2401, 18.2401, 18.2401, 18.24014, 18.24013, 18.24015, 18.24017, 
    18.24018, 18.24019, 18.24019, 18.24018, 18.24018, 18.24017, 18.24016, 
    18.24015, 18.24015, 18.24013, 18.24012, 18.24011, 18.24011, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24009, 18.2401, 18.24009, 18.24011, 
    18.24011, 18.24015, 18.24016, 18.24017, 18.24017, 18.24019, 18.24018, 
    18.24018, 18.24017, 18.24017, 18.24017, 18.24015, 18.24016, 18.24012, 
    18.24014, 18.2401, 18.24011, 18.2401, 18.2401, 18.24009, 18.2401, 
    18.24009, 18.24008, 18.24008, 18.24008, 18.2401, 18.24009, 18.24017, 
    18.24017, 18.24017, 18.24018, 18.24018, 18.24018, 18.24018, 18.24017, 
    18.24017, 18.24016, 18.24016, 18.24015, 18.24014, 18.24012, 18.24011, 
    18.2401, 18.2401, 18.2401, 18.2401, 18.24011, 18.24008, 18.2401, 
    18.24008, 18.24008, 18.24009, 18.24008, 18.24017, 18.24017, 18.24018, 
    18.24017, 18.24019, 18.24018, 18.24018, 18.24016, 18.24015, 18.24015, 
    18.24014, 18.24014, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.2401, 18.24008, 18.24008, 
    18.24008, 18.24008, 18.24017, 18.24017, 18.24017, 18.24016, 18.24017, 
    18.24015, 18.24015, 18.24013, 18.24014, 18.24012, 18.24014, 18.24013, 
    18.24012, 18.24014, 18.24011, 18.24013, 18.2401, 18.24011, 18.2401, 
    18.2401, 18.24009, 18.24009, 18.24008, 18.24007, 18.24007, 18.24006, 
    18.24016, 18.24015, 18.24015, 18.24015, 18.24014, 18.24013, 18.24012, 
    18.24012, 18.24011, 18.24011, 18.24013, 18.24012, 18.24015, 18.24014, 
    18.24015, 18.24016, 18.24012, 18.24014, 18.24011, 18.24012, 18.24009, 
    18.2401, 18.24007, 18.24006, 18.24005, 18.24004, 18.24015, 18.24015, 
    18.24015, 18.24014, 18.24013, 18.24012, 18.24012, 18.24011, 18.24011, 
    18.2401, 18.24011, 18.2401, 18.24014, 18.24012, 18.24016, 18.24014, 
    18.24014, 18.24014, 18.24013, 18.24012, 18.24011, 18.24011, 18.24007, 
    18.24009, 18.24003, 18.24004, 18.24016, 18.24015, 18.24013, 18.24014, 
    18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24012, 18.24011, 18.24014, 18.24013, 18.24013, 18.24013, 18.24012, 
    18.24011, 18.24011, 18.24011, 18.2401, 18.24012, 18.24006, 18.2401, 
    18.24014, 18.24014, 18.24013, 18.24014, 18.24011, 18.24012, 18.2401, 
    18.2401, 18.24009, 18.2401, 18.2401, 18.2401, 18.24011, 18.24012, 
    18.24013, 18.24014, 18.24014, 18.24013, 18.24011, 18.2401, 18.2401, 
    18.24009, 18.24012, 18.24011, 18.24011, 18.2401, 18.24012, 18.2401, 
    18.24013, 18.24013, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.24011, 18.24012, 18.24012, 18.24013, 18.24013, 18.24013, 
    18.24012, 18.24011, 18.2401, 18.24009, 18.24009, 18.24007, 18.24008, 
    18.24006, 18.24008, 18.24005, 18.2401, 18.24008, 18.24012, 18.24012, 
    18.24011, 18.24009, 18.2401, 18.24009, 18.24011, 18.24013, 18.24013, 
    18.24014, 18.24013, 18.24013, 18.24012, 18.24013, 18.24011, 18.24012, 
    18.2401, 18.24009, 18.24006, 18.24005, 18.24004, 18.24003, 18.24003, 
    18.24003 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976235e-05, 5.97622e-05, 5.976223e-05, 5.976211e-05, 5.976218e-05, 
    5.97621e-05, 5.976232e-05, 5.97622e-05, 5.976228e-05, 5.976234e-05, 
    5.976188e-05, 5.976211e-05, 5.976165e-05, 5.976179e-05, 5.976143e-05, 
    5.976167e-05, 5.976138e-05, 5.976143e-05, 5.976127e-05, 5.976131e-05, 
    5.97611e-05, 5.976125e-05, 5.976099e-05, 5.976114e-05, 5.976111e-05, 
    5.976125e-05, 5.976206e-05, 5.976191e-05, 5.976207e-05, 5.976205e-05, 
    5.976206e-05, 5.976218e-05, 5.976224e-05, 5.976236e-05, 5.976234e-05, 
    5.976225e-05, 5.976204e-05, 5.976211e-05, 5.976193e-05, 5.976194e-05, 
    5.976174e-05, 5.976183e-05, 5.976149e-05, 5.976159e-05, 5.976131e-05, 
    5.976138e-05, 5.976131e-05, 5.976134e-05, 5.976131e-05, 5.976142e-05, 
    5.976137e-05, 5.976146e-05, 5.976181e-05, 5.976171e-05, 5.976201e-05, 
    5.976219e-05, 5.976231e-05, 5.97624e-05, 5.976239e-05, 5.976237e-05, 
    5.976225e-05, 5.976214e-05, 5.976205e-05, 5.976199e-05, 5.976194e-05, 
    5.976177e-05, 5.976167e-05, 5.976147e-05, 5.976151e-05, 5.976145e-05, 
    5.976139e-05, 5.976129e-05, 5.976131e-05, 5.976126e-05, 5.976145e-05, 
    5.976133e-05, 5.976153e-05, 5.976147e-05, 5.976192e-05, 5.976209e-05, 
    5.976216e-05, 5.976223e-05, 5.976238e-05, 5.976227e-05, 5.976231e-05, 
    5.976222e-05, 5.976215e-05, 5.976218e-05, 5.976199e-05, 5.976207e-05, 
    5.976167e-05, 5.976184e-05, 5.976139e-05, 5.97615e-05, 5.976137e-05, 
    5.976144e-05, 5.976132e-05, 5.976143e-05, 5.976125e-05, 5.976121e-05, 
    5.976123e-05, 5.976113e-05, 5.976143e-05, 5.976131e-05, 5.976218e-05, 
    5.976218e-05, 5.976215e-05, 5.976226e-05, 5.976227e-05, 5.976237e-05, 
    5.976228e-05, 5.976224e-05, 5.976215e-05, 5.976209e-05, 5.976204e-05, 
    5.976193e-05, 5.97618e-05, 5.976162e-05, 5.97615e-05, 5.976141e-05, 
    5.976146e-05, 5.976142e-05, 5.976147e-05, 5.976149e-05, 5.976122e-05, 
    5.976137e-05, 5.976115e-05, 5.976116e-05, 5.976126e-05, 5.976116e-05, 
    5.976218e-05, 5.976221e-05, 5.976231e-05, 5.976223e-05, 5.976237e-05, 
    5.976229e-05, 5.976225e-05, 5.976206e-05, 5.976202e-05, 5.976199e-05, 
    5.976191e-05, 5.976182e-05, 5.976166e-05, 5.976151e-05, 5.976138e-05, 
    5.976139e-05, 5.976139e-05, 5.976136e-05, 5.976143e-05, 5.976135e-05, 
    5.976134e-05, 5.976137e-05, 5.976116e-05, 5.976122e-05, 5.976116e-05, 
    5.97612e-05, 5.976219e-05, 5.976215e-05, 5.976217e-05, 5.976212e-05, 
    5.976216e-05, 5.9762e-05, 5.976195e-05, 5.976173e-05, 5.976182e-05, 
    5.976168e-05, 5.976181e-05, 5.976178e-05, 5.976167e-05, 5.97618e-05, 
    5.976152e-05, 5.976171e-05, 5.976136e-05, 5.976155e-05, 5.976135e-05, 
    5.976139e-05, 5.976133e-05, 5.976127e-05, 5.976121e-05, 5.976108e-05, 
    5.976111e-05, 5.976101e-05, 5.976207e-05, 5.976201e-05, 5.976201e-05, 
    5.976195e-05, 5.97619e-05, 5.976179e-05, 5.976162e-05, 5.976168e-05, 
    5.976156e-05, 5.976154e-05, 5.976172e-05, 5.976161e-05, 5.976197e-05, 
    5.976191e-05, 5.976194e-05, 5.976207e-05, 5.976167e-05, 5.976187e-05, 
    5.976149e-05, 5.976161e-05, 5.976128e-05, 5.976144e-05, 5.976113e-05, 
    5.976099e-05, 5.976086e-05, 5.976071e-05, 5.976197e-05, 5.976202e-05, 
    5.976194e-05, 5.976183e-05, 5.976173e-05, 5.97616e-05, 5.976158e-05, 
    5.976156e-05, 5.976149e-05, 5.976144e-05, 5.976155e-05, 5.976143e-05, 
    5.976189e-05, 5.976165e-05, 5.976203e-05, 5.976192e-05, 5.976184e-05, 
    5.976187e-05, 5.976169e-05, 5.976165e-05, 5.976147e-05, 5.976156e-05, 
    5.976102e-05, 5.976126e-05, 5.97606e-05, 5.976078e-05, 5.976203e-05, 
    5.976197e-05, 5.976177e-05, 5.976187e-05, 5.976159e-05, 5.976152e-05, 
    5.976146e-05, 5.976139e-05, 5.976139e-05, 5.976134e-05, 5.976141e-05, 
    5.976135e-05, 5.97616e-05, 5.976149e-05, 5.976179e-05, 5.976172e-05, 
    5.976175e-05, 5.976179e-05, 5.976167e-05, 5.976155e-05, 5.976155e-05, 
    5.976151e-05, 5.976139e-05, 5.976159e-05, 5.976099e-05, 5.976136e-05, 
    5.976191e-05, 5.976179e-05, 5.976178e-05, 5.976182e-05, 5.976153e-05, 
    5.976163e-05, 5.976134e-05, 5.976142e-05, 5.97613e-05, 5.976136e-05, 
    5.976137e-05, 5.976145e-05, 5.97615e-05, 5.976163e-05, 5.976173e-05, 
    5.976182e-05, 5.97618e-05, 5.976171e-05, 5.976154e-05, 5.976138e-05, 
    5.976142e-05, 5.97613e-05, 5.976161e-05, 5.976148e-05, 5.976153e-05, 
    5.97614e-05, 5.976168e-05, 5.976145e-05, 5.976174e-05, 5.976172e-05, 
    5.976164e-05, 5.976147e-05, 5.976143e-05, 5.97614e-05, 5.976142e-05, 
    5.976154e-05, 5.976155e-05, 5.976164e-05, 5.976166e-05, 5.976173e-05, 
    5.976178e-05, 5.976173e-05, 5.976168e-05, 5.976154e-05, 5.976141e-05, 
    5.976127e-05, 5.976124e-05, 5.976107e-05, 5.976121e-05, 5.976099e-05, 
    5.976118e-05, 5.976086e-05, 5.976143e-05, 5.976118e-05, 5.976163e-05, 
    5.976158e-05, 5.97615e-05, 5.976129e-05, 5.97614e-05, 5.976127e-05, 
    5.976156e-05, 5.97617e-05, 5.976174e-05, 5.976181e-05, 5.976174e-05, 
    5.976175e-05, 5.976168e-05, 5.97617e-05, 5.976153e-05, 5.976162e-05, 
    5.976137e-05, 5.976127e-05, 5.976102e-05, 5.976086e-05, 5.976069e-05, 
    5.976062e-05, 5.97606e-05, 5.976059e-05 ;

 TOTLITC_1m =
  5.976235e-05, 5.97622e-05, 5.976223e-05, 5.976211e-05, 5.976218e-05, 
    5.97621e-05, 5.976232e-05, 5.97622e-05, 5.976228e-05, 5.976234e-05, 
    5.976188e-05, 5.976211e-05, 5.976165e-05, 5.976179e-05, 5.976143e-05, 
    5.976167e-05, 5.976138e-05, 5.976143e-05, 5.976127e-05, 5.976131e-05, 
    5.97611e-05, 5.976125e-05, 5.976099e-05, 5.976114e-05, 5.976111e-05, 
    5.976125e-05, 5.976206e-05, 5.976191e-05, 5.976207e-05, 5.976205e-05, 
    5.976206e-05, 5.976218e-05, 5.976224e-05, 5.976236e-05, 5.976234e-05, 
    5.976225e-05, 5.976204e-05, 5.976211e-05, 5.976193e-05, 5.976194e-05, 
    5.976174e-05, 5.976183e-05, 5.976149e-05, 5.976159e-05, 5.976131e-05, 
    5.976138e-05, 5.976131e-05, 5.976134e-05, 5.976131e-05, 5.976142e-05, 
    5.976137e-05, 5.976146e-05, 5.976181e-05, 5.976171e-05, 5.976201e-05, 
    5.976219e-05, 5.976231e-05, 5.97624e-05, 5.976239e-05, 5.976237e-05, 
    5.976225e-05, 5.976214e-05, 5.976205e-05, 5.976199e-05, 5.976194e-05, 
    5.976177e-05, 5.976167e-05, 5.976147e-05, 5.976151e-05, 5.976145e-05, 
    5.976139e-05, 5.976129e-05, 5.976131e-05, 5.976126e-05, 5.976145e-05, 
    5.976133e-05, 5.976153e-05, 5.976147e-05, 5.976192e-05, 5.976209e-05, 
    5.976216e-05, 5.976223e-05, 5.976238e-05, 5.976227e-05, 5.976231e-05, 
    5.976222e-05, 5.976215e-05, 5.976218e-05, 5.976199e-05, 5.976207e-05, 
    5.976167e-05, 5.976184e-05, 5.976139e-05, 5.97615e-05, 5.976137e-05, 
    5.976144e-05, 5.976132e-05, 5.976143e-05, 5.976125e-05, 5.976121e-05, 
    5.976123e-05, 5.976113e-05, 5.976143e-05, 5.976131e-05, 5.976218e-05, 
    5.976218e-05, 5.976215e-05, 5.976226e-05, 5.976227e-05, 5.976237e-05, 
    5.976228e-05, 5.976224e-05, 5.976215e-05, 5.976209e-05, 5.976204e-05, 
    5.976193e-05, 5.97618e-05, 5.976162e-05, 5.97615e-05, 5.976141e-05, 
    5.976146e-05, 5.976142e-05, 5.976147e-05, 5.976149e-05, 5.976122e-05, 
    5.976137e-05, 5.976115e-05, 5.976116e-05, 5.976126e-05, 5.976116e-05, 
    5.976218e-05, 5.976221e-05, 5.976231e-05, 5.976223e-05, 5.976237e-05, 
    5.976229e-05, 5.976225e-05, 5.976206e-05, 5.976202e-05, 5.976199e-05, 
    5.976191e-05, 5.976182e-05, 5.976166e-05, 5.976151e-05, 5.976138e-05, 
    5.976139e-05, 5.976139e-05, 5.976136e-05, 5.976143e-05, 5.976135e-05, 
    5.976134e-05, 5.976137e-05, 5.976116e-05, 5.976122e-05, 5.976116e-05, 
    5.97612e-05, 5.976219e-05, 5.976215e-05, 5.976217e-05, 5.976212e-05, 
    5.976216e-05, 5.9762e-05, 5.976195e-05, 5.976173e-05, 5.976182e-05, 
    5.976168e-05, 5.976181e-05, 5.976178e-05, 5.976167e-05, 5.97618e-05, 
    5.976152e-05, 5.976171e-05, 5.976136e-05, 5.976155e-05, 5.976135e-05, 
    5.976139e-05, 5.976133e-05, 5.976127e-05, 5.976121e-05, 5.976108e-05, 
    5.976111e-05, 5.976101e-05, 5.976207e-05, 5.976201e-05, 5.976201e-05, 
    5.976195e-05, 5.97619e-05, 5.976179e-05, 5.976162e-05, 5.976168e-05, 
    5.976156e-05, 5.976154e-05, 5.976172e-05, 5.976161e-05, 5.976197e-05, 
    5.976191e-05, 5.976194e-05, 5.976207e-05, 5.976167e-05, 5.976187e-05, 
    5.976149e-05, 5.976161e-05, 5.976128e-05, 5.976144e-05, 5.976113e-05, 
    5.976099e-05, 5.976086e-05, 5.976071e-05, 5.976197e-05, 5.976202e-05, 
    5.976194e-05, 5.976183e-05, 5.976173e-05, 5.97616e-05, 5.976158e-05, 
    5.976156e-05, 5.976149e-05, 5.976144e-05, 5.976155e-05, 5.976143e-05, 
    5.976189e-05, 5.976165e-05, 5.976203e-05, 5.976192e-05, 5.976184e-05, 
    5.976187e-05, 5.976169e-05, 5.976165e-05, 5.976147e-05, 5.976156e-05, 
    5.976102e-05, 5.976126e-05, 5.97606e-05, 5.976078e-05, 5.976203e-05, 
    5.976197e-05, 5.976177e-05, 5.976187e-05, 5.976159e-05, 5.976152e-05, 
    5.976146e-05, 5.976139e-05, 5.976139e-05, 5.976134e-05, 5.976141e-05, 
    5.976135e-05, 5.97616e-05, 5.976149e-05, 5.976179e-05, 5.976172e-05, 
    5.976175e-05, 5.976179e-05, 5.976167e-05, 5.976155e-05, 5.976155e-05, 
    5.976151e-05, 5.976139e-05, 5.976159e-05, 5.976099e-05, 5.976136e-05, 
    5.976191e-05, 5.976179e-05, 5.976178e-05, 5.976182e-05, 5.976153e-05, 
    5.976163e-05, 5.976134e-05, 5.976142e-05, 5.97613e-05, 5.976136e-05, 
    5.976137e-05, 5.976145e-05, 5.97615e-05, 5.976163e-05, 5.976173e-05, 
    5.976182e-05, 5.97618e-05, 5.976171e-05, 5.976154e-05, 5.976138e-05, 
    5.976142e-05, 5.97613e-05, 5.976161e-05, 5.976148e-05, 5.976153e-05, 
    5.97614e-05, 5.976168e-05, 5.976145e-05, 5.976174e-05, 5.976172e-05, 
    5.976164e-05, 5.976147e-05, 5.976143e-05, 5.97614e-05, 5.976142e-05, 
    5.976154e-05, 5.976155e-05, 5.976164e-05, 5.976166e-05, 5.976173e-05, 
    5.976178e-05, 5.976173e-05, 5.976168e-05, 5.976154e-05, 5.976141e-05, 
    5.976127e-05, 5.976124e-05, 5.976107e-05, 5.976121e-05, 5.976099e-05, 
    5.976118e-05, 5.976086e-05, 5.976143e-05, 5.976118e-05, 5.976163e-05, 
    5.976158e-05, 5.97615e-05, 5.976129e-05, 5.97614e-05, 5.976127e-05, 
    5.976156e-05, 5.97617e-05, 5.976174e-05, 5.976181e-05, 5.976174e-05, 
    5.976175e-05, 5.976168e-05, 5.97617e-05, 5.976153e-05, 5.976162e-05, 
    5.976137e-05, 5.976127e-05, 5.976102e-05, 5.976086e-05, 5.976069e-05, 
    5.976062e-05, 5.97606e-05, 5.976059e-05 ;

 TOTLITN =
  1.375938e-06, 1.375934e-06, 1.375935e-06, 1.375931e-06, 1.375933e-06, 
    1.375931e-06, 1.375937e-06, 1.375934e-06, 1.375936e-06, 1.375938e-06, 
    1.375925e-06, 1.375931e-06, 1.375918e-06, 1.375922e-06, 1.375912e-06, 
    1.375919e-06, 1.375911e-06, 1.375912e-06, 1.375908e-06, 1.375909e-06, 
    1.375903e-06, 1.375907e-06, 1.3759e-06, 1.375904e-06, 1.375903e-06, 
    1.375907e-06, 1.37593e-06, 1.375926e-06, 1.37593e-06, 1.37593e-06, 
    1.37593e-06, 1.375933e-06, 1.375935e-06, 1.375938e-06, 1.375938e-06, 
    1.375935e-06, 1.375929e-06, 1.375931e-06, 1.375926e-06, 1.375926e-06, 
    1.375921e-06, 1.375923e-06, 1.375914e-06, 1.375917e-06, 1.375909e-06, 
    1.375911e-06, 1.375909e-06, 1.37591e-06, 1.375909e-06, 1.375912e-06, 
    1.375911e-06, 1.375913e-06, 1.375923e-06, 1.37592e-06, 1.375928e-06, 
    1.375934e-06, 1.375937e-06, 1.37594e-06, 1.375939e-06, 1.375938e-06, 
    1.375935e-06, 1.375932e-06, 1.37593e-06, 1.375928e-06, 1.375926e-06, 
    1.375922e-06, 1.375919e-06, 1.375913e-06, 1.375914e-06, 1.375913e-06, 
    1.375911e-06, 1.375908e-06, 1.375909e-06, 1.375907e-06, 1.375913e-06, 
    1.375909e-06, 1.375915e-06, 1.375913e-06, 1.375926e-06, 1.375931e-06, 
    1.375933e-06, 1.375935e-06, 1.375939e-06, 1.375936e-06, 1.375937e-06, 
    1.375934e-06, 1.375932e-06, 1.375933e-06, 1.375928e-06, 1.37593e-06, 
    1.375919e-06, 1.375924e-06, 1.375911e-06, 1.375914e-06, 1.37591e-06, 
    1.375912e-06, 1.375909e-06, 1.375912e-06, 1.375907e-06, 1.375906e-06, 
    1.375907e-06, 1.375904e-06, 1.375912e-06, 1.375909e-06, 1.375933e-06, 
    1.375933e-06, 1.375933e-06, 1.375936e-06, 1.375936e-06, 1.375938e-06, 
    1.375936e-06, 1.375935e-06, 1.375932e-06, 1.375931e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.375918e-06, 1.375914e-06, 1.375912e-06, 
    1.375913e-06, 1.375912e-06, 1.375913e-06, 1.375914e-06, 1.375906e-06, 
    1.375911e-06, 1.375904e-06, 1.375905e-06, 1.375907e-06, 1.375904e-06, 
    1.375933e-06, 1.375934e-06, 1.375937e-06, 1.375935e-06, 1.375939e-06, 
    1.375936e-06, 1.375935e-06, 1.37593e-06, 1.375929e-06, 1.375928e-06, 
    1.375926e-06, 1.375923e-06, 1.375918e-06, 1.375915e-06, 1.375911e-06, 
    1.375911e-06, 1.375911e-06, 1.37591e-06, 1.375912e-06, 1.37591e-06, 
    1.37591e-06, 1.375911e-06, 1.375905e-06, 1.375906e-06, 1.375905e-06, 
    1.375906e-06, 1.375934e-06, 1.375932e-06, 1.375933e-06, 1.375932e-06, 
    1.375933e-06, 1.375928e-06, 1.375927e-06, 1.375921e-06, 1.375923e-06, 
    1.375919e-06, 1.375923e-06, 1.375922e-06, 1.375919e-06, 1.375923e-06, 
    1.375915e-06, 1.37592e-06, 1.37591e-06, 1.375916e-06, 1.37591e-06, 
    1.375911e-06, 1.375909e-06, 1.375908e-06, 1.375906e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.37593e-06, 1.375928e-06, 1.375929e-06, 
    1.375927e-06, 1.375925e-06, 1.375922e-06, 1.375917e-06, 1.375919e-06, 
    1.375916e-06, 1.375915e-06, 1.37592e-06, 1.375917e-06, 1.375927e-06, 
    1.375926e-06, 1.375927e-06, 1.37593e-06, 1.375919e-06, 1.375925e-06, 
    1.375914e-06, 1.375917e-06, 1.375908e-06, 1.375912e-06, 1.375903e-06, 
    1.3759e-06, 1.375896e-06, 1.375892e-06, 1.375927e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.375921e-06, 1.375917e-06, 1.375916e-06, 
    1.375916e-06, 1.375914e-06, 1.375912e-06, 1.375916e-06, 1.375912e-06, 
    1.375925e-06, 1.375918e-06, 1.375929e-06, 1.375926e-06, 1.375924e-06, 
    1.375925e-06, 1.375919e-06, 1.375918e-06, 1.375913e-06, 1.375916e-06, 
    1.375901e-06, 1.375907e-06, 1.375889e-06, 1.375894e-06, 1.375929e-06, 
    1.375927e-06, 1.375922e-06, 1.375924e-06, 1.375917e-06, 1.375915e-06, 
    1.375913e-06, 1.375911e-06, 1.375911e-06, 1.37591e-06, 1.375912e-06, 
    1.37591e-06, 1.375917e-06, 1.375914e-06, 1.375922e-06, 1.37592e-06, 
    1.375921e-06, 1.375922e-06, 1.375919e-06, 1.375915e-06, 1.375915e-06, 
    1.375914e-06, 1.375911e-06, 1.375917e-06, 1.3759e-06, 1.37591e-06, 
    1.375926e-06, 1.375922e-06, 1.375922e-06, 1.375923e-06, 1.375915e-06, 
    1.375918e-06, 1.37591e-06, 1.375912e-06, 1.375908e-06, 1.37591e-06, 
    1.37591e-06, 1.375913e-06, 1.375914e-06, 1.375918e-06, 1.375921e-06, 
    1.375923e-06, 1.375922e-06, 1.37592e-06, 1.375915e-06, 1.375911e-06, 
    1.375912e-06, 1.375909e-06, 1.375917e-06, 1.375914e-06, 1.375915e-06, 
    1.375911e-06, 1.375919e-06, 1.375912e-06, 1.375921e-06, 1.37592e-06, 
    1.375918e-06, 1.375913e-06, 1.375912e-06, 1.375911e-06, 1.375912e-06, 
    1.375915e-06, 1.375916e-06, 1.375918e-06, 1.375919e-06, 1.37592e-06, 
    1.375922e-06, 1.375921e-06, 1.375919e-06, 1.375915e-06, 1.375912e-06, 
    1.375908e-06, 1.375907e-06, 1.375902e-06, 1.375906e-06, 1.3759e-06, 
    1.375905e-06, 1.375896e-06, 1.375912e-06, 1.375905e-06, 1.375918e-06, 
    1.375916e-06, 1.375914e-06, 1.375908e-06, 1.375911e-06, 1.375908e-06, 
    1.375916e-06, 1.37592e-06, 1.375921e-06, 1.375923e-06, 1.375921e-06, 
    1.375921e-06, 1.375919e-06, 1.37592e-06, 1.375915e-06, 1.375917e-06, 
    1.37591e-06, 1.375908e-06, 1.3759e-06, 1.375896e-06, 1.375891e-06, 
    1.375889e-06, 1.375889e-06, 1.375888e-06 ;

 TOTLITN_1m =
  1.375938e-06, 1.375934e-06, 1.375935e-06, 1.375931e-06, 1.375933e-06, 
    1.375931e-06, 1.375937e-06, 1.375934e-06, 1.375936e-06, 1.375938e-06, 
    1.375925e-06, 1.375931e-06, 1.375918e-06, 1.375922e-06, 1.375912e-06, 
    1.375919e-06, 1.375911e-06, 1.375912e-06, 1.375908e-06, 1.375909e-06, 
    1.375903e-06, 1.375907e-06, 1.3759e-06, 1.375904e-06, 1.375903e-06, 
    1.375907e-06, 1.37593e-06, 1.375926e-06, 1.37593e-06, 1.37593e-06, 
    1.37593e-06, 1.375933e-06, 1.375935e-06, 1.375938e-06, 1.375938e-06, 
    1.375935e-06, 1.375929e-06, 1.375931e-06, 1.375926e-06, 1.375926e-06, 
    1.375921e-06, 1.375923e-06, 1.375914e-06, 1.375917e-06, 1.375909e-06, 
    1.375911e-06, 1.375909e-06, 1.37591e-06, 1.375909e-06, 1.375912e-06, 
    1.375911e-06, 1.375913e-06, 1.375923e-06, 1.37592e-06, 1.375928e-06, 
    1.375934e-06, 1.375937e-06, 1.37594e-06, 1.375939e-06, 1.375938e-06, 
    1.375935e-06, 1.375932e-06, 1.37593e-06, 1.375928e-06, 1.375926e-06, 
    1.375922e-06, 1.375919e-06, 1.375913e-06, 1.375914e-06, 1.375913e-06, 
    1.375911e-06, 1.375908e-06, 1.375909e-06, 1.375907e-06, 1.375913e-06, 
    1.375909e-06, 1.375915e-06, 1.375913e-06, 1.375926e-06, 1.375931e-06, 
    1.375933e-06, 1.375935e-06, 1.375939e-06, 1.375936e-06, 1.375937e-06, 
    1.375934e-06, 1.375932e-06, 1.375933e-06, 1.375928e-06, 1.37593e-06, 
    1.375919e-06, 1.375924e-06, 1.375911e-06, 1.375914e-06, 1.37591e-06, 
    1.375912e-06, 1.375909e-06, 1.375912e-06, 1.375907e-06, 1.375906e-06, 
    1.375907e-06, 1.375904e-06, 1.375912e-06, 1.375909e-06, 1.375933e-06, 
    1.375933e-06, 1.375933e-06, 1.375936e-06, 1.375936e-06, 1.375938e-06, 
    1.375936e-06, 1.375935e-06, 1.375932e-06, 1.375931e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.375918e-06, 1.375914e-06, 1.375912e-06, 
    1.375913e-06, 1.375912e-06, 1.375913e-06, 1.375914e-06, 1.375906e-06, 
    1.375911e-06, 1.375904e-06, 1.375905e-06, 1.375907e-06, 1.375904e-06, 
    1.375933e-06, 1.375934e-06, 1.375937e-06, 1.375935e-06, 1.375939e-06, 
    1.375936e-06, 1.375935e-06, 1.37593e-06, 1.375929e-06, 1.375928e-06, 
    1.375926e-06, 1.375923e-06, 1.375918e-06, 1.375915e-06, 1.375911e-06, 
    1.375911e-06, 1.375911e-06, 1.37591e-06, 1.375912e-06, 1.37591e-06, 
    1.37591e-06, 1.375911e-06, 1.375905e-06, 1.375906e-06, 1.375905e-06, 
    1.375906e-06, 1.375934e-06, 1.375932e-06, 1.375933e-06, 1.375932e-06, 
    1.375933e-06, 1.375928e-06, 1.375927e-06, 1.375921e-06, 1.375923e-06, 
    1.375919e-06, 1.375923e-06, 1.375922e-06, 1.375919e-06, 1.375923e-06, 
    1.375915e-06, 1.37592e-06, 1.37591e-06, 1.375916e-06, 1.37591e-06, 
    1.375911e-06, 1.375909e-06, 1.375908e-06, 1.375906e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.37593e-06, 1.375928e-06, 1.375929e-06, 
    1.375927e-06, 1.375925e-06, 1.375922e-06, 1.375917e-06, 1.375919e-06, 
    1.375916e-06, 1.375915e-06, 1.37592e-06, 1.375917e-06, 1.375927e-06, 
    1.375926e-06, 1.375927e-06, 1.37593e-06, 1.375919e-06, 1.375925e-06, 
    1.375914e-06, 1.375917e-06, 1.375908e-06, 1.375912e-06, 1.375903e-06, 
    1.3759e-06, 1.375896e-06, 1.375892e-06, 1.375927e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.375921e-06, 1.375917e-06, 1.375916e-06, 
    1.375916e-06, 1.375914e-06, 1.375912e-06, 1.375916e-06, 1.375912e-06, 
    1.375925e-06, 1.375918e-06, 1.375929e-06, 1.375926e-06, 1.375924e-06, 
    1.375925e-06, 1.375919e-06, 1.375918e-06, 1.375913e-06, 1.375916e-06, 
    1.375901e-06, 1.375907e-06, 1.375889e-06, 1.375894e-06, 1.375929e-06, 
    1.375927e-06, 1.375922e-06, 1.375924e-06, 1.375917e-06, 1.375915e-06, 
    1.375913e-06, 1.375911e-06, 1.375911e-06, 1.37591e-06, 1.375912e-06, 
    1.37591e-06, 1.375917e-06, 1.375914e-06, 1.375922e-06, 1.37592e-06, 
    1.375921e-06, 1.375922e-06, 1.375919e-06, 1.375915e-06, 1.375915e-06, 
    1.375914e-06, 1.375911e-06, 1.375917e-06, 1.3759e-06, 1.37591e-06, 
    1.375926e-06, 1.375922e-06, 1.375922e-06, 1.375923e-06, 1.375915e-06, 
    1.375918e-06, 1.37591e-06, 1.375912e-06, 1.375908e-06, 1.37591e-06, 
    1.37591e-06, 1.375913e-06, 1.375914e-06, 1.375918e-06, 1.375921e-06, 
    1.375923e-06, 1.375922e-06, 1.37592e-06, 1.375915e-06, 1.375911e-06, 
    1.375912e-06, 1.375909e-06, 1.375917e-06, 1.375914e-06, 1.375915e-06, 
    1.375911e-06, 1.375919e-06, 1.375912e-06, 1.375921e-06, 1.37592e-06, 
    1.375918e-06, 1.375913e-06, 1.375912e-06, 1.375911e-06, 1.375912e-06, 
    1.375915e-06, 1.375916e-06, 1.375918e-06, 1.375919e-06, 1.37592e-06, 
    1.375922e-06, 1.375921e-06, 1.375919e-06, 1.375915e-06, 1.375912e-06, 
    1.375908e-06, 1.375907e-06, 1.375902e-06, 1.375906e-06, 1.3759e-06, 
    1.375905e-06, 1.375896e-06, 1.375912e-06, 1.375905e-06, 1.375918e-06, 
    1.375916e-06, 1.375914e-06, 1.375908e-06, 1.375911e-06, 1.375908e-06, 
    1.375916e-06, 1.37592e-06, 1.375921e-06, 1.375923e-06, 1.375921e-06, 
    1.375921e-06, 1.375919e-06, 1.37592e-06, 1.375915e-06, 1.375917e-06, 
    1.37591e-06, 1.375908e-06, 1.3759e-06, 1.375896e-06, 1.375891e-06, 
    1.375889e-06, 1.375889e-06, 1.375888e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.3448, 17.34479, 17.34479, 17.34478, 17.34479, 17.34478, 17.3448, 
    17.34479, 17.3448, 17.3448, 17.34476, 17.34478, 17.34474, 17.34475, 
    17.34472, 17.34474, 17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34468, 17.3447, 17.34469, 17.34471, 17.34478, 17.34476, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.34479, 17.3448, 17.3448, 
    17.3448, 17.34478, 17.34478, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34471, 17.34472, 17.34471, 17.34471, 17.34471, 
    17.34472, 17.34472, 17.34472, 17.34476, 17.34475, 17.34477, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 
    17.34477, 17.34477, 17.34475, 17.34474, 17.34472, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.34471, 17.34472, 17.34471, 17.34473, 
    17.34472, 17.34476, 17.34478, 17.34479, 17.34479, 17.34481, 17.3448, 
    17.3448, 17.34479, 17.34479, 17.34479, 17.34477, 17.34478, 17.34474, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34472, 17.34471, 17.34472, 
    17.34471, 17.3447, 17.3447, 17.34469, 17.34472, 17.34471, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.3448, 17.3448, 17.34479, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34472, 17.34473, 17.3447, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.3448, 17.34479, 17.34478, 17.34477, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34472, 17.3447, 17.3447, 
    17.3447, 17.3447, 17.34479, 17.34479, 17.34479, 17.34478, 17.34479, 
    17.34477, 17.34477, 17.34475, 17.34476, 17.34474, 17.34476, 17.34475, 
    17.34474, 17.34476, 17.34473, 17.34475, 17.34472, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.34469, 17.34469, 17.34468, 
    17.34478, 17.34477, 17.34477, 17.34477, 17.34476, 17.34475, 17.34474, 
    17.34474, 17.34473, 17.34473, 17.34475, 17.34474, 17.34477, 17.34476, 
    17.34477, 17.34478, 17.34474, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34472, 17.34469, 17.34468, 17.34467, 17.34466, 17.34477, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34476, 17.34474, 17.34478, 17.34476, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34472, 17.34473, 17.34468, 
    17.34471, 17.34465, 17.34466, 17.34478, 17.34477, 17.34475, 17.34476, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34471, 17.34472, 
    17.34471, 17.34474, 17.34473, 17.34475, 17.34475, 17.34475, 17.34475, 
    17.34474, 17.34473, 17.34473, 17.34473, 17.34472, 17.34474, 17.34468, 
    17.34472, 17.34476, 17.34476, 17.34475, 17.34476, 17.34473, 17.34474, 
    17.34471, 17.34472, 17.34471, 17.34472, 17.34472, 17.34472, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34474, 17.34473, 17.34473, 17.34472, 17.34474, 
    17.34472, 17.34475, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 
    17.34475, 17.34474, 17.34473, 17.34472, 17.34471, 17.3447, 17.34469, 
    17.3447, 17.34468, 17.3447, 17.34467, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34473, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34468, 17.34467, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 TOTSOMC_1m =
  17.3448, 17.34479, 17.34479, 17.34478, 17.34479, 17.34478, 17.3448, 
    17.34479, 17.3448, 17.3448, 17.34476, 17.34478, 17.34474, 17.34475, 
    17.34472, 17.34474, 17.34472, 17.34472, 17.34471, 17.34471, 17.34469, 
    17.34471, 17.34468, 17.3447, 17.34469, 17.34471, 17.34478, 17.34476, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.34479, 17.3448, 17.3448, 
    17.3448, 17.34478, 17.34478, 17.34477, 17.34477, 17.34475, 17.34476, 
    17.34473, 17.34474, 17.34471, 17.34472, 17.34471, 17.34471, 17.34471, 
    17.34472, 17.34472, 17.34472, 17.34476, 17.34475, 17.34477, 17.34479, 
    17.3448, 17.34481, 17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 
    17.34477, 17.34477, 17.34475, 17.34474, 17.34472, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.34471, 17.34472, 17.34471, 17.34473, 
    17.34472, 17.34476, 17.34478, 17.34479, 17.34479, 17.34481, 17.3448, 
    17.3448, 17.34479, 17.34479, 17.34479, 17.34477, 17.34478, 17.34474, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34472, 17.34471, 17.34472, 
    17.34471, 17.3447, 17.3447, 17.34469, 17.34472, 17.34471, 17.34479, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.3448, 17.3448, 17.34479, 
    17.34479, 17.34478, 17.34478, 17.34477, 17.34476, 17.34474, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34472, 17.34473, 17.3447, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.34479, 17.3448, 
    17.34479, 17.3448, 17.3448, 17.34479, 17.34478, 17.34477, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34472, 17.3447, 17.3447, 
    17.3447, 17.3447, 17.34479, 17.34479, 17.34479, 17.34478, 17.34479, 
    17.34477, 17.34477, 17.34475, 17.34476, 17.34474, 17.34476, 17.34475, 
    17.34474, 17.34476, 17.34473, 17.34475, 17.34472, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.34469, 17.34469, 17.34468, 
    17.34478, 17.34477, 17.34477, 17.34477, 17.34476, 17.34475, 17.34474, 
    17.34474, 17.34473, 17.34473, 17.34475, 17.34474, 17.34477, 17.34476, 
    17.34477, 17.34478, 17.34474, 17.34476, 17.34473, 17.34474, 17.34471, 
    17.34472, 17.34469, 17.34468, 17.34467, 17.34466, 17.34477, 17.34477, 
    17.34477, 17.34476, 17.34475, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34472, 17.34473, 17.34472, 17.34476, 17.34474, 17.34478, 17.34476, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34472, 17.34473, 17.34468, 
    17.34471, 17.34465, 17.34466, 17.34478, 17.34477, 17.34475, 17.34476, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34471, 17.34472, 
    17.34471, 17.34474, 17.34473, 17.34475, 17.34475, 17.34475, 17.34475, 
    17.34474, 17.34473, 17.34473, 17.34473, 17.34472, 17.34474, 17.34468, 
    17.34472, 17.34476, 17.34476, 17.34475, 17.34476, 17.34473, 17.34474, 
    17.34471, 17.34472, 17.34471, 17.34472, 17.34472, 17.34472, 17.34473, 
    17.34474, 17.34475, 17.34476, 17.34476, 17.34475, 17.34473, 17.34472, 
    17.34472, 17.34471, 17.34474, 17.34473, 17.34473, 17.34472, 17.34474, 
    17.34472, 17.34475, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 
    17.34472, 17.34473, 17.34473, 17.34474, 17.34474, 17.34475, 17.34475, 
    17.34475, 17.34474, 17.34473, 17.34472, 17.34471, 17.3447, 17.34469, 
    17.3447, 17.34468, 17.3447, 17.34467, 17.34472, 17.3447, 17.34474, 
    17.34474, 17.34473, 17.34471, 17.34472, 17.34471, 17.34473, 17.34475, 
    17.34475, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 17.34473, 
    17.34474, 17.34472, 17.34471, 17.34468, 17.34467, 17.34466, 17.34465, 
    17.34465, 17.34465 ;

 TOTSOMN =
  1.773786, 1.773784, 1.773784, 1.773783, 1.773783, 1.773782, 1.773785, 
    1.773784, 1.773785, 1.773785, 1.77378, 1.773782, 1.773777, 1.773779, 
    1.773774, 1.773777, 1.773773, 1.773774, 1.773772, 1.773773, 1.77377, 
    1.773772, 1.773769, 1.77377, 1.77377, 1.773772, 1.773782, 1.77378, 
    1.773782, 1.773782, 1.773782, 1.773783, 1.773784, 1.773786, 1.773785, 
    1.773784, 1.773782, 1.773783, 1.77378, 1.77378, 1.773778, 1.773779, 
    1.773775, 1.773776, 1.773773, 1.773773, 1.773773, 1.773773, 1.773773, 
    1.773774, 1.773773, 1.773775, 1.773779, 1.773777, 1.773781, 1.773784, 
    1.773785, 1.773786, 1.773786, 1.773786, 1.773784, 1.773783, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773777, 1.773775, 1.773775, 1.773774, 
    1.773774, 1.773772, 1.773772, 1.773772, 1.773774, 1.773773, 1.773775, 
    1.773775, 1.77378, 1.773782, 1.773783, 1.773784, 1.773786, 1.773785, 
    1.773785, 1.773784, 1.773783, 1.773783, 1.773781, 1.773782, 1.773777, 
    1.773779, 1.773774, 1.773775, 1.773773, 1.773774, 1.773773, 1.773774, 
    1.773772, 1.773771, 1.773772, 1.77377, 1.773774, 1.773773, 1.773784, 
    1.773783, 1.773783, 1.773785, 1.773785, 1.773786, 1.773785, 1.773784, 
    1.773783, 1.773782, 1.773782, 1.77378, 1.773779, 1.773776, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773775, 1.773775, 1.773771, 1.773773, 
    1.77377, 1.773771, 1.773772, 1.773771, 1.773783, 1.773784, 1.773785, 
    1.773784, 1.773786, 1.773785, 1.773784, 1.773782, 1.773782, 1.773781, 
    1.77378, 1.773779, 1.773777, 1.773775, 1.773773, 1.773774, 1.773774, 
    1.773773, 1.773774, 1.773773, 1.773773, 1.773773, 1.773771, 1.773771, 
    1.773771, 1.773771, 1.773784, 1.773783, 1.773783, 1.773783, 1.773783, 
    1.773781, 1.773781, 1.773778, 1.773779, 1.773777, 1.773779, 1.773779, 
    1.773777, 1.773779, 1.773775, 1.773778, 1.773773, 1.773776, 1.773773, 
    1.773774, 1.773773, 1.773772, 1.773771, 1.77377, 1.77377, 1.773769, 
    1.773782, 1.773781, 1.773781, 1.773781, 1.77378, 1.773779, 1.773776, 
    1.773777, 1.773776, 1.773775, 1.773778, 1.773776, 1.773781, 1.77378, 
    1.77378, 1.773782, 1.773777, 1.77378, 1.773775, 1.773776, 1.773772, 
    1.773774, 1.77377, 1.773769, 1.773767, 1.773765, 1.773781, 1.773781, 
    1.77378, 1.773779, 1.773778, 1.773776, 1.773776, 1.773776, 1.773775, 
    1.773774, 1.773776, 1.773774, 1.77378, 1.773777, 1.773782, 1.77378, 
    1.773779, 1.77378, 1.773777, 1.773777, 1.773775, 1.773776, 1.773769, 
    1.773772, 1.773764, 1.773766, 1.773782, 1.773781, 1.773778, 1.77378, 
    1.773776, 1.773775, 1.773775, 1.773774, 1.773774, 1.773773, 1.773774, 
    1.773773, 1.773776, 1.773775, 1.773779, 1.773778, 1.773778, 1.773779, 
    1.773777, 1.773776, 1.773775, 1.773775, 1.773774, 1.773776, 1.773769, 
    1.773773, 1.77378, 1.773779, 1.773778, 1.773779, 1.773775, 1.773777, 
    1.773773, 1.773774, 1.773772, 1.773773, 1.773773, 1.773774, 1.773775, 
    1.773777, 1.773778, 1.773779, 1.773779, 1.773777, 1.773775, 1.773773, 
    1.773774, 1.773772, 1.773776, 1.773775, 1.773775, 1.773774, 1.773777, 
    1.773774, 1.773778, 1.773778, 1.773777, 1.773775, 1.773774, 1.773774, 
    1.773774, 1.773775, 1.773776, 1.773777, 1.773777, 1.773778, 1.773778, 
    1.773778, 1.773777, 1.773775, 1.773774, 1.773772, 1.773772, 1.77377, 
    1.773771, 1.773769, 1.773771, 1.773767, 1.773774, 1.773771, 1.773777, 
    1.773776, 1.773775, 1.773772, 1.773774, 1.773772, 1.773776, 1.773777, 
    1.773778, 1.773779, 1.773778, 1.773778, 1.773777, 1.773777, 1.773775, 
    1.773776, 1.773773, 1.773772, 1.773769, 1.773767, 1.773765, 1.773764, 
    1.773764, 1.773763 ;

 TOTSOMN_1m =
  1.773786, 1.773784, 1.773784, 1.773783, 1.773783, 1.773782, 1.773785, 
    1.773784, 1.773785, 1.773785, 1.77378, 1.773782, 1.773777, 1.773779, 
    1.773774, 1.773777, 1.773773, 1.773774, 1.773772, 1.773773, 1.77377, 
    1.773772, 1.773769, 1.77377, 1.77377, 1.773772, 1.773782, 1.77378, 
    1.773782, 1.773782, 1.773782, 1.773783, 1.773784, 1.773786, 1.773785, 
    1.773784, 1.773782, 1.773783, 1.77378, 1.77378, 1.773778, 1.773779, 
    1.773775, 1.773776, 1.773773, 1.773773, 1.773773, 1.773773, 1.773773, 
    1.773774, 1.773773, 1.773775, 1.773779, 1.773777, 1.773781, 1.773784, 
    1.773785, 1.773786, 1.773786, 1.773786, 1.773784, 1.773783, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773777, 1.773775, 1.773775, 1.773774, 
    1.773774, 1.773772, 1.773772, 1.773772, 1.773774, 1.773773, 1.773775, 
    1.773775, 1.77378, 1.773782, 1.773783, 1.773784, 1.773786, 1.773785, 
    1.773785, 1.773784, 1.773783, 1.773783, 1.773781, 1.773782, 1.773777, 
    1.773779, 1.773774, 1.773775, 1.773773, 1.773774, 1.773773, 1.773774, 
    1.773772, 1.773771, 1.773772, 1.77377, 1.773774, 1.773773, 1.773784, 
    1.773783, 1.773783, 1.773785, 1.773785, 1.773786, 1.773785, 1.773784, 
    1.773783, 1.773782, 1.773782, 1.77378, 1.773779, 1.773776, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773775, 1.773775, 1.773771, 1.773773, 
    1.77377, 1.773771, 1.773772, 1.773771, 1.773783, 1.773784, 1.773785, 
    1.773784, 1.773786, 1.773785, 1.773784, 1.773782, 1.773782, 1.773781, 
    1.77378, 1.773779, 1.773777, 1.773775, 1.773773, 1.773774, 1.773774, 
    1.773773, 1.773774, 1.773773, 1.773773, 1.773773, 1.773771, 1.773771, 
    1.773771, 1.773771, 1.773784, 1.773783, 1.773783, 1.773783, 1.773783, 
    1.773781, 1.773781, 1.773778, 1.773779, 1.773777, 1.773779, 1.773779, 
    1.773777, 1.773779, 1.773775, 1.773778, 1.773773, 1.773776, 1.773773, 
    1.773774, 1.773773, 1.773772, 1.773771, 1.77377, 1.77377, 1.773769, 
    1.773782, 1.773781, 1.773781, 1.773781, 1.77378, 1.773779, 1.773776, 
    1.773777, 1.773776, 1.773775, 1.773778, 1.773776, 1.773781, 1.77378, 
    1.77378, 1.773782, 1.773777, 1.77378, 1.773775, 1.773776, 1.773772, 
    1.773774, 1.77377, 1.773769, 1.773767, 1.773765, 1.773781, 1.773781, 
    1.77378, 1.773779, 1.773778, 1.773776, 1.773776, 1.773776, 1.773775, 
    1.773774, 1.773776, 1.773774, 1.77378, 1.773777, 1.773782, 1.77378, 
    1.773779, 1.77378, 1.773777, 1.773777, 1.773775, 1.773776, 1.773769, 
    1.773772, 1.773764, 1.773766, 1.773782, 1.773781, 1.773778, 1.77378, 
    1.773776, 1.773775, 1.773775, 1.773774, 1.773774, 1.773773, 1.773774, 
    1.773773, 1.773776, 1.773775, 1.773779, 1.773778, 1.773778, 1.773779, 
    1.773777, 1.773776, 1.773775, 1.773775, 1.773774, 1.773776, 1.773769, 
    1.773773, 1.77378, 1.773779, 1.773778, 1.773779, 1.773775, 1.773777, 
    1.773773, 1.773774, 1.773772, 1.773773, 1.773773, 1.773774, 1.773775, 
    1.773777, 1.773778, 1.773779, 1.773779, 1.773777, 1.773775, 1.773773, 
    1.773774, 1.773772, 1.773776, 1.773775, 1.773775, 1.773774, 1.773777, 
    1.773774, 1.773778, 1.773778, 1.773777, 1.773775, 1.773774, 1.773774, 
    1.773774, 1.773775, 1.773776, 1.773777, 1.773777, 1.773778, 1.773778, 
    1.773778, 1.773777, 1.773775, 1.773774, 1.773772, 1.773772, 1.77377, 
    1.773771, 1.773769, 1.773771, 1.773767, 1.773774, 1.773771, 1.773777, 
    1.773776, 1.773775, 1.773772, 1.773774, 1.773772, 1.773776, 1.773777, 
    1.773778, 1.773779, 1.773778, 1.773778, 1.773777, 1.773777, 1.773775, 
    1.773776, 1.773773, 1.773772, 1.773769, 1.773767, 1.773765, 1.773764, 
    1.773764, 1.773763 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9785, 249.9788, 249.9788, 249.979, 249.9789, 249.979, 249.9786, 
    249.9788, 249.9787, 249.9786, 249.9794, 249.979, 249.9799, 249.9796, 
    249.9803, 249.9798, 249.9804, 249.9803, 249.9806, 249.9805, 249.9809, 
    249.9806, 249.9811, 249.9808, 249.9809, 249.9806, 249.9791, 249.9794, 
    249.9791, 249.9791, 249.9791, 249.9789, 249.9787, 249.9785, 249.9786, 
    249.9787, 249.9791, 249.979, 249.9793, 249.9793, 249.9797, 249.9795, 
    249.9802, 249.98, 249.9805, 249.9804, 249.9805, 249.9805, 249.9805, 
    249.9803, 249.9804, 249.9802, 249.9796, 249.9798, 249.9792, 249.9788, 
    249.9786, 249.9785, 249.9785, 249.9785, 249.9787, 249.9789, 249.9791, 
    249.9792, 249.9793, 249.9796, 249.9798, 249.9802, 249.9801, 249.9802, 
    249.9804, 249.9805, 249.9805, 249.9806, 249.9802, 249.9805, 249.9801, 
    249.9802, 249.9793, 249.979, 249.9789, 249.9788, 249.9785, 249.9787, 
    249.9786, 249.9788, 249.9789, 249.9789, 249.9792, 249.9791, 249.9798, 
    249.9795, 249.9803, 249.9801, 249.9804, 249.9803, 249.9805, 249.9803, 
    249.9806, 249.9807, 249.9807, 249.9809, 249.9803, 249.9805, 249.9789, 
    249.9789, 249.9789, 249.9787, 249.9787, 249.9785, 249.9787, 249.9787, 
    249.9789, 249.979, 249.9791, 249.9793, 249.9796, 249.9799, 249.9802, 
    249.9803, 249.9802, 249.9803, 249.9802, 249.9802, 249.9807, 249.9804, 
    249.9808, 249.9808, 249.9806, 249.9808, 249.9789, 249.9788, 249.9786, 
    249.9788, 249.9785, 249.9787, 249.9787, 249.9791, 249.9792, 249.9792, 
    249.9794, 249.9795, 249.9798, 249.9801, 249.9804, 249.9803, 249.9804, 
    249.9804, 249.9803, 249.9804, 249.9805, 249.9804, 249.9808, 249.9807, 
    249.9808, 249.9807, 249.9788, 249.9789, 249.9789, 249.979, 249.9789, 
    249.9792, 249.9793, 249.9797, 249.9795, 249.9798, 249.9796, 249.9796, 
    249.9798, 249.9796, 249.9801, 249.9797, 249.9804, 249.98, 249.9804, 
    249.9804, 249.9805, 249.9806, 249.9807, 249.9809, 249.9809, 249.9811, 
    249.9791, 249.9792, 249.9792, 249.9793, 249.9794, 249.9796, 249.9799, 
    249.9798, 249.98, 249.9801, 249.9797, 249.9799, 249.9793, 249.9794, 
    249.9793, 249.9791, 249.9798, 249.9794, 249.9802, 249.9799, 249.9806, 
    249.9803, 249.9809, 249.9811, 249.9814, 249.9816, 249.9792, 249.9792, 
    249.9793, 249.9795, 249.9797, 249.98, 249.98, 249.98, 249.9802, 249.9803, 
    249.98, 249.9803, 249.9794, 249.9799, 249.9791, 249.9794, 249.9795, 
    249.9794, 249.9798, 249.9799, 249.9802, 249.98, 249.981, 249.9806, 
    249.9819, 249.9815, 249.9791, 249.9792, 249.9796, 249.9794, 249.98, 
    249.9801, 249.9802, 249.9803, 249.9804, 249.9804, 249.9803, 249.9804, 
    249.98, 249.9802, 249.9796, 249.9797, 249.9797, 249.9796, 249.9798, 
    249.9801, 249.9801, 249.9801, 249.9803, 249.98, 249.9811, 249.9804, 
    249.9794, 249.9796, 249.9796, 249.9795, 249.9801, 249.9799, 249.9804, 
    249.9803, 249.9805, 249.9804, 249.9804, 249.9802, 249.9801, 249.9799, 
    249.9797, 249.9796, 249.9796, 249.9798, 249.9801, 249.9804, 249.9803, 
    249.9805, 249.9799, 249.9802, 249.9801, 249.9803, 249.9798, 249.9802, 
    249.9797, 249.9797, 249.9799, 249.9802, 249.9803, 249.9803, 249.9803, 
    249.9801, 249.98, 249.9799, 249.9798, 249.9797, 249.9796, 249.9797, 
    249.9798, 249.9801, 249.9803, 249.9806, 249.9807, 249.9809, 249.9807, 
    249.9811, 249.9807, 249.9814, 249.9803, 249.9807, 249.9799, 249.98, 
    249.9801, 249.9805, 249.9803, 249.9806, 249.98, 249.9798, 249.9797, 
    249.9796, 249.9797, 249.9797, 249.9798, 249.9798, 249.9801, 249.9799, 
    249.9804, 249.9806, 249.9811, 249.9814, 249.9817, 249.9818, 249.9819, 
    249.9819 ;

 TREFMNAV_R =
  249.9785, 249.9788, 249.9788, 249.979, 249.9789, 249.979, 249.9786, 
    249.9788, 249.9787, 249.9786, 249.9794, 249.979, 249.9799, 249.9796, 
    249.9803, 249.9798, 249.9804, 249.9803, 249.9806, 249.9805, 249.9809, 
    249.9806, 249.9811, 249.9808, 249.9809, 249.9806, 249.9791, 249.9794, 
    249.9791, 249.9791, 249.9791, 249.9789, 249.9787, 249.9785, 249.9786, 
    249.9787, 249.9791, 249.979, 249.9793, 249.9793, 249.9797, 249.9795, 
    249.9802, 249.98, 249.9805, 249.9804, 249.9805, 249.9805, 249.9805, 
    249.9803, 249.9804, 249.9802, 249.9796, 249.9798, 249.9792, 249.9788, 
    249.9786, 249.9785, 249.9785, 249.9785, 249.9787, 249.9789, 249.9791, 
    249.9792, 249.9793, 249.9796, 249.9798, 249.9802, 249.9801, 249.9802, 
    249.9804, 249.9805, 249.9805, 249.9806, 249.9802, 249.9805, 249.9801, 
    249.9802, 249.9793, 249.979, 249.9789, 249.9788, 249.9785, 249.9787, 
    249.9786, 249.9788, 249.9789, 249.9789, 249.9792, 249.9791, 249.9798, 
    249.9795, 249.9803, 249.9801, 249.9804, 249.9803, 249.9805, 249.9803, 
    249.9806, 249.9807, 249.9807, 249.9809, 249.9803, 249.9805, 249.9789, 
    249.9789, 249.9789, 249.9787, 249.9787, 249.9785, 249.9787, 249.9787, 
    249.9789, 249.979, 249.9791, 249.9793, 249.9796, 249.9799, 249.9802, 
    249.9803, 249.9802, 249.9803, 249.9802, 249.9802, 249.9807, 249.9804, 
    249.9808, 249.9808, 249.9806, 249.9808, 249.9789, 249.9788, 249.9786, 
    249.9788, 249.9785, 249.9787, 249.9787, 249.9791, 249.9792, 249.9792, 
    249.9794, 249.9795, 249.9798, 249.9801, 249.9804, 249.9803, 249.9804, 
    249.9804, 249.9803, 249.9804, 249.9805, 249.9804, 249.9808, 249.9807, 
    249.9808, 249.9807, 249.9788, 249.9789, 249.9789, 249.979, 249.9789, 
    249.9792, 249.9793, 249.9797, 249.9795, 249.9798, 249.9796, 249.9796, 
    249.9798, 249.9796, 249.9801, 249.9797, 249.9804, 249.98, 249.9804, 
    249.9804, 249.9805, 249.9806, 249.9807, 249.9809, 249.9809, 249.9811, 
    249.9791, 249.9792, 249.9792, 249.9793, 249.9794, 249.9796, 249.9799, 
    249.9798, 249.98, 249.9801, 249.9797, 249.9799, 249.9793, 249.9794, 
    249.9793, 249.9791, 249.9798, 249.9794, 249.9802, 249.9799, 249.9806, 
    249.9803, 249.9809, 249.9811, 249.9814, 249.9816, 249.9792, 249.9792, 
    249.9793, 249.9795, 249.9797, 249.98, 249.98, 249.98, 249.9802, 249.9803, 
    249.98, 249.9803, 249.9794, 249.9799, 249.9791, 249.9794, 249.9795, 
    249.9794, 249.9798, 249.9799, 249.9802, 249.98, 249.981, 249.9806, 
    249.9819, 249.9815, 249.9791, 249.9792, 249.9796, 249.9794, 249.98, 
    249.9801, 249.9802, 249.9803, 249.9804, 249.9804, 249.9803, 249.9804, 
    249.98, 249.9802, 249.9796, 249.9797, 249.9797, 249.9796, 249.9798, 
    249.9801, 249.9801, 249.9801, 249.9803, 249.98, 249.9811, 249.9804, 
    249.9794, 249.9796, 249.9796, 249.9795, 249.9801, 249.9799, 249.9804, 
    249.9803, 249.9805, 249.9804, 249.9804, 249.9802, 249.9801, 249.9799, 
    249.9797, 249.9796, 249.9796, 249.9798, 249.9801, 249.9804, 249.9803, 
    249.9805, 249.9799, 249.9802, 249.9801, 249.9803, 249.9798, 249.9802, 
    249.9797, 249.9797, 249.9799, 249.9802, 249.9803, 249.9803, 249.9803, 
    249.9801, 249.98, 249.9799, 249.9798, 249.9797, 249.9796, 249.9797, 
    249.9798, 249.9801, 249.9803, 249.9806, 249.9807, 249.9809, 249.9807, 
    249.9811, 249.9807, 249.9814, 249.9803, 249.9807, 249.9799, 249.98, 
    249.9801, 249.9805, 249.9803, 249.9806, 249.98, 249.9798, 249.9797, 
    249.9796, 249.9797, 249.9797, 249.9798, 249.9798, 249.9801, 249.9799, 
    249.9804, 249.9806, 249.9811, 249.9814, 249.9817, 249.9818, 249.9819, 
    249.9819 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.6035, 258.6039, 258.6038, 258.6041, 258.6039, 258.6041, 258.6036, 
    258.6039, 258.6037, 258.6036, 258.6046, 258.6041, 258.6052, 258.6049, 
    258.6057, 258.6051, 258.6058, 258.6057, 258.6061, 258.606, 258.6064, 
    258.6061, 258.6067, 258.6064, 258.6064, 258.6061, 258.6042, 258.6046, 
    258.6042, 258.6042, 258.6042, 258.6039, 258.6038, 258.6035, 258.6036, 
    258.6038, 258.6043, 258.6041, 258.6045, 258.6045, 258.605, 258.6048, 
    258.6055, 258.6053, 258.606, 258.6058, 258.606, 258.6059, 258.606, 
    258.6057, 258.6058, 258.6056, 258.6048, 258.605, 258.6043, 258.6039, 
    258.6036, 258.6034, 258.6035, 258.6035, 258.6038, 258.604, 258.6042, 
    258.6044, 258.6045, 258.6049, 258.6051, 258.6056, 258.6055, 258.6057, 
    258.6058, 258.606, 258.606, 258.6061, 258.6057, 258.6059, 258.6055, 
    258.6056, 258.6045, 258.6042, 258.604, 258.6038, 258.6035, 258.6037, 
    258.6036, 258.6039, 258.604, 258.6039, 258.6044, 258.6042, 258.6051, 
    258.6047, 258.6058, 258.6055, 258.6058, 258.6057, 258.6059, 258.6057, 
    258.6061, 258.6062, 258.6061, 258.6064, 258.6057, 258.606, 258.6039, 
    258.6039, 258.604, 258.6038, 258.6037, 258.6035, 258.6037, 258.6038, 
    258.604, 258.6042, 258.6042, 258.6045, 258.6048, 258.6052, 258.6055, 
    258.6057, 258.6056, 258.6057, 258.6056, 258.6056, 258.6062, 258.6058, 
    258.6064, 258.6063, 258.6061, 258.6063, 258.6039, 258.6039, 258.6036, 
    258.6038, 258.6035, 258.6037, 258.6038, 258.6042, 258.6043, 258.6044, 
    258.6046, 258.6048, 258.6052, 258.6055, 258.6058, 258.6058, 258.6058, 
    258.6058, 258.6057, 258.6059, 258.6059, 258.6058, 258.6063, 258.6062, 
    258.6063, 258.6062, 258.6039, 258.604, 258.604, 258.6041, 258.604, 
    258.6043, 258.6045, 258.605, 258.6048, 258.6051, 258.6048, 258.6049, 
    258.6051, 258.6048, 258.6055, 258.605, 258.6059, 258.6054, 258.6059, 
    258.6058, 258.6059, 258.606, 258.6062, 258.6065, 258.6064, 258.6067, 
    258.6042, 258.6043, 258.6043, 258.6045, 258.6046, 258.6049, 258.6053, 
    258.6051, 258.6054, 258.6054, 258.605, 258.6053, 258.6044, 258.6046, 
    258.6045, 258.6042, 258.6051, 258.6046, 258.6055, 258.6053, 258.606, 
    258.6057, 258.6064, 258.6067, 258.607, 258.6074, 258.6044, 258.6043, 
    258.6045, 258.6047, 258.605, 258.6053, 258.6053, 258.6054, 258.6055, 
    258.6057, 258.6054, 258.6057, 258.6046, 258.6052, 258.6043, 258.6046, 
    258.6047, 258.6046, 258.6051, 258.6052, 258.6056, 258.6054, 258.6066, 
    258.6061, 258.6076, 258.6072, 258.6043, 258.6044, 258.6049, 258.6047, 
    258.6053, 258.6055, 258.6056, 258.6058, 258.6058, 258.6059, 258.6057, 
    258.6059, 258.6053, 258.6056, 258.6049, 258.605, 258.6049, 258.6049, 
    258.6051, 258.6054, 258.6054, 258.6055, 258.6057, 258.6053, 258.6067, 
    258.6058, 258.6046, 258.6048, 258.6049, 258.6048, 258.6055, 258.6052, 
    258.6059, 258.6057, 258.606, 258.6059, 258.6058, 258.6057, 258.6055, 
    258.6052, 258.605, 258.6048, 258.6048, 258.605, 258.6054, 258.6058, 
    258.6057, 258.606, 258.6053, 258.6056, 258.6054, 258.6057, 258.6051, 
    258.6057, 258.6049, 258.605, 258.6052, 258.6056, 258.6057, 258.6058, 
    258.6057, 258.6054, 258.6054, 258.6052, 258.6051, 258.605, 258.6049, 
    258.605, 258.6051, 258.6054, 258.6057, 258.606, 258.6061, 258.6065, 
    258.6062, 258.6067, 258.6063, 258.607, 258.6057, 258.6063, 258.6052, 
    258.6053, 258.6055, 258.606, 258.6057, 258.606, 258.6054, 258.605, 
    258.6049, 258.6048, 258.605, 258.6049, 258.6051, 258.6051, 258.6054, 
    258.6053, 258.6058, 258.606, 258.6067, 258.607, 258.6074, 258.6076, 
    258.6077, 258.6077 ;

 TREFMXAV_R =
  258.6035, 258.6039, 258.6038, 258.6041, 258.6039, 258.6041, 258.6036, 
    258.6039, 258.6037, 258.6036, 258.6046, 258.6041, 258.6052, 258.6049, 
    258.6057, 258.6051, 258.6058, 258.6057, 258.6061, 258.606, 258.6064, 
    258.6061, 258.6067, 258.6064, 258.6064, 258.6061, 258.6042, 258.6046, 
    258.6042, 258.6042, 258.6042, 258.6039, 258.6038, 258.6035, 258.6036, 
    258.6038, 258.6043, 258.6041, 258.6045, 258.6045, 258.605, 258.6048, 
    258.6055, 258.6053, 258.606, 258.6058, 258.606, 258.6059, 258.606, 
    258.6057, 258.6058, 258.6056, 258.6048, 258.605, 258.6043, 258.6039, 
    258.6036, 258.6034, 258.6035, 258.6035, 258.6038, 258.604, 258.6042, 
    258.6044, 258.6045, 258.6049, 258.6051, 258.6056, 258.6055, 258.6057, 
    258.6058, 258.606, 258.606, 258.6061, 258.6057, 258.6059, 258.6055, 
    258.6056, 258.6045, 258.6042, 258.604, 258.6038, 258.6035, 258.6037, 
    258.6036, 258.6039, 258.604, 258.6039, 258.6044, 258.6042, 258.6051, 
    258.6047, 258.6058, 258.6055, 258.6058, 258.6057, 258.6059, 258.6057, 
    258.6061, 258.6062, 258.6061, 258.6064, 258.6057, 258.606, 258.6039, 
    258.6039, 258.604, 258.6038, 258.6037, 258.6035, 258.6037, 258.6038, 
    258.604, 258.6042, 258.6042, 258.6045, 258.6048, 258.6052, 258.6055, 
    258.6057, 258.6056, 258.6057, 258.6056, 258.6056, 258.6062, 258.6058, 
    258.6064, 258.6063, 258.6061, 258.6063, 258.6039, 258.6039, 258.6036, 
    258.6038, 258.6035, 258.6037, 258.6038, 258.6042, 258.6043, 258.6044, 
    258.6046, 258.6048, 258.6052, 258.6055, 258.6058, 258.6058, 258.6058, 
    258.6058, 258.6057, 258.6059, 258.6059, 258.6058, 258.6063, 258.6062, 
    258.6063, 258.6062, 258.6039, 258.604, 258.604, 258.6041, 258.604, 
    258.6043, 258.6045, 258.605, 258.6048, 258.6051, 258.6048, 258.6049, 
    258.6051, 258.6048, 258.6055, 258.605, 258.6059, 258.6054, 258.6059, 
    258.6058, 258.6059, 258.606, 258.6062, 258.6065, 258.6064, 258.6067, 
    258.6042, 258.6043, 258.6043, 258.6045, 258.6046, 258.6049, 258.6053, 
    258.6051, 258.6054, 258.6054, 258.605, 258.6053, 258.6044, 258.6046, 
    258.6045, 258.6042, 258.6051, 258.6046, 258.6055, 258.6053, 258.606, 
    258.6057, 258.6064, 258.6067, 258.607, 258.6074, 258.6044, 258.6043, 
    258.6045, 258.6047, 258.605, 258.6053, 258.6053, 258.6054, 258.6055, 
    258.6057, 258.6054, 258.6057, 258.6046, 258.6052, 258.6043, 258.6046, 
    258.6047, 258.6046, 258.6051, 258.6052, 258.6056, 258.6054, 258.6066, 
    258.6061, 258.6076, 258.6072, 258.6043, 258.6044, 258.6049, 258.6047, 
    258.6053, 258.6055, 258.6056, 258.6058, 258.6058, 258.6059, 258.6057, 
    258.6059, 258.6053, 258.6056, 258.6049, 258.605, 258.6049, 258.6049, 
    258.6051, 258.6054, 258.6054, 258.6055, 258.6057, 258.6053, 258.6067, 
    258.6058, 258.6046, 258.6048, 258.6049, 258.6048, 258.6055, 258.6052, 
    258.6059, 258.6057, 258.606, 258.6059, 258.6058, 258.6057, 258.6055, 
    258.6052, 258.605, 258.6048, 258.6048, 258.605, 258.6054, 258.6058, 
    258.6057, 258.606, 258.6053, 258.6056, 258.6054, 258.6057, 258.6051, 
    258.6057, 258.6049, 258.605, 258.6052, 258.6056, 258.6057, 258.6058, 
    258.6057, 258.6054, 258.6054, 258.6052, 258.6051, 258.605, 258.6049, 
    258.605, 258.6051, 258.6054, 258.6057, 258.606, 258.6061, 258.6065, 
    258.6062, 258.6067, 258.6063, 258.607, 258.6057, 258.6063, 258.6052, 
    258.6053, 258.6055, 258.606, 258.6057, 258.606, 258.6054, 258.605, 
    258.6049, 258.6048, 258.605, 258.6049, 258.6051, 258.6051, 258.6054, 
    258.6053, 258.6058, 258.606, 258.6067, 258.607, 258.6074, 258.6076, 
    258.6077, 258.6077 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9705, 253.9706, 253.9706, 253.9708, 253.9707, 253.9708, 253.9705, 
    253.9707, 253.9706, 253.9705, 253.971, 253.9708, 253.9713, 253.9712, 
    253.9716, 253.9713, 253.9717, 253.9716, 253.9718, 253.9718, 253.972, 
    253.9718, 253.9722, 253.972, 253.972, 253.9718, 253.9708, 253.971, 
    253.9708, 253.9708, 253.9708, 253.9707, 253.9706, 253.9705, 253.9705, 
    253.9706, 253.9709, 253.9708, 253.971, 253.971, 253.9712, 253.9711, 
    253.9715, 253.9714, 253.9718, 253.9717, 253.9717, 253.9717, 253.9717, 
    253.9716, 253.9717, 253.9716, 253.9711, 253.9713, 253.9709, 253.9707, 
    253.9705, 253.9704, 253.9704, 253.9704, 253.9706, 253.9707, 253.9708, 
    253.9709, 253.971, 253.9712, 253.9713, 253.9716, 253.9715, 253.9716, 
    253.9717, 253.9718, 253.9718, 253.9718, 253.9716, 253.9717, 253.9715, 
    253.9716, 253.971, 253.9708, 253.9707, 253.9706, 253.9704, 253.9706, 
    253.9705, 253.9706, 253.9707, 253.9707, 253.9709, 253.9708, 253.9713, 
    253.9711, 253.9716, 253.9715, 253.9717, 253.9716, 253.9717, 253.9716, 
    253.9718, 253.9719, 253.9718, 253.972, 253.9716, 253.9717, 253.9707, 
    253.9707, 253.9707, 253.9706, 253.9706, 253.9705, 253.9706, 253.9706, 
    253.9707, 253.9708, 253.9708, 253.971, 253.9711, 253.9714, 253.9715, 
    253.9716, 253.9716, 253.9716, 253.9716, 253.9715, 253.9719, 253.9717, 
    253.972, 253.9719, 253.9718, 253.972, 253.9707, 253.9706, 253.9705, 
    253.9706, 253.9704, 253.9705, 253.9706, 253.9708, 253.9709, 253.9709, 
    253.971, 253.9711, 253.9713, 253.9715, 253.9717, 253.9716, 253.9716, 
    253.9717, 253.9716, 253.9717, 253.9717, 253.9717, 253.9719, 253.9719, 
    253.9719, 253.9719, 253.9707, 253.9707, 253.9707, 253.9707, 253.9707, 
    253.9709, 253.9709, 253.9712, 253.9711, 253.9713, 253.9711, 253.9712, 
    253.9713, 253.9711, 253.9715, 253.9713, 253.9717, 253.9715, 253.9717, 
    253.9717, 253.9717, 253.9718, 253.9719, 253.972, 253.972, 253.9721, 
    253.9708, 253.9709, 253.9709, 253.971, 253.971, 253.9712, 253.9714, 
    253.9713, 253.9714, 253.9715, 253.9713, 253.9714, 253.9709, 253.971, 
    253.971, 253.9708, 253.9713, 253.9711, 253.9715, 253.9714, 253.9718, 
    253.9716, 253.972, 253.9722, 253.9723, 253.9725, 253.9709, 253.9709, 
    253.971, 253.9711, 253.9712, 253.9714, 253.9714, 253.9715, 253.9715, 
    253.9716, 253.9715, 253.9716, 253.971, 253.9713, 253.9709, 253.971, 
    253.9711, 253.9711, 253.9713, 253.9713, 253.9716, 253.9715, 253.9721, 
    253.9718, 253.9726, 253.9724, 253.9709, 253.9709, 253.9712, 253.9711, 
    253.9714, 253.9715, 253.9716, 253.9716, 253.9717, 253.9717, 253.9716, 
    253.9717, 253.9714, 253.9715, 253.9712, 253.9713, 253.9712, 253.9712, 
    253.9713, 253.9715, 253.9715, 253.9715, 253.9716, 253.9714, 253.9721, 
    253.9717, 253.971, 253.9711, 253.9712, 253.9711, 253.9715, 253.9713, 
    253.9717, 253.9716, 253.9718, 253.9717, 253.9717, 253.9716, 253.9715, 
    253.9714, 253.9712, 253.9711, 253.9711, 253.9713, 253.9715, 253.9717, 
    253.9716, 253.9718, 253.9714, 253.9715, 253.9715, 253.9716, 253.9713, 
    253.9716, 253.9712, 253.9713, 253.9713, 253.9715, 253.9716, 253.9716, 
    253.9716, 253.9715, 253.9715, 253.9713, 253.9713, 253.9712, 253.9712, 
    253.9712, 253.9713, 253.9715, 253.9716, 253.9718, 253.9718, 253.972, 
    253.9719, 253.9721, 253.9719, 253.9723, 253.9716, 253.9719, 253.9714, 
    253.9714, 253.9715, 253.9718, 253.9716, 253.9718, 253.9715, 253.9713, 
    253.9712, 253.9711, 253.9712, 253.9712, 253.9713, 253.9713, 253.9715, 
    253.9714, 253.9717, 253.9718, 253.9721, 253.9723, 253.9725, 253.9726, 
    253.9727, 253.9727 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9705, 253.9706, 253.9706, 253.9708, 253.9707, 253.9708, 253.9705, 
    253.9707, 253.9706, 253.9705, 253.971, 253.9708, 253.9713, 253.9712, 
    253.9716, 253.9713, 253.9717, 253.9716, 253.9718, 253.9718, 253.972, 
    253.9718, 253.9722, 253.972, 253.972, 253.9718, 253.9708, 253.971, 
    253.9708, 253.9708, 253.9708, 253.9707, 253.9706, 253.9705, 253.9705, 
    253.9706, 253.9709, 253.9708, 253.971, 253.971, 253.9712, 253.9711, 
    253.9715, 253.9714, 253.9718, 253.9717, 253.9717, 253.9717, 253.9717, 
    253.9716, 253.9717, 253.9716, 253.9711, 253.9713, 253.9709, 253.9707, 
    253.9705, 253.9704, 253.9704, 253.9704, 253.9706, 253.9707, 253.9708, 
    253.9709, 253.971, 253.9712, 253.9713, 253.9716, 253.9715, 253.9716, 
    253.9717, 253.9718, 253.9718, 253.9718, 253.9716, 253.9717, 253.9715, 
    253.9716, 253.971, 253.9708, 253.9707, 253.9706, 253.9704, 253.9706, 
    253.9705, 253.9706, 253.9707, 253.9707, 253.9709, 253.9708, 253.9713, 
    253.9711, 253.9716, 253.9715, 253.9717, 253.9716, 253.9717, 253.9716, 
    253.9718, 253.9719, 253.9718, 253.972, 253.9716, 253.9717, 253.9707, 
    253.9707, 253.9707, 253.9706, 253.9706, 253.9705, 253.9706, 253.9706, 
    253.9707, 253.9708, 253.9708, 253.971, 253.9711, 253.9714, 253.9715, 
    253.9716, 253.9716, 253.9716, 253.9716, 253.9715, 253.9719, 253.9717, 
    253.972, 253.9719, 253.9718, 253.972, 253.9707, 253.9706, 253.9705, 
    253.9706, 253.9704, 253.9705, 253.9706, 253.9708, 253.9709, 253.9709, 
    253.971, 253.9711, 253.9713, 253.9715, 253.9717, 253.9716, 253.9716, 
    253.9717, 253.9716, 253.9717, 253.9717, 253.9717, 253.9719, 253.9719, 
    253.9719, 253.9719, 253.9707, 253.9707, 253.9707, 253.9707, 253.9707, 
    253.9709, 253.9709, 253.9712, 253.9711, 253.9713, 253.9711, 253.9712, 
    253.9713, 253.9711, 253.9715, 253.9713, 253.9717, 253.9715, 253.9717, 
    253.9717, 253.9717, 253.9718, 253.9719, 253.972, 253.972, 253.9721, 
    253.9708, 253.9709, 253.9709, 253.971, 253.971, 253.9712, 253.9714, 
    253.9713, 253.9714, 253.9715, 253.9713, 253.9714, 253.9709, 253.971, 
    253.971, 253.9708, 253.9713, 253.9711, 253.9715, 253.9714, 253.9718, 
    253.9716, 253.972, 253.9722, 253.9723, 253.9725, 253.9709, 253.9709, 
    253.971, 253.9711, 253.9712, 253.9714, 253.9714, 253.9715, 253.9715, 
    253.9716, 253.9715, 253.9716, 253.971, 253.9713, 253.9709, 253.971, 
    253.9711, 253.9711, 253.9713, 253.9713, 253.9716, 253.9715, 253.9721, 
    253.9718, 253.9726, 253.9724, 253.9709, 253.9709, 253.9712, 253.9711, 
    253.9714, 253.9715, 253.9716, 253.9716, 253.9717, 253.9717, 253.9716, 
    253.9717, 253.9714, 253.9715, 253.9712, 253.9713, 253.9712, 253.9712, 
    253.9713, 253.9715, 253.9715, 253.9715, 253.9716, 253.9714, 253.9721, 
    253.9717, 253.971, 253.9711, 253.9712, 253.9711, 253.9715, 253.9713, 
    253.9717, 253.9716, 253.9718, 253.9717, 253.9717, 253.9716, 253.9715, 
    253.9714, 253.9712, 253.9711, 253.9711, 253.9713, 253.9715, 253.9717, 
    253.9716, 253.9718, 253.9714, 253.9715, 253.9715, 253.9716, 253.9713, 
    253.9716, 253.9712, 253.9713, 253.9713, 253.9715, 253.9716, 253.9716, 
    253.9716, 253.9715, 253.9715, 253.9713, 253.9713, 253.9712, 253.9712, 
    253.9712, 253.9713, 253.9715, 253.9716, 253.9718, 253.9718, 253.972, 
    253.9719, 253.9721, 253.9719, 253.9723, 253.9716, 253.9719, 253.9714, 
    253.9714, 253.9715, 253.9718, 253.9716, 253.9718, 253.9715, 253.9713, 
    253.9712, 253.9711, 253.9712, 253.9712, 253.9713, 253.9713, 253.9715, 
    253.9714, 253.9717, 253.9718, 253.9721, 253.9723, 253.9725, 253.9726, 
    253.9727, 253.9727 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.4901, 254.4918, 254.4915, 254.4928, 254.4921, 254.493, 254.4905, 
    254.4919, 254.491, 254.4903, 254.4954, 254.4929, 254.4982, 254.4965, 
    254.5007, 254.4979, 254.5012, 254.5006, 254.5026, 254.502, 254.5044, 
    254.5028, 254.5057, 254.5041, 254.5043, 254.5027, 254.4934, 254.4951, 
    254.4933, 254.4936, 254.4935, 254.4921, 254.4914, 254.49, 254.4903, 
    254.4913, 254.4937, 254.4929, 254.4949, 254.4949, 254.4971, 254.4961, 
    254.5, 254.4989, 254.502, 254.5012, 254.502, 254.5018, 254.502, 254.5008, 
    254.5013, 254.5003, 254.4963, 254.4975, 254.494, 254.4919, 254.4906, 
    254.4896, 254.4897, 254.49, 254.4913, 254.4926, 254.4936, 254.4942, 
    254.4949, 254.4967, 254.4978, 254.5002, 254.4998, 254.5004, 254.5011, 
    254.5023, 254.5021, 254.5026, 254.5004, 254.5019, 254.4995, 254.5002, 
    254.4949, 254.4931, 254.4922, 254.4916, 254.4898, 254.491, 254.4905, 
    254.4917, 254.4924, 254.4921, 254.4942, 254.4934, 254.4979, 254.4959, 
    254.5011, 254.4998, 254.5014, 254.5006, 254.5019, 254.5007, 254.5028, 
    254.5032, 254.5029, 254.5041, 254.5007, 254.502, 254.492, 254.4921, 
    254.4924, 254.4912, 254.4911, 254.49, 254.491, 254.4914, 254.4924, 
    254.4931, 254.4937, 254.4949, 254.4964, 254.4984, 254.4999, 254.5009, 
    254.5003, 254.5008, 254.5002, 254.5, 254.5031, 254.5013, 254.504, 
    254.5038, 254.5026, 254.5038, 254.4921, 254.4918, 254.4906, 254.4916, 
    254.4899, 254.4908, 254.4913, 254.4934, 254.4939, 254.4943, 254.4951, 
    254.4962, 254.498, 254.4997, 254.5012, 254.5011, 254.5011, 254.5014, 
    254.5006, 254.5016, 254.5017, 254.5013, 254.5038, 254.5031, 254.5038, 
    254.5034, 254.4919, 254.4925, 254.4922, 254.4927, 254.4923, 254.4941, 
    254.4946, 254.4972, 254.4962, 254.4978, 254.4963, 254.4966, 254.4978, 
    254.4964, 254.4996, 254.4974, 254.5015, 254.4992, 254.5016, 254.5012, 
    254.5019, 254.5025, 254.5033, 254.5047, 254.5044, 254.5056, 254.4933, 
    254.494, 254.494, 254.4948, 254.4953, 254.4965, 254.4985, 254.4978, 
    254.4991, 254.4994, 254.4973, 254.4986, 254.4945, 254.4952, 254.4948, 
    254.4934, 254.4979, 254.4956, 254.4999, 254.4987, 254.5024, 254.5005, 
    254.5042, 254.5057, 254.5073, 254.509, 254.4944, 254.494, 254.4948, 
    254.496, 254.4972, 254.4987, 254.4989, 254.4992, 254.4999, 254.5006, 
    254.4993, 254.5007, 254.4953, 254.4981, 254.4937, 254.495, 254.496, 
    254.4956, 254.4977, 254.4982, 254.5002, 254.4992, 254.5053, 254.5026, 
    254.5103, 254.5081, 254.4938, 254.4944, 254.4967, 254.4957, 254.4989, 
    254.4996, 254.5003, 254.5011, 254.5012, 254.5017, 254.5009, 254.5016, 
    254.4987, 254.5, 254.4965, 254.4974, 254.497, 254.4965, 254.4979, 
    254.4993, 254.4993, 254.4998, 254.501, 254.4989, 254.5056, 254.5014, 
    254.4952, 254.4964, 254.4966, 254.4962, 254.4995, 254.4983, 254.5016, 
    254.5007, 254.5022, 254.5015, 254.5014, 254.5004, 254.4998, 254.4984, 
    254.4972, 254.4962, 254.4964, 254.4975, 254.4994, 254.5012, 254.5008, 
    254.5021, 254.4986, 254.5001, 254.4995, 254.501, 254.4978, 254.5004, 
    254.4971, 254.4974, 254.4983, 254.5002, 254.5006, 254.501, 254.5008, 
    254.4994, 254.4992, 254.4983, 254.498, 254.4973, 254.4967, 254.4972, 
    254.4978, 254.4994, 254.5009, 254.5025, 254.5029, 254.5047, 254.5032, 
    254.5056, 254.5035, 254.5073, 254.5006, 254.5035, 254.4983, 254.4989, 
    254.4999, 254.5022, 254.501, 254.5024, 254.4992, 254.4975, 254.4971, 
    254.4963, 254.4971, 254.497, 254.4978, 254.4976, 254.4995, 254.4985, 
    254.5014, 254.5024, 254.5055, 254.5073, 254.5092, 254.5101, 254.5103, 
    254.5105,
  255.5812, 255.5831, 255.5827, 255.5842, 255.5834, 255.5844, 255.5816, 
    255.5831, 255.5821, 255.5814, 255.5871, 255.5843, 255.5902, 255.5883, 
    255.593, 255.5899, 255.5936, 255.5929, 255.5951, 255.5945, 255.5972, 
    255.5954, 255.5987, 255.5968, 255.5971, 255.5954, 255.5849, 255.5867, 
    255.5848, 255.585, 255.5849, 255.5834, 255.5826, 255.5811, 255.5813, 
    255.5825, 255.5851, 255.5843, 255.5865, 255.5865, 255.589, 255.5879, 
    255.5922, 255.591, 255.5945, 255.5936, 255.5945, 255.5942, 255.5945, 
    255.5932, 255.5937, 255.5926, 255.5881, 255.5894, 255.5855, 255.5831, 
    255.5816, 255.5806, 255.5807, 255.581, 255.5825, 255.5839, 255.585, 
    255.5858, 255.5865, 255.5886, 255.5898, 255.5924, 255.592, 255.5928, 
    255.5935, 255.5948, 255.5946, 255.5952, 255.5928, 255.5943, 255.5917, 
    255.5924, 255.5866, 255.5845, 255.5835, 255.5828, 255.5808, 255.5822, 
    255.5816, 255.5829, 255.5837, 255.5833, 255.5858, 255.5848, 255.5899, 
    255.5877, 255.5934, 255.5921, 255.5938, 255.5929, 255.5944, 255.5931, 
    255.5954, 255.5959, 255.5956, 255.5969, 255.593, 255.5945, 255.5833, 
    255.5834, 255.5837, 255.5823, 255.5822, 255.581, 255.5821, 255.5826, 
    255.5838, 255.5845, 255.5851, 255.5866, 255.5882, 255.5905, 255.5921, 
    255.5933, 255.5926, 255.5932, 255.5925, 255.5922, 255.5957, 255.5937, 
    255.5967, 255.5965, 255.5952, 255.5966, 255.5834, 255.5831, 255.5817, 
    255.5828, 255.5809, 255.5819, 255.5825, 255.5848, 255.5854, 255.5858, 
    255.5867, 255.588, 255.59, 255.5919, 255.5936, 255.5935, 255.5935, 
    255.5939, 255.5929, 255.594, 255.5942, 255.5937, 255.5965, 255.5957, 
    255.5965, 255.596, 255.5832, 255.5838, 255.5835, 255.5841, 255.5836, 
    255.5856, 255.5862, 255.5891, 255.5879, 255.5898, 255.5881, 255.5884, 
    255.5898, 255.5882, 255.5918, 255.5893, 255.5939, 255.5914, 255.594, 
    255.5936, 255.5944, 255.595, 255.5959, 255.5976, 255.5972, 255.5986, 
    255.5847, 255.5855, 255.5855, 255.5863, 255.587, 255.5884, 255.5906, 
    255.5898, 255.5913, 255.5916, 255.5893, 255.5907, 255.5861, 255.5868, 
    255.5864, 255.5848, 255.5899, 255.5873, 255.5922, 255.5907, 255.595, 
    255.5928, 255.597, 255.5987, 255.6004, 255.6024, 255.586, 255.5854, 
    255.5865, 255.5878, 255.5891, 255.5908, 255.591, 255.5913, 255.5922, 
    255.5929, 255.5914, 255.593, 255.5869, 255.5901, 255.5852, 255.5867, 
    255.5877, 255.5873, 255.5897, 255.5902, 255.5925, 255.5913, 255.5983, 
    255.5952, 255.6039, 255.6014, 255.5853, 255.586, 255.5886, 255.5874, 
    255.591, 255.5918, 255.5926, 255.5935, 255.5936, 255.5941, 255.5932, 
    255.5941, 255.5908, 255.5923, 255.5883, 255.5893, 255.5888, 255.5884, 
    255.5899, 255.5914, 255.5915, 255.592, 255.5934, 255.591, 255.5986, 
    255.5938, 255.5868, 255.5882, 255.5885, 255.5879, 255.5917, 255.5903, 
    255.5941, 255.5931, 255.5948, 255.5939, 255.5938, 255.5927, 255.5921, 
    255.5904, 255.5891, 255.588, 255.5883, 255.5894, 255.5915, 255.5936, 
    255.5931, 255.5946, 255.5907, 255.5923, 255.5917, 255.5934, 255.5897, 
    255.5927, 255.5889, 255.5893, 255.5903, 255.5924, 255.5929, 255.5934, 
    255.5931, 255.5916, 255.5914, 255.5903, 255.59, 255.5892, 255.5885, 
    255.5891, 255.5898, 255.5916, 255.5932, 255.5951, 255.5955, 255.5976, 
    255.5959, 255.5986, 255.5962, 255.6004, 255.593, 255.5962, 255.5904, 
    255.591, 255.5921, 255.5947, 255.5934, 255.595, 255.5914, 255.5894, 
    255.589, 255.5881, 255.589, 255.5889, 255.5898, 255.5895, 255.5917, 
    255.5905, 255.5938, 255.595, 255.5984, 255.6005, 255.6027, 255.6036, 
    255.6039, 255.604,
  257.1418, 257.1438, 257.1434, 257.145, 257.1441, 257.1452, 257.1422, 
    257.1439, 257.1428, 257.142, 257.1481, 257.1451, 257.1514, 257.1494, 
    257.1545, 257.1511, 257.1552, 257.1544, 257.1568, 257.1561, 257.1591, 
    257.1571, 257.1606, 257.1586, 257.1589, 257.157, 257.1457, 257.1477, 
    257.1456, 257.1459, 257.1458, 257.1441, 257.1433, 257.1416, 257.1419, 
    257.1432, 257.146, 257.1451, 257.1475, 257.1475, 257.1502, 257.149, 
    257.1536, 257.1523, 257.1561, 257.1552, 257.1561, 257.1558, 257.1561, 
    257.1547, 257.1552, 257.154, 257.1492, 257.1506, 257.1464, 257.1439, 
    257.1422, 257.1411, 257.1412, 257.1416, 257.1432, 257.1447, 257.1459, 
    257.1467, 257.1475, 257.1497, 257.151, 257.1538, 257.1534, 257.1542, 
    257.1551, 257.1564, 257.1562, 257.1568, 257.1542, 257.1559, 257.1531, 
    257.1538, 257.1476, 257.1453, 257.1443, 257.1435, 257.1414, 257.1428, 
    257.1422, 257.1436, 257.1445, 257.144, 257.1467, 257.1457, 257.1511, 
    257.1487, 257.1549, 257.1535, 257.1553, 257.1544, 257.156, 257.1545, 
    257.157, 257.1576, 257.1572, 257.1587, 257.1544, 257.1561, 257.144, 
    257.1441, 257.1444, 257.143, 257.1429, 257.1416, 257.1428, 257.1432, 
    257.1445, 257.1453, 257.146, 257.1476, 257.1493, 257.1518, 257.1536, 
    257.1548, 257.154, 257.1547, 257.154, 257.1536, 257.1574, 257.1552, 
    257.1585, 257.1583, 257.1568, 257.1583, 257.1442, 257.1438, 257.1424, 
    257.1435, 257.1415, 257.1426, 257.1432, 257.1457, 257.1462, 257.1467, 
    257.1477, 257.149, 257.1513, 257.1533, 257.1551, 257.155, 257.155, 
    257.1554, 257.1544, 257.1556, 257.1558, 257.1553, 257.1583, 257.1574, 
    257.1583, 257.1577, 257.1439, 257.1446, 257.1442, 257.1449, 257.1444, 
    257.1465, 257.1472, 257.1502, 257.149, 257.151, 257.1492, 257.1495, 
    257.151, 257.1493, 257.1531, 257.1505, 257.1554, 257.1527, 257.1556, 
    257.1551, 257.1559, 257.1567, 257.1577, 257.1594, 257.159, 257.1605, 
    257.1456, 257.1464, 257.1464, 257.1473, 257.148, 257.1495, 257.1519, 
    257.151, 257.1526, 257.153, 257.1504, 257.1519, 257.147, 257.1478, 
    257.1474, 257.1456, 257.1512, 257.1483, 257.1536, 257.152, 257.1566, 
    257.1543, 257.1588, 257.1607, 257.1625, 257.1646, 257.1469, 257.1463, 
    257.1474, 257.1489, 257.1503, 257.1521, 257.1523, 257.1527, 257.1536, 
    257.1543, 257.1528, 257.1545, 257.1479, 257.1514, 257.1461, 257.1477, 
    257.1488, 257.1483, 257.1508, 257.1515, 257.1539, 257.1526, 257.1602, 
    257.1568, 257.1663, 257.1636, 257.1461, 257.1469, 257.1497, 257.1484, 
    257.1523, 257.1532, 257.154, 257.155, 257.1551, 257.1557, 257.1547, 
    257.1556, 257.1521, 257.1537, 257.1494, 257.1505, 257.15, 257.1495, 
    257.1511, 257.1528, 257.1528, 257.1534, 257.1549, 257.1523, 257.1606, 
    257.1554, 257.1478, 257.1494, 257.1496, 257.149, 257.1531, 257.1516, 
    257.1557, 257.1546, 257.1564, 257.1555, 257.1553, 257.1542, 257.1535, 
    257.1517, 257.1502, 257.1491, 257.1494, 257.1506, 257.1529, 257.1551, 
    257.1546, 257.1562, 257.152, 257.1537, 257.153, 257.1549, 257.1509, 
    257.1542, 257.1501, 257.1505, 257.1516, 257.1538, 257.1544, 257.1549, 
    257.1546, 257.153, 257.1527, 257.1516, 257.1512, 257.1504, 257.1497, 
    257.1503, 257.151, 257.153, 257.1548, 257.1567, 257.1572, 257.1594, 
    257.1576, 257.1606, 257.158, 257.1625, 257.1544, 257.1579, 257.1516, 
    257.1523, 257.1535, 257.1564, 257.1548, 257.1566, 257.1527, 257.1506, 
    257.1501, 257.1491, 257.1501, 257.1501, 257.151, 257.1507, 257.153, 
    257.1518, 257.1553, 257.1566, 257.1603, 257.1626, 257.1649, 257.166, 
    257.1663, 257.1664,
  259.1952, 259.1971, 259.1967, 259.1983, 259.1974, 259.1985, 259.1956, 
    259.1972, 259.1962, 259.1954, 259.2014, 259.1984, 259.2046, 259.2026, 
    259.2075, 259.2043, 259.2082, 259.2075, 259.2097, 259.2091, 259.212, 
    259.2101, 259.2135, 259.2115, 259.2118, 259.21, 259.199, 259.201, 
    259.1989, 259.1992, 259.199, 259.1975, 259.1967, 259.195, 259.1953, 
    259.1965, 259.1993, 259.1984, 259.2007, 259.2007, 259.2033, 259.2021, 
    259.2067, 259.2054, 259.2091, 259.2082, 259.2091, 259.2088, 259.2091, 
    259.2077, 259.2083, 259.2071, 259.2024, 259.2037, 259.1997, 259.1972, 
    259.1956, 259.1945, 259.1947, 259.195, 259.1966, 259.198, 259.1992, 
    259.2, 259.2007, 259.2029, 259.2042, 259.2069, 259.2064, 259.2072, 
    259.2081, 259.2094, 259.2092, 259.2098, 259.2072, 259.2089, 259.2061, 
    259.2069, 259.2008, 259.1986, 259.1976, 259.1968, 259.1948, 259.1962, 
    259.1956, 259.197, 259.1978, 259.1974, 259.2, 259.1989, 259.2042, 
    259.202, 259.208, 259.2065, 259.2083, 259.2074, 259.209, 259.2076, 
    259.21, 259.2105, 259.2102, 259.2116, 259.2075, 259.209, 259.1974, 
    259.1974, 259.1978, 259.1964, 259.1963, 259.195, 259.1962, 259.1966, 
    259.1978, 259.1986, 259.1993, 259.2008, 259.2025, 259.2049, 259.2066, 
    259.2078, 259.2071, 259.2077, 259.207, 259.2067, 259.2104, 259.2083, 
    259.2114, 259.2112, 259.2098, 259.2112, 259.1975, 259.1971, 259.1958, 
    259.1968, 259.1949, 259.196, 259.1966, 259.199, 259.1995, 259.2, 259.201, 
    259.2022, 259.2044, 259.2063, 259.2081, 259.208, 259.208, 259.2084, 
    259.2075, 259.2086, 259.2088, 259.2083, 259.2112, 259.2104, 259.2112, 
    259.2107, 259.1972, 259.1979, 259.1975, 259.1982, 259.1977, 259.1998, 
    259.2004, 259.2034, 259.2022, 259.2041, 259.2024, 259.2027, 259.2042, 
    259.2025, 259.2062, 259.2037, 259.2084, 259.2058, 259.2086, 259.2081, 
    259.2089, 259.2097, 259.2106, 259.2123, 259.2119, 259.2134, 259.1989, 
    259.1997, 259.1996, 259.2005, 259.2012, 259.2026, 259.205, 259.2041, 
    259.2057, 259.206, 259.2036, 259.2051, 259.2003, 259.201, 259.2006, 
    259.1989, 259.2043, 259.2015, 259.2066, 259.2051, 259.2096, 259.2073, 
    259.2117, 259.2136, 259.2154, 259.2174, 259.2002, 259.1996, 259.2007, 
    259.2021, 259.2034, 259.2052, 259.2054, 259.2057, 259.2066, 259.2074, 
    259.2058, 259.2076, 259.2012, 259.2045, 259.1994, 259.2009, 259.202, 
    259.2015, 259.204, 259.2046, 259.2069, 259.2057, 259.2131, 259.2098, 
    259.219, 259.2164, 259.1994, 259.2002, 259.2029, 259.2016, 259.2054, 
    259.2063, 259.207, 259.208, 259.2081, 259.2087, 259.2077, 259.2086, 
    259.2052, 259.2068, 259.2026, 259.2036, 259.2032, 259.2026, 259.2042, 
    259.2059, 259.2059, 259.2065, 259.2079, 259.2054, 259.2135, 259.2084, 
    259.201, 259.2025, 259.2028, 259.2022, 259.2062, 259.2047, 259.2087, 
    259.2076, 259.2094, 259.2085, 259.2083, 259.2072, 259.2065, 259.2048, 
    259.2034, 259.2023, 259.2025, 259.2037, 259.206, 259.2081, 259.2076, 
    259.2092, 259.2051, 259.2068, 259.2061, 259.2079, 259.2041, 259.2073, 
    259.2032, 259.2036, 259.2047, 259.2069, 259.2074, 259.2079, 259.2076, 
    259.206, 259.2058, 259.2047, 259.2043, 259.2035, 259.2028, 259.2035, 
    259.2041, 259.2061, 259.2078, 259.2097, 259.2101, 259.2123, 259.2105, 
    259.2135, 259.2109, 259.2154, 259.2075, 259.2109, 259.2047, 259.2054, 
    259.2066, 259.2094, 259.2079, 259.2096, 259.2058, 259.2038, 259.2033, 
    259.2023, 259.2033, 259.2032, 259.2042, 259.2039, 259.2061, 259.2049, 
    259.2083, 259.2096, 259.2132, 259.2154, 259.2177, 259.2188, 259.2191, 
    259.2192,
  261.3474, 261.3488, 261.3485, 261.3497, 261.349, 261.3498, 261.3477, 
    261.3488, 261.3481, 261.3475, 261.352, 261.3497, 261.3543, 261.3529, 
    261.3565, 261.3541, 261.357, 261.3565, 261.3582, 261.3577, 261.3599, 
    261.3584, 261.361, 261.3595, 261.3597, 261.3584, 261.3502, 261.3517, 
    261.3501, 261.3503, 261.3502, 261.3491, 261.3484, 261.3472, 261.3475, 
    261.3484, 261.3504, 261.3497, 261.3515, 261.3514, 261.3534, 261.3525, 
    261.3559, 261.3549, 261.3577, 261.357, 261.3577, 261.3575, 261.3577, 
    261.3567, 261.3571, 261.3562, 261.3527, 261.3537, 261.3507, 261.3489, 
    261.3477, 261.3469, 261.347, 261.3472, 261.3484, 261.3495, 261.3503, 
    261.3509, 261.3514, 261.3531, 261.354, 261.3561, 261.3557, 261.3563, 
    261.3569, 261.3579, 261.3578, 261.3582, 261.3563, 261.3576, 261.3555, 
    261.3561, 261.3516, 261.3499, 261.3492, 261.3486, 261.3471, 261.3481, 
    261.3477, 261.3487, 261.3493, 261.349, 261.3509, 261.3502, 261.3541, 
    261.3524, 261.3569, 261.3558, 261.3571, 261.3564, 261.3576, 261.3566, 
    261.3584, 261.3588, 261.3585, 261.3596, 261.3565, 261.3577, 261.349, 
    261.349, 261.3492, 261.3482, 261.3482, 261.3472, 261.3481, 261.3484, 
    261.3493, 261.3499, 261.3504, 261.3515, 261.3528, 261.3546, 261.3559, 
    261.3567, 261.3562, 261.3567, 261.3561, 261.3559, 261.3586, 261.3571, 
    261.3594, 261.3593, 261.3582, 261.3593, 261.3491, 261.3488, 261.3478, 
    261.3485, 261.3471, 261.3479, 261.3484, 261.3502, 261.3506, 261.3509, 
    261.3517, 261.3526, 261.3542, 261.3557, 261.357, 261.3569, 261.3569, 
    261.3572, 261.3565, 261.3573, 261.3575, 261.3571, 261.3593, 261.3586, 
    261.3593, 261.3589, 261.3489, 261.3494, 261.3491, 261.3496, 261.3492, 
    261.3508, 261.3513, 261.3535, 261.3525, 261.354, 261.3527, 261.3529, 
    261.354, 261.3528, 261.3556, 261.3536, 261.3572, 261.3553, 261.3573, 
    261.357, 261.3576, 261.3581, 261.3588, 261.3601, 261.3598, 261.3609, 
    261.3501, 261.3507, 261.3506, 261.3513, 261.3518, 261.3529, 261.3546, 
    261.354, 261.3552, 261.3554, 261.3536, 261.3547, 261.3511, 261.3517, 
    261.3514, 261.3501, 261.3541, 261.3521, 261.3559, 261.3547, 261.3581, 
    261.3564, 261.3596, 261.3611, 261.3624, 261.364, 261.351, 261.3506, 
    261.3514, 261.3525, 261.3535, 261.3548, 261.3549, 261.3552, 261.3559, 
    261.3564, 261.3553, 261.3565, 261.3518, 261.3543, 261.3505, 261.3516, 
    261.3524, 261.3521, 261.3539, 261.3543, 261.3561, 261.3552, 261.3607, 
    261.3582, 261.3651, 261.3632, 261.3505, 261.351, 261.3531, 261.3521, 
    261.3549, 261.3556, 261.3562, 261.3569, 261.357, 261.3574, 261.3567, 
    261.3574, 261.3548, 261.356, 261.3528, 261.3536, 261.3533, 261.3529, 
    261.3541, 261.3553, 261.3553, 261.3557, 261.3568, 261.3549, 261.361, 
    261.3572, 261.3517, 261.3528, 261.353, 261.3525, 261.3555, 261.3544, 
    261.3574, 261.3566, 261.3579, 261.3572, 261.3571, 261.3563, 261.3558, 
    261.3545, 261.3534, 261.3526, 261.3528, 261.3537, 261.3554, 261.357, 
    261.3566, 261.3578, 261.3547, 261.356, 261.3555, 261.3568, 261.3539, 
    261.3564, 261.3533, 261.3536, 261.3544, 261.3561, 261.3564, 261.3568, 
    261.3566, 261.3554, 261.3552, 261.3544, 261.3542, 261.3535, 261.353, 
    261.3535, 261.354, 261.3554, 261.3567, 261.3581, 261.3585, 261.3601, 
    261.3588, 261.361, 261.3591, 261.3624, 261.3565, 261.3591, 261.3545, 
    261.3549, 261.3558, 261.3579, 261.3568, 261.3581, 261.3552, 261.3537, 
    261.3534, 261.3527, 261.3534, 261.3533, 261.354, 261.3538, 261.3555, 
    261.3546, 261.3571, 261.3581, 261.3608, 261.3625, 261.3642, 261.3649, 
    261.3652, 261.3653,
  262.7316, 262.7321, 262.7321, 262.7325, 262.7323, 262.7326, 262.7317, 
    262.7322, 262.7319, 262.7316, 262.7334, 262.7325, 262.7344, 262.7338, 
    262.7353, 262.7343, 262.7355, 262.7352, 262.7359, 262.7357, 262.7366, 
    262.736, 262.7371, 262.7365, 262.7366, 262.736, 262.7327, 262.7333, 
    262.7327, 262.7328, 262.7327, 262.7323, 262.732, 262.7315, 262.7316, 
    262.732, 262.7328, 262.7325, 262.7332, 262.7332, 262.734, 262.7336, 
    262.735, 262.7346, 262.7357, 262.7355, 262.7357, 262.7357, 262.7357, 
    262.7353, 262.7355, 262.7351, 262.7337, 262.7341, 262.7329, 262.7322, 
    262.7317, 262.7314, 262.7314, 262.7315, 262.732, 262.7324, 262.7328, 
    262.733, 262.7332, 262.7339, 262.7343, 262.7351, 262.7349, 262.7352, 
    262.7354, 262.7358, 262.7358, 262.736, 262.7352, 262.7357, 262.7349, 
    262.7351, 262.7333, 262.7326, 262.7323, 262.7321, 262.7315, 262.7319, 
    262.7317, 262.7321, 262.7324, 262.7322, 262.733, 262.7327, 262.7343, 
    262.7336, 262.7354, 262.735, 262.7355, 262.7352, 262.7357, 262.7353, 
    262.736, 262.7362, 262.7361, 262.7365, 262.7353, 262.7357, 262.7322, 
    262.7322, 262.7324, 262.7319, 262.7319, 262.7315, 262.7319, 262.732, 
    262.7324, 262.7326, 262.7328, 262.7332, 262.7338, 262.7345, 262.735, 
    262.7354, 262.7351, 262.7353, 262.7351, 262.735, 262.7361, 262.7355, 
    262.7365, 262.7364, 262.736, 262.7364, 262.7323, 262.7321, 262.7318, 
    262.7321, 262.7315, 262.7318, 262.732, 262.7327, 262.7329, 262.733, 
    262.7333, 262.7337, 262.7343, 262.7349, 262.7354, 262.7354, 262.7354, 
    262.7355, 262.7352, 262.7356, 262.7357, 262.7355, 262.7364, 262.7361, 
    262.7364, 262.7362, 262.7322, 262.7324, 262.7323, 262.7325, 262.7323, 
    262.733, 262.7332, 262.734, 262.7337, 262.7343, 262.7337, 262.7338, 
    262.7343, 262.7338, 262.7349, 262.7341, 262.7355, 262.7348, 262.7356, 
    262.7354, 262.7357, 262.7359, 262.7362, 262.7367, 262.7366, 262.737, 
    262.7327, 262.7329, 262.7329, 262.7332, 262.7334, 262.7338, 262.7345, 
    262.7342, 262.7347, 262.7348, 262.7341, 262.7345, 262.7331, 262.7333, 
    262.7332, 262.7327, 262.7343, 262.7335, 262.735, 262.7346, 262.7359, 
    262.7352, 262.7365, 262.7371, 262.7376, 262.7383, 262.7331, 262.7329, 
    262.7332, 262.7336, 262.734, 262.7346, 262.7346, 262.7347, 262.735, 
    262.7352, 262.7348, 262.7353, 262.7334, 262.7344, 262.7328, 262.7333, 
    262.7336, 262.7335, 262.7342, 262.7344, 262.7351, 262.7347, 262.7369, 
    262.736, 262.7387, 262.7379, 262.7328, 262.7331, 262.7339, 262.7335, 
    262.7346, 262.7349, 262.7351, 262.7354, 262.7354, 262.7356, 262.7353, 
    262.7356, 262.7346, 262.735, 262.7338, 262.7341, 262.7339, 262.7338, 
    262.7343, 262.7348, 262.7348, 262.735, 262.7354, 262.7346, 262.7371, 
    262.7355, 262.7333, 262.7338, 262.7338, 262.7337, 262.7349, 262.7344, 
    262.7356, 262.7353, 262.7358, 262.7356, 262.7355, 262.7352, 262.735, 
    262.7344, 262.734, 262.7337, 262.7338, 262.7341, 262.7348, 262.7354, 
    262.7353, 262.7358, 262.7345, 262.735, 262.7349, 262.7354, 262.7342, 
    262.7352, 262.734, 262.7341, 262.7344, 262.7351, 262.7352, 262.7354, 
    262.7353, 262.7348, 262.7347, 262.7344, 262.7343, 262.7341, 262.7339, 
    262.734, 262.7343, 262.7348, 262.7354, 262.7359, 262.7361, 262.7367, 
    262.7362, 262.7371, 262.7363, 262.7377, 262.7353, 262.7363, 262.7344, 
    262.7346, 262.735, 262.7358, 262.7354, 262.7359, 262.7347, 262.7341, 
    262.734, 262.7337, 262.734, 262.734, 262.7343, 262.7342, 262.7348, 
    262.7345, 262.7355, 262.7359, 262.737, 262.7377, 262.7383, 262.7387, 
    262.7388, 262.7388,
  263.1134, 263.1135, 263.1135, 263.1136, 263.1135, 263.1136, 263.1134, 
    263.1135, 263.1135, 263.1134, 263.1137, 263.1136, 263.1138, 263.1137, 
    263.114, 263.1138, 263.114, 263.114, 263.1141, 263.114, 263.1142, 
    263.1141, 263.1143, 263.1142, 263.1142, 263.1141, 263.1136, 263.1137, 
    263.1136, 263.1136, 263.1136, 263.1135, 263.1135, 263.1134, 263.1134, 
    263.1135, 263.1136, 263.1136, 263.1137, 263.1137, 263.1138, 263.1137, 
    263.1139, 263.1139, 263.114, 263.114, 263.114, 263.114, 263.114, 263.114, 
    263.114, 263.114, 263.1137, 263.1138, 263.1136, 263.1135, 263.1134, 
    263.1134, 263.1134, 263.1134, 263.1135, 263.1136, 263.1136, 263.1136, 
    263.1137, 263.1138, 263.1138, 263.114, 263.1139, 263.114, 263.114, 
    263.1141, 263.114, 263.1141, 263.114, 263.114, 263.1139, 263.114, 
    263.1137, 263.1136, 263.1135, 263.1135, 263.1134, 263.1135, 263.1134, 
    263.1135, 263.1135, 263.1135, 263.1136, 263.1136, 263.1138, 263.1137, 
    263.114, 263.1139, 263.114, 263.114, 263.114, 263.114, 263.1141, 
    263.1141, 263.1141, 263.1142, 263.114, 263.114, 263.1135, 263.1135, 
    263.1135, 263.1135, 263.1135, 263.1134, 263.1135, 263.1135, 263.1135, 
    263.1136, 263.1136, 263.1137, 263.1137, 263.1139, 263.1139, 263.114, 
    263.114, 263.114, 263.114, 263.1139, 263.1141, 263.114, 263.1142, 
    263.1141, 263.1141, 263.1141, 263.1135, 263.1135, 263.1134, 263.1135, 
    263.1134, 263.1135, 263.1135, 263.1136, 263.1136, 263.1136, 263.1137, 
    263.1137, 263.1138, 263.1139, 263.114, 263.114, 263.114, 263.114, 
    263.114, 263.114, 263.114, 263.114, 263.1141, 263.1141, 263.1141, 
    263.1141, 263.1135, 263.1135, 263.1135, 263.1136, 263.1135, 263.1136, 
    263.1136, 263.1138, 263.1137, 263.1138, 263.1137, 263.1138, 263.1138, 
    263.1137, 263.1139, 263.1138, 263.114, 263.1139, 263.114, 263.114, 
    263.114, 263.1141, 263.1141, 263.1142, 263.1142, 263.1143, 263.1136, 
    263.1136, 263.1136, 263.1136, 263.1137, 263.1137, 263.1139, 263.1138, 
    263.1139, 263.1139, 263.1138, 263.1139, 263.1136, 263.1137, 263.1136, 
    263.1136, 263.1138, 263.1137, 263.1139, 263.1139, 263.1141, 263.114, 
    263.1142, 263.1143, 263.1143, 263.1144, 263.1136, 263.1136, 263.1136, 
    263.1137, 263.1138, 263.1139, 263.1139, 263.1139, 263.1139, 263.114, 
    263.1139, 263.114, 263.1137, 263.1138, 263.1136, 263.1137, 263.1137, 
    263.1137, 263.1138, 263.1138, 263.114, 263.1139, 263.1142, 263.1141, 
    263.1145, 263.1144, 263.1136, 263.1136, 263.1138, 263.1137, 263.1139, 
    263.1139, 263.114, 263.114, 263.114, 263.114, 263.114, 263.114, 263.1139, 
    263.114, 263.1137, 263.1138, 263.1138, 263.1137, 263.1138, 263.1139, 
    263.1139, 263.1139, 263.114, 263.1139, 263.1143, 263.114, 263.1137, 
    263.1137, 263.1138, 263.1137, 263.1139, 263.1139, 263.114, 263.114, 
    263.1141, 263.114, 263.114, 263.114, 263.1139, 263.1139, 263.1138, 
    263.1137, 263.1137, 263.1138, 263.1139, 263.114, 263.114, 263.114, 
    263.1139, 263.114, 263.1139, 263.114, 263.1138, 263.114, 263.1138, 
    263.1138, 263.1139, 263.114, 263.114, 263.114, 263.114, 263.1139, 
    263.1139, 263.1138, 263.1138, 263.1138, 263.1138, 263.1138, 263.1138, 
    263.1139, 263.114, 263.1141, 263.1141, 263.1142, 263.1141, 263.1143, 
    263.1141, 263.1143, 263.114, 263.1141, 263.1139, 263.1139, 263.1139, 
    263.1141, 263.114, 263.1141, 263.1139, 263.1138, 263.1138, 263.1137, 
    263.1138, 263.1138, 263.1138, 263.1138, 263.1139, 263.1139, 263.114, 
    263.1141, 263.1142, 263.1143, 263.1144, 263.1145, 263.1145, 263.1145,
  263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 263.149, 
    263.149, 263.149,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.0269, 263.0419, 263.039, 263.051, 263.0444, 263.0522, 263.03, 263.0425, 
    263.0345, 263.0283, 263.0743, 263.0516, 263.0979, 263.0835, 263.1196, 
    263.0956, 263.1245, 263.119, 263.1356, 263.1308, 263.152, 263.1378, 
    263.163, 263.1486, 263.1508, 263.1373, 263.0562, 263.0715, 263.0553, 
    263.0575, 263.0565, 263.0445, 263.0385, 263.0258, 263.0281, 263.0374, 
    263.0584, 263.0513, 263.0693, 263.0689, 263.0888, 263.0798, 263.1132, 
    263.1037, 263.131, 263.1242, 263.1307, 263.1287, 263.1307, 263.1207, 
    263.125, 263.1161, 263.0815, 263.0917, 263.0612, 263.0428, 263.0305, 
    263.0218, 263.023, 263.0254, 263.0374, 263.0488, 263.0574, 263.0631, 
    263.0688, 263.0859, 263.0949, 263.1151, 263.1115, 263.1176, 263.1235, 
    263.1333, 263.1317, 263.136, 263.1175, 263.1298, 263.1094, 263.115, 
    263.0703, 263.0533, 263.0459, 263.0396, 263.024, 263.0347, 263.0305, 
    263.0406, 263.047, 263.0438, 263.0633, 263.0558, 263.0955, 263.0784, 
    263.1228, 263.1122, 263.1253, 263.1187, 263.1301, 263.1198, 263.1377, 
    263.1415, 263.1389, 263.1491, 263.1192, 263.1307, 263.0437, 263.0443, 
    263.0467, 263.0361, 263.0354, 263.0258, 263.0344, 263.038, 263.0474, 
    263.0529, 263.0581, 263.0695, 263.0823, 263.1001, 263.1129, 263.1214, 
    263.1162, 263.1208, 263.1157, 263.1132, 263.1401, 263.125, 263.1476, 
    263.1464, 263.1361, 263.1465, 263.0446, 263.0417, 263.0313, 263.0394, 
    263.0247, 263.0329, 263.0377, 263.0559, 263.0599, 263.0636, 263.0709, 
    263.0803, 263.0967, 263.1109, 263.1238, 263.1229, 263.1232, 263.1261, 
    263.1189, 263.1273, 263.1287, 263.125, 263.1462, 263.1402, 263.1464, 
    263.1424, 263.0426, 263.0476, 263.0449, 263.05, 263.0464, 263.0623, 
    263.067, 263.0892, 263.0801, 263.0945, 263.0816, 263.0839, 263.095, 
    263.0823, 263.1101, 263.0912, 263.1262, 263.1074, 263.1274, 263.1238, 
    263.1298, 263.1351, 263.1418, 263.1543, 263.1514, 263.1618, 263.0551, 
    263.0615, 263.0609, 263.0677, 263.0727, 263.0835, 263.1007, 263.0943, 
    263.1061, 263.1085, 263.0905, 263.1016, 263.0658, 263.0716, 263.0681, 
    263.0555, 263.0958, 263.0752, 263.1131, 263.102, 263.1343, 263.1183, 
    263.1498, 263.1632, 263.1759, 263.1906, 263.065, 263.0606, 263.0685, 
    263.0793, 263.0894, 263.1027, 263.104, 263.1065, 263.113, 263.1184, 
    263.1073, 263.1198, 263.0729, 263.0975, 263.059, 263.0706, 263.0787, 
    263.0752, 263.0935, 263.0978, 263.1153, 263.1063, 263.1599, 263.1362, 
    263.2018, 263.1836, 263.0591, 263.065, 263.0855, 263.0758, 263.1036, 
    263.1104, 263.1159, 263.123, 263.1237, 263.128, 263.1211, 263.1277, 
    263.1027, 263.1139, 263.0832, 263.0907, 263.0872, 263.0835, 263.0951, 
    263.1075, 263.1078, 263.1117, 263.1228, 263.1037, 263.1629, 263.1263, 
    263.0714, 263.0828, 263.0844, 263.08, 263.1097, 263.099, 263.1278, 
    263.1201, 263.1328, 263.1265, 263.1255, 263.1174, 263.1123, 263.0995, 
    263.089, 263.0807, 263.0826, 263.0918, 263.1082, 263.1238, 263.1204, 
    263.1319, 263.1016, 263.1143, 263.1093, 263.1222, 263.0941, 263.1179, 
    263.088, 263.0906, 263.0988, 263.1151, 263.1187, 263.1226, 263.1202, 
    263.1086, 263.1068, 263.0986, 263.0963, 263.0901, 263.0849, 263.0896, 
    263.0946, 263.1087, 263.1214, 263.1352, 263.1386, 263.1546, 263.1415, 
    263.1631, 263.1447, 263.1766, 263.1194, 263.1442, 263.0991, 263.104, 
    263.1128, 263.133, 263.1221, 263.1348, 263.1067, 263.092, 263.0883, 
    263.0812, 263.0884, 263.0879, 263.0948, 263.0926, 263.1091, 263.1002, 
    263.1255, 263.1347, 263.1607, 263.1765, 263.1927, 263.1998, 263.202, 
    263.2029 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9618, 253.9627, 253.9626, 253.9633, 253.9629, 253.9634, 253.962, 
    253.9628, 253.9623, 253.9619, 253.9647, 253.9633, 253.9662, 253.9653, 
    253.9675, 253.966, 253.9679, 253.9675, 253.9686, 253.9683, 253.9696, 
    253.9687, 253.9703, 253.9694, 253.9695, 253.9687, 253.9636, 253.9645, 
    253.9636, 253.9637, 253.9636, 253.9629, 253.9625, 253.9618, 253.9619, 
    253.9624, 253.9637, 253.9633, 253.9644, 253.9644, 253.9656, 253.9651, 
    253.9672, 253.9666, 253.9683, 253.9678, 253.9683, 253.9681, 253.9683, 
    253.9676, 253.9679, 253.9673, 253.9652, 253.9658, 253.9639, 253.9628, 
    253.962, 253.9615, 253.9616, 253.9617, 253.9624, 253.9632, 253.9637, 
    253.9641, 253.9644, 253.9654, 253.966, 253.9673, 253.9671, 253.9674, 
    253.9678, 253.9684, 253.9683, 253.9686, 253.9674, 253.9682, 253.9669, 
    253.9673, 253.9644, 253.9634, 253.963, 253.9626, 253.9616, 253.9623, 
    253.962, 253.9627, 253.963, 253.9629, 253.9641, 253.9636, 253.966, 
    253.965, 253.9678, 253.9671, 253.9679, 253.9675, 253.9682, 253.9676, 
    253.9687, 253.9689, 253.9688, 253.9694, 253.9675, 253.9683, 253.9628, 
    253.9629, 253.963, 253.9624, 253.9623, 253.9617, 253.9623, 253.9625, 
    253.9631, 253.9634, 253.9637, 253.9644, 253.9652, 253.9663, 253.9671, 
    253.9677, 253.9674, 253.9677, 253.9673, 253.9672, 253.9689, 253.9679, 
    253.9693, 253.9693, 253.9686, 253.9693, 253.9629, 253.9627, 253.9621, 
    253.9626, 253.9617, 253.9622, 253.9625, 253.9636, 253.9639, 253.9641, 
    253.9645, 253.9651, 253.9661, 253.967, 253.9678, 253.9678, 253.9678, 
    253.968, 253.9675, 253.968, 253.9681, 253.9679, 253.9693, 253.9689, 
    253.9693, 253.969, 253.9628, 253.9631, 253.9629, 253.9632, 253.963, 
    253.964, 253.9643, 253.9656, 253.9651, 253.966, 253.9652, 253.9653, 
    253.966, 253.9652, 253.9669, 253.9658, 253.968, 253.9668, 253.9681, 
    253.9678, 253.9682, 253.9685, 253.969, 253.9698, 253.9696, 253.9702, 
    253.9635, 253.9639, 253.9639, 253.9643, 253.9646, 253.9653, 253.9664, 
    253.966, 253.9667, 253.9669, 253.9657, 253.9664, 253.9642, 253.9646, 
    253.9644, 253.9636, 253.966, 253.9648, 253.9671, 253.9665, 253.9685, 
    253.9675, 253.9695, 253.9703, 253.9711, 253.9721, 253.9642, 253.9639, 
    253.9644, 253.965, 253.9657, 253.9665, 253.9666, 253.9667, 253.9671, 
    253.9675, 253.9668, 253.9676, 253.9646, 253.9662, 253.9638, 253.9645, 
    253.965, 253.9648, 253.9659, 253.9662, 253.9673, 253.9667, 253.9701, 
    253.9686, 253.9728, 253.9716, 253.9638, 253.9642, 253.9654, 253.9648, 
    253.9666, 253.967, 253.9673, 253.9678, 253.9678, 253.9681, 253.9677, 
    253.9681, 253.9665, 253.9672, 253.9653, 253.9657, 253.9655, 253.9653, 
    253.966, 253.9668, 253.9668, 253.9671, 253.9677, 253.9666, 253.9702, 
    253.9679, 253.9646, 253.9652, 253.9654, 253.9651, 253.9669, 253.9663, 
    253.9681, 253.9676, 253.9684, 253.968, 253.9679, 253.9674, 253.9671, 
    253.9663, 253.9656, 253.9651, 253.9653, 253.9658, 253.9668, 253.9678, 
    253.9676, 253.9683, 253.9664, 253.9672, 253.9669, 253.9677, 253.966, 
    253.9674, 253.9656, 253.9657, 253.9662, 253.9673, 253.9675, 253.9677, 
    253.9676, 253.9669, 253.9668, 253.9662, 253.9661, 253.9657, 253.9654, 
    253.9657, 253.966, 253.9669, 253.9677, 253.9686, 253.9688, 253.9697, 
    253.9689, 253.9703, 253.9691, 253.9711, 253.9675, 253.9691, 253.9663, 
    253.9666, 253.9671, 253.9684, 253.9677, 253.9685, 253.9668, 253.9658, 
    253.9656, 253.9652, 253.9656, 253.9656, 253.966, 253.9659, 253.9669, 
    253.9664, 253.9679, 253.9685, 253.9702, 253.9712, 253.9722, 253.9727, 
    253.9728, 253.9729 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1405833, 0.1405927, 0.1405909, 0.1405984, 0.1405943, 0.1405992, 
    0.1405853, 0.140593, 0.1405881, 0.1405843, 0.1406128, 0.1405988, 
    0.1406282, 0.1406191, 0.1406423, 0.1406267, 0.1406454, 0.140642, 
    0.1406528, 0.1406497, 0.1406633, 0.1406543, 0.1406706, 0.1406612, 
    0.1406626, 0.1406539, 0.1406018, 0.140611, 0.1406012, 0.1406025, 
    0.140602, 0.1405944, 0.1405904, 0.1405827, 0.1405842, 0.1405899, 
    0.1406031, 0.1405987, 0.1406101, 0.1406099, 0.1406225, 0.1406168, 
    0.1406382, 0.1406322, 0.1406499, 0.1406454, 0.1406496, 0.1406484, 
    0.1406496, 0.1406431, 0.1406459, 0.1406402, 0.1406178, 0.1406243, 
    0.1406049, 0.1405931, 0.1405856, 0.1405802, 0.140581, 0.1405824, 
    0.1405899, 0.1405971, 0.1406026, 0.1406062, 0.1406098, 0.1406204, 
    0.1406263, 0.1406394, 0.1406372, 0.140641, 0.1406449, 0.1406513, 
    0.1406503, 0.1406531, 0.140641, 0.140649, 0.1406359, 0.1406394, 
    0.1406102, 0.1405999, 0.1405951, 0.1405913, 0.1405815, 0.1405882, 
    0.1405856, 0.140592, 0.140596, 0.140594, 0.1406063, 0.1406015, 0.1406267, 
    0.1406158, 0.1406445, 0.1406376, 0.1406462, 0.1406418, 0.1406492, 
    0.1406426, 0.1406541, 0.1406566, 0.1406549, 0.1406616, 0.1406422, 
    0.1406496, 0.140594, 0.1405943, 0.1405958, 0.140589, 0.1405887, 
    0.1405827, 0.1405881, 0.1405903, 0.1405963, 0.1405997, 0.140603, 
    0.1406103, 0.1406183, 0.1406297, 0.1406381, 0.1406436, 0.1406403, 
    0.1406432, 0.1406399, 0.1406383, 0.1406557, 0.1406459, 0.1406607, 
    0.1406599, 0.1406531, 0.14066, 0.1405945, 0.1405927, 0.1405861, 
    0.1405912, 0.140582, 0.1405871, 0.14059, 0.1406015, 0.1406042, 0.1406065, 
    0.1406112, 0.1406171, 0.1406275, 0.1406367, 0.1406452, 0.1406446, 
    0.1406448, 0.1406466, 0.140642, 0.1406474, 0.1406482, 0.1406459, 
    0.1406597, 0.1406558, 0.1406599, 0.1406573, 0.1405933, 0.1405964, 
    0.1405947, 0.1405979, 0.1405956, 0.1406055, 0.1406085, 0.1406226, 
    0.140617, 0.1406261, 0.1406179, 0.1406194, 0.1406262, 0.1406184, 
    0.1406361, 0.1406239, 0.1406467, 0.1406342, 0.1406475, 0.1406452, 
    0.1406491, 0.1406525, 0.1406569, 0.1406649, 0.1406631, 0.1406699, 
    0.1406011, 0.1406051, 0.1406048, 0.1406091, 0.1406122, 0.1406192, 
    0.1406302, 0.1406261, 0.1406337, 0.1406353, 0.1406237, 0.1406307, 
    0.1406078, 0.1406114, 0.1406094, 0.1406013, 0.1406269, 0.1406137, 
    0.1406382, 0.140631, 0.140652, 0.1406414, 0.1406621, 0.1406706, 
    0.1406792, 0.1406887, 0.1406074, 0.1406047, 0.1406096, 0.1406163, 
    0.1406229, 0.1406315, 0.1406324, 0.140634, 0.1406382, 0.1406417, 
    0.1406343, 0.1406425, 0.140612, 0.1406281, 0.1406035, 0.1406108, 
    0.140616, 0.1406138, 0.1406256, 0.1406284, 0.1406396, 0.1406338, 
    0.1406684, 0.1406531, 0.1406963, 0.1406841, 0.1406037, 0.1406074, 
    0.1406204, 0.1406142, 0.1406321, 0.1406364, 0.1406401, 0.1406446, 
    0.1406451, 0.1406478, 0.1406434, 0.1406477, 0.1406315, 0.1406387, 
    0.140619, 0.1406237, 0.1406216, 0.1406192, 0.1406266, 0.1406344, 
    0.1406348, 0.1406372, 0.1406439, 0.1406322, 0.1406701, 0.1406463, 
    0.1406115, 0.1406185, 0.1406197, 0.140617, 0.140636, 0.1406291, 
    0.1406478, 0.1406427, 0.140651, 0.1406469, 0.1406463, 0.140641, 
    0.1406377, 0.1406294, 0.1406226, 0.1406174, 0.1406186, 0.1406244, 
    0.140635, 0.1406451, 0.1406429, 0.1406504, 0.1406308, 0.1406389, 
    0.1406357, 0.1406441, 0.1406259, 0.1406409, 0.1406221, 0.1406237, 
    0.1406289, 0.1406393, 0.1406419, 0.1406443, 0.1406429, 0.1406353, 
    0.1406341, 0.1406288, 0.1406273, 0.1406234, 0.1406201, 0.140623, 
    0.1406262, 0.1406353, 0.1406435, 0.1406525, 0.1406548, 0.1406649, 
    0.1406564, 0.1406702, 0.1406581, 0.1406792, 0.140642, 0.1406581, 
    0.1406292, 0.1406324, 0.1406379, 0.1406509, 0.140644, 0.1406521, 
    0.1406341, 0.1406245, 0.1406222, 0.1406177, 0.1406223, 0.140622, 
    0.1406264, 0.140625, 0.1406356, 0.1406299, 0.1406462, 0.1406521, 
    0.1406691, 0.1406795, 0.1406903, 0.140695, 0.1406965, 0.1406971,
  0.1468979, 0.146909, 0.1469069, 0.1469157, 0.1469109, 0.1469167, 0.1469003, 
    0.1469094, 0.1469036, 0.146899, 0.1469328, 0.1469162, 0.1469509, 
    0.1469401, 0.1469675, 0.1469491, 0.1469713, 0.1469672, 0.14698, 
    0.1469764, 0.1469925, 0.1469817, 0.1470011, 0.14699, 0.1469917, 
    0.1469813, 0.1469197, 0.1469307, 0.146919, 0.1469206, 0.1469199, 
    0.1469109, 0.1469063, 0.1468972, 0.1468989, 0.1469056, 0.1469213, 
    0.1469161, 0.1469295, 0.1469292, 0.1469442, 0.1469374, 0.1469627, 
    0.1469556, 0.1469765, 0.1469712, 0.1469762, 0.1469747, 0.1469762, 
    0.1469685, 0.1469718, 0.146965, 0.1469387, 0.1469463, 0.1469234, 
    0.1469094, 0.1469006, 0.1468942, 0.1468951, 0.1468968, 0.1469057, 
    0.1469142, 0.1469206, 0.1469249, 0.1469292, 0.1469417, 0.1469487, 
    0.1469641, 0.1469615, 0.1469661, 0.1469707, 0.1469782, 0.146977, 
    0.1469803, 0.1469661, 0.1469755, 0.1469599, 0.1469641, 0.1469298, 
    0.1469175, 0.1469118, 0.1469073, 0.1468958, 0.1469037, 0.1469006, 
    0.1469081, 0.1469128, 0.1469105, 0.146925, 0.1469194, 0.1469491, 
    0.1469363, 0.1469701, 0.146962, 0.1469721, 0.146967, 0.1469757, 
    0.1469679, 0.1469816, 0.1469845, 0.1469825, 0.1469905, 0.1469674, 
    0.1469762, 0.1469104, 0.1469108, 0.1469126, 0.1469047, 0.1469042, 
    0.1468971, 0.1469035, 0.1469062, 0.1469132, 0.1469172, 0.1469211, 
    0.1469297, 0.1469392, 0.1469527, 0.1469625, 0.1469691, 0.1469651, 
    0.1469687, 0.1469647, 0.1469629, 0.1469834, 0.1469718, 0.1469893, 
    0.1469884, 0.1469804, 0.1469885, 0.1469111, 0.1469089, 0.1469012, 
    0.1469072, 0.1468964, 0.1469024, 0.1469058, 0.1469194, 0.1469225, 
    0.1469252, 0.1469307, 0.1469378, 0.1469501, 0.1469609, 0.146971, 
    0.1469702, 0.1469705, 0.1469727, 0.1469672, 0.1469736, 0.1469746, 
    0.1469719, 0.1469882, 0.1469835, 0.1469883, 0.1469853, 0.1469096, 
    0.1469133, 0.1469113, 0.146915, 0.1469124, 0.1469241, 0.1469276, 
    0.1469443, 0.1469376, 0.1469484, 0.1469387, 0.1469404, 0.1469486, 
    0.1469393, 0.1469602, 0.1469458, 0.1469728, 0.1469581, 0.1469737, 
    0.1469709, 0.1469755, 0.1469796, 0.1469849, 0.1469944, 0.1469922, 
    0.1470003, 0.1469188, 0.1469236, 0.1469233, 0.1469283, 0.146932, 
    0.1469402, 0.1469532, 0.1469484, 0.1469574, 0.1469592, 0.1469455, 
    0.1469538, 0.1469268, 0.1469311, 0.1469286, 0.1469192, 0.1469493, 
    0.1469337, 0.1469627, 0.1469542, 0.146979, 0.1469666, 0.146991, 
    0.1470012, 0.1470114, 0.1470227, 0.1469263, 0.1469231, 0.1469289, 
    0.1469369, 0.1469446, 0.1469547, 0.1469558, 0.1469577, 0.1469627, 
    0.1469668, 0.1469582, 0.1469678, 0.1469318, 0.1469507, 0.1469217, 
    0.1469303, 0.1469365, 0.1469339, 0.1469478, 0.1469511, 0.1469643, 
    0.1469575, 0.1469986, 0.1469803, 0.1470317, 0.1470172, 0.1469219, 
    0.1469263, 0.1469416, 0.1469343, 0.1469554, 0.1469606, 0.1469649, 
    0.1469703, 0.1469709, 0.1469741, 0.1469689, 0.1469739, 0.1469547, 
    0.1469633, 0.14694, 0.1469456, 0.146943, 0.1469402, 0.146949, 0.1469583, 
    0.1469586, 0.1469616, 0.1469696, 0.1469555, 0.1470006, 0.1469724, 
    0.1469312, 0.1469395, 0.1469409, 0.1469376, 0.1469601, 0.1469519, 
    0.146974, 0.1469681, 0.1469779, 0.146973, 0.1469723, 0.146966, 0.1469621, 
    0.1469522, 0.1469443, 0.1469381, 0.1469395, 0.1469464, 0.1469589, 
    0.1469709, 0.1469682, 0.1469771, 0.1469539, 0.1469635, 0.1469598, 
    0.1469697, 0.1469482, 0.1469659, 0.1469436, 0.1469456, 0.1469517, 
    0.1469641, 0.1469671, 0.14697, 0.1469682, 0.1469592, 0.1469578, 
    0.1469516, 0.1469498, 0.1469452, 0.1469412, 0.1469448, 0.1469485, 
    0.1469593, 0.146969, 0.1469796, 0.1469823, 0.1469944, 0.1469843, 
    0.1470007, 0.1469864, 0.1470114, 0.1469672, 0.1469864, 0.1469521, 
    0.1469558, 0.1469623, 0.1469778, 0.1469696, 0.1469793, 0.1469578, 
    0.1469465, 0.1469438, 0.1469384, 0.1469439, 0.1469435, 0.1469488, 
    0.1469471, 0.1469597, 0.1469529, 0.1469722, 0.1469792, 0.1469994, 
    0.1470117, 0.1470245, 0.1470301, 0.1470319, 0.1470326,
  0.1564216, 0.1564342, 0.1564318, 0.1564419, 0.1564364, 0.1564429, 
    0.1564243, 0.1564347, 0.1564281, 0.1564229, 0.1564614, 0.1564424, 
    0.156482, 0.1564696, 0.156501, 0.15648, 0.1565053, 0.1565006, 0.1565152, 
    0.156511, 0.1565295, 0.1565172, 0.1565394, 0.1565267, 0.1565286, 
    0.1565167, 0.1564464, 0.156459, 0.1564456, 0.1564474, 0.1564466, 
    0.1564364, 0.1564312, 0.1564208, 0.1564227, 0.1564304, 0.1564482, 
    0.1564422, 0.1564576, 0.1564572, 0.1564743, 0.1564666, 0.1564955, 
    0.1564873, 0.1565112, 0.1565051, 0.1565109, 0.1565092, 0.1565109, 
    0.156502, 0.1565058, 0.1564981, 0.156468, 0.1564767, 0.1564506, 
    0.1564348, 0.1564247, 0.1564174, 0.1564185, 0.1564204, 0.1564305, 
    0.1564401, 0.1564474, 0.1564523, 0.1564572, 0.1564715, 0.1564794, 
    0.1564971, 0.156494, 0.1564993, 0.1565045, 0.1565132, 0.1565118, 
    0.1565156, 0.1564993, 0.15651, 0.1564922, 0.1564971, 0.156458, 0.1564439, 
    0.1564375, 0.1564323, 0.1564192, 0.1564282, 0.1564246, 0.1564332, 
    0.1564386, 0.1564359, 0.1564524, 0.156446, 0.1564799, 0.1564653, 
    0.1565039, 0.1564946, 0.1565062, 0.1565003, 0.1565103, 0.1565013, 
    0.156517, 0.1565204, 0.1565181, 0.1565272, 0.1565008, 0.1565108, 
    0.1564358, 0.1564363, 0.1564383, 0.1564293, 0.1564288, 0.1564207, 
    0.1564279, 0.156431, 0.1564389, 0.1564435, 0.156448, 0.1564577, 
    0.1564686, 0.156484, 0.1564952, 0.1565028, 0.1564982, 0.1565022, 
    0.1564977, 0.1564956, 0.1565191, 0.1565058, 0.1565259, 0.1565248, 
    0.1565157, 0.1565249, 0.1564366, 0.1564341, 0.1564254, 0.1564322, 
    0.1564198, 0.1564267, 0.1564306, 0.156446, 0.1564495, 0.1564527, 
    0.1564589, 0.1564669, 0.156481, 0.1564934, 0.1565049, 0.156504, 
    0.1565043, 0.1565068, 0.1565006, 0.1565079, 0.1565091, 0.1565059, 
    0.1565246, 0.1565193, 0.1565247, 0.1565213, 0.1564349, 0.1564391, 
    0.1564368, 0.1564411, 0.1564381, 0.1564514, 0.1564554, 0.1564745, 
    0.1564668, 0.1564792, 0.1564681, 0.15647, 0.1564793, 0.1564687, 
    0.1564926, 0.1564762, 0.1565069, 0.1564902, 0.156508, 0.1565048, 
    0.1565101, 0.1565148, 0.1565208, 0.1565317, 0.1565292, 0.1565384, 
    0.1564454, 0.1564508, 0.1564504, 0.1564562, 0.1564604, 0.1564697, 
    0.1564846, 0.156479, 0.1564894, 0.1564914, 0.1564758, 0.1564853, 
    0.1564545, 0.1564594, 0.1564565, 0.1564458, 0.1564802, 0.1564624, 
    0.1564954, 0.1564857, 0.1565141, 0.1564999, 0.1565278, 0.1565395, 
    0.1565511, 0.1565642, 0.1564539, 0.1564502, 0.1564569, 0.156466, 
    0.1564748, 0.1564863, 0.1564875, 0.1564897, 0.1564953, 0.1565001, 
    0.1564903, 0.1565013, 0.1564603, 0.1564818, 0.1564487, 0.1564585, 
    0.1564655, 0.1564625, 0.1564784, 0.1564821, 0.1564973, 0.1564895, 
    0.1565365, 0.1565156, 0.1565745, 0.1565579, 0.1564489, 0.1564539, 
    0.1564714, 0.1564631, 0.1564871, 0.156493, 0.1564979, 0.1565041, 
    0.1565048, 0.1565084, 0.1565025, 0.1565082, 0.1564863, 0.1564961, 
    0.1564695, 0.1564759, 0.156473, 0.1564697, 0.1564798, 0.1564904, 
    0.1564908, 0.1564942, 0.1565034, 0.1564872, 0.156539, 0.1565066, 
    0.1564594, 0.1564689, 0.1564705, 0.1564668, 0.1564924, 0.1564831, 
    0.1565084, 0.1565015, 0.1565128, 0.1565072, 0.1565063, 0.1564992, 
    0.1564947, 0.1564835, 0.1564744, 0.1564673, 0.156469, 0.1564768, 
    0.1564911, 0.1565048, 0.1565018, 0.1565119, 0.1564854, 0.1564964, 
    0.1564921, 0.1565034, 0.1564789, 0.1564992, 0.1564736, 0.1564759, 
    0.1564829, 0.156497, 0.1565004, 0.1565037, 0.1565017, 0.1564915, 
    0.1564899, 0.1564828, 0.1564807, 0.1564754, 0.1564709, 0.156475, 
    0.1564792, 0.1564915, 0.1565026, 0.1565148, 0.1565179, 0.1565318, 
    0.1565202, 0.1565391, 0.1565228, 0.1565513, 0.1565007, 0.1565226, 
    0.1564833, 0.1564875, 0.156495, 0.1565127, 0.1565033, 0.1565144, 
    0.1564898, 0.156477, 0.1564738, 0.1564677, 0.156474, 0.1564735, 
    0.1564795, 0.1564776, 0.156492, 0.1564842, 0.1565063, 0.1565143, 
    0.1565374, 0.1565516, 0.1565663, 0.1565727, 0.1565747, 0.1565755,
  0.1697581, 0.1697711, 0.1697686, 0.1697791, 0.1697733, 0.1697801, 
    0.1697607, 0.1697716, 0.1697647, 0.1697593, 0.1697994, 0.1697796, 
    0.1698208, 0.1698079, 0.1698406, 0.1698187, 0.1698451, 0.1698401, 
    0.1698554, 0.169851, 0.1698704, 0.1698574, 0.1698808, 0.1698674, 
    0.1698694, 0.169857, 0.1697837, 0.1697969, 0.1697829, 0.1697848, 
    0.1697839, 0.1697734, 0.169768, 0.1697571, 0.1697591, 0.1697671, 
    0.1697856, 0.1697794, 0.1697953, 0.1697949, 0.1698127, 0.1698047, 
    0.1698348, 0.1698262, 0.1698512, 0.1698449, 0.1698509, 0.1698491, 
    0.1698509, 0.1698416, 0.1698456, 0.1698375, 0.1698061, 0.1698153, 
    0.1697881, 0.1697717, 0.1697612, 0.1697537, 0.1697547, 0.1697567, 
    0.1697672, 0.1697772, 0.1697848, 0.1697899, 0.1697949, 0.1698099, 
    0.1698181, 0.1698365, 0.1698333, 0.1698388, 0.1698443, 0.1698533, 
    0.1698518, 0.1698558, 0.1698387, 0.16985, 0.1698314, 0.1698365, 
    0.1697959, 0.1697811, 0.1697745, 0.169769, 0.1697555, 0.1697648, 
    0.1697612, 0.16977, 0.1697756, 0.1697728, 0.16979, 0.1697833, 0.1698186, 
    0.1698033, 0.1698436, 0.1698339, 0.169846, 0.1698398, 0.1698503, 
    0.1698409, 0.1698573, 0.1698608, 0.1698584, 0.1698679, 0.1698404, 
    0.1698508, 0.1697727, 0.1697732, 0.1697753, 0.169766, 0.1697654, 
    0.1697571, 0.1697646, 0.1697677, 0.1697759, 0.1697807, 0.1697854, 
    0.1697955, 0.1698068, 0.1698229, 0.1698346, 0.1698424, 0.1698376, 
    0.1698418, 0.1698371, 0.1698349, 0.1698595, 0.1698456, 0.1698665, 
    0.1698654, 0.1698559, 0.1698655, 0.1697735, 0.1697709, 0.1697619, 
    0.169769, 0.1697562, 0.1697633, 0.1697673, 0.1697833, 0.169787, 
    0.1697902, 0.1697967, 0.1698051, 0.1698198, 0.1698327, 0.1698446, 
    0.1698437, 0.169844, 0.1698466, 0.1698401, 0.1698477, 0.169849, 
    0.1698457, 0.1698652, 0.1698596, 0.1698654, 0.1698617, 0.1697718, 
    0.1697761, 0.1697738, 0.1697782, 0.1697751, 0.1697889, 0.1697931, 
    0.1698129, 0.1698049, 0.1698178, 0.1698062, 0.1698083, 0.1698181, 
    0.1698069, 0.1698319, 0.1698148, 0.1698467, 0.1698294, 0.1698478, 
    0.1698445, 0.16985, 0.1698549, 0.1698612, 0.1698727, 0.16987, 0.1698797, 
    0.1697827, 0.1697883, 0.1697879, 0.1697939, 0.1697983, 0.1698079, 
    0.1698235, 0.1698176, 0.1698284, 0.1698306, 0.1698142, 0.1698242, 
    0.1697922, 0.1697972, 0.1697943, 0.1697831, 0.1698189, 0.1698004, 
    0.1698347, 0.1698246, 0.1698542, 0.1698394, 0.1698686, 0.1698809, 
    0.169893, 0.1699068, 0.1697915, 0.1697876, 0.1697946, 0.1698041, 
    0.1698132, 0.1698252, 0.1698265, 0.1698288, 0.1698347, 0.1698396, 
    0.1698294, 0.1698408, 0.1697983, 0.1698205, 0.1697861, 0.1697963, 
    0.1698036, 0.1698005, 0.169817, 0.1698209, 0.1698367, 0.1698286, 
    0.1698778, 0.1698559, 0.1699175, 0.1699001, 0.1697863, 0.1697915, 
    0.1698097, 0.169801, 0.1698261, 0.1698323, 0.1698374, 0.1698438, 
    0.1698445, 0.1698483, 0.1698421, 0.1698481, 0.1698253, 0.1698354, 
    0.1698077, 0.1698144, 0.1698113, 0.1698079, 0.1698184, 0.1698295, 
    0.1698299, 0.1698334, 0.1698433, 0.1698262, 0.1698804, 0.1698466, 
    0.1697972, 0.1698072, 0.1698088, 0.1698049, 0.1698316, 0.1698219, 
    0.1698482, 0.1698411, 0.1698528, 0.169847, 0.1698461, 0.1698387, 
    0.169834, 0.1698223, 0.1698128, 0.1698055, 0.1698072, 0.1698153, 
    0.1698302, 0.1698445, 0.1698414, 0.169852, 0.1698243, 0.1698358, 
    0.1698313, 0.169843, 0.1698175, 0.1698388, 0.169812, 0.1698143, 
    0.1698217, 0.1698365, 0.1698399, 0.1698434, 0.1698413, 0.1698307, 
    0.169829, 0.1698215, 0.1698194, 0.1698138, 0.1698092, 0.1698134, 
    0.1698178, 0.1698307, 0.1698423, 0.169855, 0.1698582, 0.1698728, 
    0.1698607, 0.1698806, 0.1698635, 0.1698933, 0.1698403, 0.1698632, 
    0.1698221, 0.1698265, 0.1698344, 0.1698528, 0.169843, 0.1698546, 
    0.1698289, 0.1698155, 0.1698122, 0.1698059, 0.1698124, 0.1698119, 
    0.1698181, 0.1698161, 0.1698311, 0.1698231, 0.1698461, 0.1698545, 
    0.1698786, 0.1698935, 0.1699089, 0.1699157, 0.1699177, 0.1699186,
  0.1847913, 0.1848018, 0.1847998, 0.1848082, 0.1848036, 0.1848091, 
    0.1847935, 0.1848022, 0.1847966, 0.1847923, 0.1848248, 0.1848087, 
    0.184842, 0.1848315, 0.184858, 0.1848403, 0.1848617, 0.1848576, 0.18487, 
    0.1848665, 0.1848823, 0.1848717, 0.1848907, 0.1848798, 0.1848815, 
    0.1848713, 0.1848119, 0.1848227, 0.1848113, 0.1848128, 0.1848121, 
    0.1848036, 0.1847993, 0.1847905, 0.1847921, 0.1847986, 0.1848135, 
    0.1848085, 0.1848213, 0.184821, 0.1848354, 0.1848289, 0.1848533, 
    0.1848464, 0.1848666, 0.1848615, 0.1848664, 0.1848649, 0.1848664, 
    0.1848589, 0.1848621, 0.1848555, 0.1848301, 0.1848375, 0.1848155, 
    0.1848024, 0.1847938, 0.1847878, 0.1847886, 0.1847902, 0.1847987, 
    0.1848067, 0.1848128, 0.1848169, 0.184821, 0.1848332, 0.1848398, 
    0.1848547, 0.1848521, 0.1848566, 0.184861, 0.1848683, 0.1848671, 
    0.1848703, 0.1848565, 0.1848657, 0.1848505, 0.1848547, 0.1848219, 
    0.1848099, 0.1848046, 0.1848001, 0.1847893, 0.1847968, 0.1847938, 
    0.1848009, 0.1848054, 0.1848032, 0.184817, 0.1848116, 0.1848402, 
    0.1848278, 0.1848605, 0.1848526, 0.1848623, 0.1848574, 0.1848659, 
    0.1848582, 0.1848716, 0.1848745, 0.1848725, 0.1848802, 0.1848578, 
    0.1848663, 0.1848031, 0.1848035, 0.1848052, 0.1847977, 0.1847972, 
    0.1847905, 0.1847965, 0.1847991, 0.1848057, 0.1848096, 0.1848133, 
    0.1848215, 0.1848307, 0.1848437, 0.1848531, 0.1848595, 0.1848556, 
    0.184859, 0.1848552, 0.1848534, 0.1848734, 0.1848621, 0.1848791, 
    0.1848782, 0.1848704, 0.1848782, 0.1848037, 0.1848017, 0.1847944, 
    0.1848001, 0.1847897, 0.1847955, 0.1847988, 0.1848117, 0.1848146, 
    0.1848172, 0.1848225, 0.1848292, 0.1848411, 0.1848516, 0.1848612, 
    0.1848605, 0.1848608, 0.1848629, 0.1848576, 0.1848638, 0.1848648, 
    0.1848621, 0.184878, 0.1848735, 0.1848781, 0.1848752, 0.1848023, 
    0.1848059, 0.1848039, 0.1848075, 0.184805, 0.1848162, 0.1848196, 
    0.1848356, 0.1848291, 0.1848396, 0.1848302, 0.1848318, 0.1848398, 
    0.1848307, 0.184851, 0.1848371, 0.184863, 0.184849, 0.1848639, 0.1848612, 
    0.1848657, 0.1848697, 0.1848747, 0.1848841, 0.1848819, 0.1848898, 
    0.1848111, 0.1848157, 0.1848153, 0.1848202, 0.1848237, 0.1848316, 
    0.1848441, 0.1848394, 0.1848481, 0.1848499, 0.1848366, 0.1848447, 
    0.1848188, 0.1848229, 0.1848205, 0.1848115, 0.1848404, 0.1848255, 
    0.1848533, 0.1848451, 0.1848691, 0.1848571, 0.1848807, 0.1848909, 
    0.1849006, 0.1849119, 0.1848182, 0.1848151, 0.1848208, 0.1848285, 
    0.1848358, 0.1848456, 0.1848466, 0.1848484, 0.1848532, 0.1848572, 
    0.1848489, 0.1848582, 0.1848238, 0.1848418, 0.1848139, 0.1848222, 
    0.1848281, 0.1848255, 0.1848389, 0.184842, 0.1848549, 0.1848482, 
    0.1848883, 0.1848705, 0.1849207, 0.1849065, 0.184814, 0.1848183, 
    0.184833, 0.184826, 0.1848462, 0.1848512, 0.1848554, 0.1848606, 
    0.1848612, 0.1848643, 0.1848592, 0.1848641, 0.1848456, 0.1848538, 
    0.1848314, 0.1848368, 0.1848343, 0.1848315, 0.18484, 0.1848491, 
    0.1848493, 0.1848522, 0.1848603, 0.1848463, 0.1848905, 0.184863, 
    0.1848229, 0.184831, 0.1848322, 0.1848291, 0.1848507, 0.1848428, 
    0.1848642, 0.1848584, 0.1848679, 0.1848632, 0.1848625, 0.1848565, 
    0.1848527, 0.1848432, 0.1848355, 0.1848295, 0.1848309, 0.1848375, 
    0.1848496, 0.1848612, 0.1848587, 0.1848672, 0.1848448, 0.1848541, 
    0.1848505, 0.18486, 0.1848393, 0.1848567, 0.1848348, 0.1848367, 
    0.1848427, 0.1848547, 0.1848575, 0.1848603, 0.1848586, 0.18485, 
    0.1848486, 0.1848426, 0.1848409, 0.1848363, 0.1848325, 0.184836, 
    0.1848396, 0.18485, 0.1848594, 0.1848697, 0.1848723, 0.1848843, 
    0.1848744, 0.1848906, 0.1848767, 0.184901, 0.1848578, 0.1848764, 
    0.184843, 0.1848466, 0.184853, 0.184868, 0.1848599, 0.1848694, 0.1848485, 
    0.1848377, 0.184835, 0.1848299, 0.1848352, 0.1848347, 0.1848398, 
    0.1848382, 0.1848503, 0.1848438, 0.1848625, 0.1848693, 0.184889, 
    0.1849011, 0.1849136, 0.1849191, 0.1849208, 0.1849215,
  0.195208, 0.1952125, 0.1952117, 0.1952153, 0.1952133, 0.1952157, 0.1952089, 
    0.1952127, 0.1952103, 0.1952084, 0.1952224, 0.1952155, 0.1952299, 
    0.1952253, 0.1952368, 0.1952291, 0.1952384, 0.1952366, 0.195242, 
    0.1952404, 0.1952473, 0.1952427, 0.1952509, 0.1952462, 0.1952469, 
    0.1952425, 0.1952169, 0.1952216, 0.1952166, 0.1952173, 0.195217, 
    0.1952133, 0.1952115, 0.1952077, 0.1952084, 0.1952112, 0.1952176, 
    0.1952154, 0.1952209, 0.1952208, 0.195227, 0.1952242, 0.1952347, 
    0.1952317, 0.1952405, 0.1952383, 0.1952404, 0.1952398, 0.1952404, 
    0.1952371, 0.1952385, 0.1952357, 0.1952247, 0.1952279, 0.1952184, 
    0.1952128, 0.1952091, 0.1952065, 0.1952069, 0.1952076, 0.1952112, 
    0.1952146, 0.1952173, 0.195219, 0.1952208, 0.1952261, 0.1952289, 
    0.1952353, 0.1952342, 0.1952361, 0.1952381, 0.1952412, 0.1952407, 
    0.1952421, 0.1952361, 0.1952401, 0.1952335, 0.1952353, 0.1952212, 
    0.195216, 0.1952137, 0.1952118, 0.1952071, 0.1952104, 0.1952091, 
    0.1952121, 0.1952141, 0.1952131, 0.1952191, 0.1952168, 0.1952291, 
    0.1952237, 0.1952378, 0.1952344, 0.1952386, 0.1952365, 0.1952402, 
    0.1952369, 0.1952426, 0.1952439, 0.195243, 0.1952464, 0.1952367, 
    0.1952404, 0.1952131, 0.1952132, 0.195214, 0.1952108, 0.1952106, 
    0.1952077, 0.1952103, 0.1952114, 0.1952142, 0.1952159, 0.1952175, 
    0.195221, 0.195225, 0.1952306, 0.1952347, 0.1952374, 0.1952357, 
    0.1952372, 0.1952355, 0.1952348, 0.1952434, 0.1952385, 0.1952459, 
    0.1952455, 0.1952422, 0.1952455, 0.1952134, 0.1952125, 0.1952093, 
    0.1952118, 0.1952074, 0.1952098, 0.1952112, 0.1952168, 0.195218, 
    0.1952192, 0.1952214, 0.1952243, 0.1952295, 0.195234, 0.1952382, 
    0.1952379, 0.195238, 0.1952389, 0.1952366, 0.1952393, 0.1952397, 
    0.1952385, 0.1952454, 0.1952435, 0.1952455, 0.1952442, 0.1952128, 
    0.1952143, 0.1952135, 0.195215, 0.1952139, 0.1952187, 0.1952202, 
    0.1952271, 0.1952243, 0.1952288, 0.1952247, 0.1952254, 0.1952289, 
    0.195225, 0.1952337, 0.1952278, 0.1952389, 0.1952329, 0.1952393, 
    0.1952381, 0.1952401, 0.1952418, 0.195244, 0.1952481, 0.1952471, 
    0.1952506, 0.1952165, 0.1952185, 0.1952184, 0.1952204, 0.195222, 
    0.1952253, 0.1952308, 0.1952287, 0.1952325, 0.1952333, 0.1952275, 
    0.195231, 0.1952198, 0.1952216, 0.1952206, 0.1952167, 0.1952292, 
    0.1952227, 0.1952347, 0.1952312, 0.1952416, 0.1952364, 0.1952466, 
    0.195251, 0.1952553, 0.1952602, 0.1952196, 0.1952183, 0.1952207, 
    0.195224, 0.1952272, 0.1952314, 0.1952318, 0.1952326, 0.1952347, 
    0.1952364, 0.1952329, 0.1952368, 0.195222, 0.1952297, 0.1952177, 
    0.1952213, 0.1952238, 0.1952227, 0.1952285, 0.1952299, 0.1952354, 
    0.1952325, 0.1952499, 0.1952422, 0.195264, 0.1952578, 0.1952178, 
    0.1952196, 0.195226, 0.1952229, 0.1952317, 0.1952338, 0.1952356, 
    0.1952379, 0.1952381, 0.1952395, 0.1952373, 0.1952394, 0.1952314, 
    0.195235, 0.1952253, 0.1952276, 0.1952265, 0.1952253, 0.195229, 
    0.1952329, 0.195233, 0.1952343, 0.1952378, 0.1952317, 0.1952509, 
    0.1952389, 0.1952216, 0.1952251, 0.1952256, 0.1952243, 0.1952336, 
    0.1952302, 0.1952395, 0.195237, 0.1952411, 0.195239, 0.1952387, 
    0.1952361, 0.1952345, 0.1952304, 0.1952271, 0.1952245, 0.1952251, 
    0.1952279, 0.1952332, 0.1952382, 0.1952371, 0.1952408, 0.1952311, 
    0.1952351, 0.1952335, 0.1952376, 0.1952287, 0.1952362, 0.1952267, 
    0.1952276, 0.1952301, 0.1952353, 0.1952365, 0.1952378, 0.195237, 
    0.1952333, 0.1952327, 0.1952301, 0.1952294, 0.1952274, 0.1952258, 
    0.1952273, 0.1952288, 0.1952333, 0.1952374, 0.1952418, 0.195243, 
    0.1952482, 0.1952439, 0.195251, 0.1952449, 0.1952554, 0.1952367, 
    0.1952448, 0.1952303, 0.1952318, 0.1952346, 0.1952411, 0.1952376, 
    0.1952417, 0.1952327, 0.195228, 0.1952268, 0.1952246, 0.1952269, 
    0.1952267, 0.1952289, 0.1952282, 0.1952334, 0.1952306, 0.1952387, 
    0.1952417, 0.1952502, 0.1952555, 0.1952609, 0.1952633, 0.195264, 0.1952644,
  0.1982284, 0.1982291, 0.198229, 0.1982296, 0.1982292, 0.1982296, 0.1982286, 
    0.1982291, 0.1982288, 0.1982285, 0.1982307, 0.1982296, 0.1982318, 
    0.1982311, 0.1982329, 0.1982317, 0.1982332, 0.1982329, 0.1982337, 
    0.1982335, 0.1982346, 0.1982338, 0.1982351, 0.1982344, 0.1982345, 
    0.1982338, 0.1982298, 0.1982305, 0.1982297, 0.1982298, 0.1982298, 
    0.1982292, 0.198229, 0.1982284, 0.1982285, 0.1982289, 0.1982299, 
    0.1982296, 0.1982304, 0.1982304, 0.1982314, 0.1982309, 0.1982326, 
    0.1982321, 0.1982335, 0.1982331, 0.1982335, 0.1982334, 0.1982335, 
    0.198233, 0.1982332, 0.1982327, 0.198231, 0.1982315, 0.19823, 0.1982292, 
    0.1982286, 0.1982282, 0.1982282, 0.1982283, 0.1982289, 0.1982294, 
    0.1982298, 0.1982301, 0.1982304, 0.1982312, 0.1982317, 0.1982327, 
    0.1982325, 0.1982328, 0.1982331, 0.1982336, 0.1982335, 0.1982337, 
    0.1982328, 0.1982334, 0.1982324, 0.1982327, 0.1982305, 0.1982297, 
    0.1982293, 0.198229, 0.1982283, 0.1982288, 0.1982286, 0.1982291, 
    0.1982294, 0.1982292, 0.1982301, 0.1982298, 0.1982317, 0.1982309, 
    0.1982331, 0.1982325, 0.1982332, 0.1982329, 0.1982334, 0.1982329, 
    0.1982338, 0.198234, 0.1982339, 0.1982344, 0.1982329, 0.1982335, 
    0.1982292, 0.1982292, 0.1982293, 0.1982289, 0.1982288, 0.1982284, 
    0.1982288, 0.1982289, 0.1982294, 0.1982296, 0.1982299, 0.1982304, 
    0.1982311, 0.1982319, 0.1982326, 0.198233, 0.1982327, 0.198233, 
    0.1982327, 0.1982326, 0.1982339, 0.1982332, 0.1982343, 0.1982343, 
    0.1982338, 0.1982343, 0.1982293, 0.1982291, 0.1982286, 0.198229, 
    0.1982283, 0.1982287, 0.1982289, 0.1982298, 0.19823, 0.1982301, 
    0.1982305, 0.198231, 0.1982318, 0.1982325, 0.1982331, 0.1982331, 
    0.1982331, 0.1982332, 0.1982329, 0.1982333, 0.1982334, 0.1982332, 
    0.1982343, 0.198234, 0.1982343, 0.1982341, 0.1982291, 0.1982294, 
    0.1982293, 0.1982295, 0.1982293, 0.1982301, 0.1982303, 0.1982314, 
    0.198231, 0.1982317, 0.198231, 0.1982311, 0.1982317, 0.1982311, 
    0.1982324, 0.1982315, 0.1982332, 0.1982323, 0.1982333, 0.1982331, 
    0.1982334, 0.1982337, 0.198234, 0.1982347, 0.1982345, 0.1982351, 
    0.1982297, 0.19823, 0.19823, 0.1982303, 0.1982306, 0.1982311, 0.198232, 
    0.1982316, 0.1982322, 0.1982324, 0.1982315, 0.198232, 0.1982303, 
    0.1982305, 0.1982304, 0.1982298, 0.1982317, 0.1982307, 0.1982326, 
    0.198232, 0.1982337, 0.1982328, 0.1982345, 0.1982352, 0.1982358, 
    0.1982366, 0.1982302, 0.19823, 0.1982304, 0.1982309, 0.1982314, 
    0.1982321, 0.1982321, 0.1982322, 0.1982326, 0.1982328, 0.1982323, 
    0.1982329, 0.1982306, 0.1982318, 0.1982299, 0.1982305, 0.1982309, 
    0.1982307, 0.1982316, 0.1982318, 0.1982327, 0.1982322, 0.198235, 
    0.1982338, 0.1982372, 0.1982362, 0.1982299, 0.1982302, 0.1982312, 
    0.1982307, 0.1982321, 0.1982324, 0.1982327, 0.1982331, 0.1982331, 
    0.1982333, 0.198233, 0.1982333, 0.1982321, 0.1982326, 0.1982311, 
    0.1982315, 0.1982313, 0.1982311, 0.1982317, 0.1982323, 0.1982323, 
    0.1982325, 0.1982331, 0.1982321, 0.1982351, 0.1982332, 0.1982305, 
    0.1982311, 0.1982312, 0.1982309, 0.1982324, 0.1982319, 0.1982333, 
    0.1982329, 0.1982336, 0.1982333, 0.1982332, 0.1982328, 0.1982325, 
    0.1982319, 0.1982314, 0.198231, 0.1982311, 0.1982315, 0.1982323, 
    0.1982331, 0.1982329, 0.1982335, 0.198232, 0.1982326, 0.1982324, 
    0.198233, 0.1982316, 0.1982328, 0.1982313, 0.1982315, 0.1982319, 
    0.1982327, 0.1982329, 0.1982331, 0.1982329, 0.1982324, 0.1982323, 
    0.1982319, 0.1982317, 0.1982314, 0.1982312, 0.1982314, 0.1982317, 
    0.1982324, 0.198233, 0.1982337, 0.1982339, 0.1982347, 0.198234, 
    0.1982351, 0.1982342, 0.1982359, 0.1982329, 0.1982342, 0.1982319, 
    0.1982321, 0.1982326, 0.1982336, 0.198233, 0.1982337, 0.1982323, 
    0.1982315, 0.1982313, 0.198231, 0.1982314, 0.1982313, 0.1982317, 
    0.1982316, 0.1982324, 0.1982319, 0.1982332, 0.1982337, 0.198235, 
    0.1982359, 0.1982367, 0.1982371, 0.1982372, 0.1982373,
  0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 
    0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985142, 0.1985141, 
    0.1985143, 0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985144, 0.1985144, 0.1985144, 0.1985144, 0.1985145, 0.1985144, 
    0.1985144, 0.1985144, 0.1985142, 0.1985142, 0.1985141, 0.1985142, 
    0.1985142, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 
    0.1985142, 0.1985141, 0.1985142, 0.1985142, 0.1985142, 0.1985142, 
    0.1985143, 0.1985143, 0.1985144, 0.1985143, 0.1985144, 0.1985144, 
    0.1985144, 0.1985143, 0.1985143, 0.1985143, 0.1985142, 0.1985143, 
    0.1985142, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 
    0.1985141, 0.1985141, 0.1985142, 0.1985142, 0.1985142, 0.1985142, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985144, 
    0.1985144, 0.1985144, 0.1985143, 0.1985144, 0.1985143, 0.1985143, 
    0.1985142, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 
    0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985142, 0.1985142, 
    0.1985143, 0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985144, 0.1985143, 0.1985144, 0.1985144, 0.1985144, 0.1985144, 
    0.1985143, 0.1985144, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 
    0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 
    0.1985142, 0.1985142, 0.1985142, 0.1985143, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985144, 0.1985143, 
    0.1985144, 0.1985144, 0.1985144, 0.1985144, 0.1985141, 0.1985141, 
    0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985142, 
    0.1985142, 0.1985142, 0.1985142, 0.1985142, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985144, 
    0.1985144, 0.1985143, 0.1985144, 0.1985144, 0.1985144, 0.1985144, 
    0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985141, 0.1985142, 
    0.1985142, 0.1985143, 0.1985142, 0.1985143, 0.1985142, 0.1985142, 
    0.1985143, 0.1985142, 0.1985143, 0.1985143, 0.1985144, 0.1985143, 
    0.1985144, 0.1985143, 0.1985144, 0.1985144, 0.1985144, 0.1985144, 
    0.1985144, 0.1985145, 0.1985141, 0.1985142, 0.1985142, 0.1985142, 
    0.1985142, 0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985142, 0.1985142, 0.1985142, 0.1985142, 
    0.1985143, 0.1985142, 0.1985143, 0.1985143, 0.1985144, 0.1985143, 
    0.1985144, 0.1985145, 0.1985145, 0.1985146, 0.1985142, 0.1985142, 
    0.1985142, 0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985142, 0.1985143, 
    0.1985142, 0.1985142, 0.1985142, 0.1985142, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985144, 0.1985144, 0.1985146, 0.1985145, 
    0.1985142, 0.1985142, 0.1985142, 0.1985142, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985143, 0.1985144, 0.1985143, 0.1985144, 
    0.1985143, 0.1985143, 0.1985142, 0.1985143, 0.1985142, 0.1985142, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985145, 0.1985144, 0.1985142, 0.1985142, 0.1985142, 0.1985142, 
    0.1985143, 0.1985143, 0.1985144, 0.1985143, 0.1985144, 0.1985144, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985142, 0.1985142, 
    0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985144, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 0.1985144, 
    0.1985144, 0.1985144, 0.1985144, 0.1985145, 0.1985144, 0.1985145, 
    0.1985143, 0.1985144, 0.1985143, 0.1985143, 0.1985143, 0.1985144, 
    0.1985143, 0.1985144, 0.1985143, 0.1985143, 0.1985142, 0.1985142, 
    0.1985142, 0.1985142, 0.1985143, 0.1985143, 0.1985143, 0.1985143, 
    0.1985143, 0.1985144, 0.1985144, 0.1985145, 0.1985146, 0.1985146, 
    0.1985146, 0.1985146,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.605145, 8.605233, 8.605217, 8.605288, 8.605248, 8.605294, 8.605163, 
    8.605236, 8.60519, 8.605153, 8.605422, 8.60529, 8.605563, 8.60548, 
    8.605692, 8.60555, 8.605721, 8.60569, 8.605787, 8.60576, 8.605881, 
    8.6058, 8.605946, 8.605862, 8.605874, 8.605797, 8.605318, 8.605405, 
    8.605313, 8.605326, 8.60532, 8.605249, 8.605212, 8.605138, 8.605152, 
    8.605206, 8.60533, 8.60529, 8.605397, 8.605394, 8.605512, 8.605459, 
    8.605656, 8.6056, 8.605761, 8.605721, 8.605759, 8.605747, 8.605759, 
    8.6057, 8.605724, 8.605673, 8.605469, 8.605528, 8.605348, 8.605237, 
    8.605166, 8.605114, 8.605122, 8.605135, 8.605206, 8.605275, 8.605326, 
    8.60536, 8.605394, 8.605492, 8.605546, 8.605666, 8.605646, 8.605681, 
    8.605717, 8.605774, 8.605764, 8.605789, 8.605681, 8.605753, 8.605634, 
    8.605666, 8.605398, 8.605301, 8.605256, 8.60522, 8.605127, 8.605191, 
    8.605165, 8.605227, 8.605265, 8.605246, 8.605361, 8.605316, 8.605549, 
    8.60545, 8.605712, 8.60565, 8.605727, 8.605688, 8.605755, 8.605695, 
    8.605799, 8.605821, 8.605806, 8.605865, 8.605691, 8.605758, 8.605246, 
    8.605248, 8.605263, 8.605199, 8.605195, 8.605138, 8.605189, 8.60521, 
    8.605267, 8.605299, 8.60533, 8.605398, 8.605473, 8.605577, 8.605654, 
    8.605704, 8.605674, 8.6057, 8.605671, 8.605657, 8.605812, 8.605724, 
    8.605857, 8.60585, 8.60579, 8.605851, 8.60525, 8.605233, 8.605171, 
    8.60522, 8.605131, 8.605181, 8.605207, 8.605316, 8.605341, 8.605362, 
    8.605407, 8.605461, 8.605557, 8.605641, 8.605719, 8.605713, 8.605715, 
    8.605732, 8.60569, 8.605739, 8.605746, 8.605725, 8.605849, 8.605814, 
    8.60585, 8.605827, 8.605239, 8.605268, 8.605252, 8.605282, 8.605261, 
    8.605353, 8.605381, 8.605513, 8.60546, 8.605544, 8.605469, 8.605482, 
    8.605545, 8.605474, 8.605636, 8.605524, 8.605732, 8.605619, 8.60574, 
    8.605719, 8.605753, 8.605784, 8.605824, 8.605895, 8.605879, 8.605939, 
    8.605312, 8.60535, 8.605347, 8.605387, 8.605416, 8.60548, 8.605582, 
    8.605544, 8.605615, 8.605628, 8.605522, 8.605586, 8.605375, 8.605409, 
    8.60539, 8.605314, 8.605551, 8.60543, 8.605655, 8.60559, 8.60578, 
    8.605684, 8.605869, 8.605946, 8.606021, 8.606104, 8.605371, 8.605345, 
    8.605392, 8.605454, 8.605515, 8.605594, 8.605602, 8.605617, 8.605655, 
    8.605686, 8.60562, 8.605695, 8.605414, 8.605562, 8.605334, 8.605403, 
    8.605452, 8.605431, 8.605539, 8.605565, 8.605668, 8.605616, 8.605926, 
    8.605789, 8.60617, 8.606064, 8.605336, 8.605371, 8.605492, 8.605434, 
    8.605599, 8.605639, 8.605673, 8.605713, 8.605718, 8.605742, 8.605702, 
    8.605742, 8.605594, 8.605659, 8.605479, 8.605522, 8.605503, 8.60548, 
    8.605549, 8.605621, 8.605624, 8.605646, 8.605707, 8.6056, 8.605941, 
    8.605728, 8.60541, 8.605474, 8.605486, 8.60546, 8.605635, 8.605572, 
    8.605742, 8.605697, 8.605771, 8.605734, 8.605728, 8.60568, 8.605651, 
    8.605575, 8.605513, 8.605464, 8.605475, 8.605528, 8.605625, 8.605718, 
    8.605698, 8.605765, 8.605587, 8.605661, 8.605633, 8.605708, 8.605542, 
    8.60568, 8.605507, 8.605522, 8.60557, 8.605665, 8.605689, 8.605711, 
    8.605698, 8.605628, 8.605618, 8.60557, 8.605556, 8.605519, 8.605489, 
    8.605516, 8.605545, 8.605629, 8.605703, 8.605784, 8.605804, 8.605895, 
    8.60582, 8.605942, 8.605834, 8.606021, 8.60569, 8.605834, 8.605573, 
    8.605602, 8.605652, 8.60577, 8.605708, 8.605782, 8.605618, 8.60553, 
    8.605509, 8.605467, 8.60551, 8.605506, 8.605547, 8.605534, 8.605632, 
    8.605579, 8.605728, 8.605781, 8.605932, 8.606023, 8.606118, 8.606158, 
    8.606172, 8.606176 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  3.987384e-15, 3.987811e-15, 3.98773e-15, 3.98807e-15, 3.987884e-15, 
    3.988105e-15, 3.987474e-15, 3.987825e-15, 3.987603e-15, 3.987427e-15, 
    3.988724e-15, 3.988086e-15, 3.989421e-15, 3.989007e-15, 3.990058e-15, 
    3.989352e-15, 3.990202e-15, 3.990045e-15, 3.990536e-15, 3.990396e-15, 
    3.991008e-15, 3.990601e-15, 3.99134e-15, 3.990915e-15, 3.990979e-15, 
    3.990586e-15, 3.988222e-15, 3.988642e-15, 3.988195e-15, 3.988255e-15, 
    3.98823e-15, 3.987885e-15, 3.987707e-15, 3.987357e-15, 3.987422e-15, 
    3.987682e-15, 3.988283e-15, 3.988084e-15, 3.988601e-15, 3.98859e-15, 
    3.989162e-15, 3.988904e-15, 3.989875e-15, 3.9896e-15, 3.990401e-15, 
    3.990199e-15, 3.990391e-15, 3.990333e-15, 3.990391e-15, 3.990094e-15, 
    3.990221e-15, 3.989962e-15, 3.988951e-15, 3.989245e-15, 3.988365e-15, 
    3.987826e-15, 3.987488e-15, 3.987242e-15, 3.987277e-15, 3.987342e-15, 
    3.987683e-15, 3.988011e-15, 3.988259e-15, 3.988424e-15, 3.988588e-15, 
    3.989064e-15, 3.989334e-15, 3.989927e-15, 3.989826e-15, 3.990002e-15, 
    3.990179e-15, 3.990468e-15, 3.990421e-15, 3.990547e-15, 3.990002e-15, 
    3.990361e-15, 3.989767e-15, 3.989929e-15, 3.988607e-15, 3.988139e-15, 
    3.987918e-15, 3.987744e-15, 3.987303e-15, 3.987606e-15, 3.987486e-15, 
    3.987778e-15, 3.987959e-15, 3.987871e-15, 3.988429e-15, 3.988211e-15, 
    3.98935e-15, 3.988859e-15, 3.990158e-15, 3.989847e-15, 3.990233e-15, 
    3.990038e-15, 3.990371e-15, 3.990071e-15, 3.990595e-15, 3.990707e-15, 
    3.99063e-15, 3.990934e-15, 3.990054e-15, 3.990388e-15, 3.987867e-15, 
    3.987881e-15, 3.987951e-15, 3.987644e-15, 3.987627e-15, 3.987353e-15, 
    3.987599e-15, 3.987701e-15, 3.987972e-15, 3.988127e-15, 3.988277e-15, 
    3.988607e-15, 3.988971e-15, 3.98949e-15, 3.989867e-15, 3.990119e-15, 
    3.989966e-15, 3.990101e-15, 3.98995e-15, 3.98988e-15, 3.990664e-15, 
    3.990221e-15, 3.99089e-15, 3.990854e-15, 3.990548e-15, 3.990858e-15, 
    3.987892e-15, 3.987808e-15, 3.987511e-15, 3.987744e-15, 3.987324e-15, 
    3.987555e-15, 3.987687e-15, 3.988209e-15, 3.98833e-15, 3.988435e-15, 
    3.988647e-15, 3.988917e-15, 3.98939e-15, 3.989806e-15, 3.99019e-15, 
    3.990162e-15, 3.990172e-15, 3.990255e-15, 3.990045e-15, 3.99029e-15, 
    3.990329e-15, 3.990224e-15, 3.990849e-15, 3.99067e-15, 3.990853e-15, 
    3.990738e-15, 3.987836e-15, 3.987977e-15, 3.987901e-15, 3.988044e-15, 
    3.987941e-15, 3.988391e-15, 3.988526e-15, 3.989167e-15, 3.98891e-15, 
    3.989326e-15, 3.988955e-15, 3.989019e-15, 3.989329e-15, 3.988976e-15, 
    3.989778e-15, 3.989224e-15, 3.990258e-15, 3.989694e-15, 3.990293e-15, 
    3.990188e-15, 3.990365e-15, 3.99052e-15, 3.99072e-15, 3.991083e-15, 
    3.991e-15, 3.991308e-15, 3.988191e-15, 3.988372e-15, 3.988361e-15, 
    3.988554e-15, 3.988696e-15, 3.989011e-15, 3.98951e-15, 3.989324e-15, 
    3.989672e-15, 3.98974e-15, 3.989214e-15, 3.989532e-15, 3.988497e-15, 
    3.988659e-15, 3.988566e-15, 3.988202e-15, 3.98936e-15, 3.988762e-15, 
    3.989872e-15, 3.989548e-15, 3.990497e-15, 3.990019e-15, 3.990953e-15, 
    3.991341e-15, 3.99173e-15, 3.992158e-15, 3.988477e-15, 3.988352e-15, 
    3.988579e-15, 3.988883e-15, 3.98918e-15, 3.989567e-15, 3.98961e-15, 
    3.989681e-15, 3.989872e-15, 3.99003e-15, 3.989699e-15, 3.99007e-15, 
    3.988687e-15, 3.989414e-15, 3.988301e-15, 3.988629e-15, 3.988867e-15, 
    3.988768e-15, 3.989304e-15, 3.989429e-15, 3.989935e-15, 3.989676e-15, 
    3.991241e-15, 3.990546e-15, 3.992502e-15, 3.99195e-15, 3.988308e-15, 
    3.988478e-15, 3.989064e-15, 3.988786e-15, 3.989596e-15, 3.989793e-15, 
    3.989958e-15, 3.990162e-15, 3.990188e-15, 3.990309e-15, 3.99011e-15, 
    3.990303e-15, 3.989568e-15, 3.989897e-15, 3.989003e-15, 3.989217e-15, 
    3.98912e-15, 3.989011e-15, 3.989349e-15, 3.989703e-15, 3.989718e-15, 
    3.98983e-15, 3.990132e-15, 3.989599e-15, 3.991316e-15, 3.99024e-15, 
    3.988663e-15, 3.988981e-15, 3.989036e-15, 3.988911e-15, 3.989773e-15, 
    3.98946e-15, 3.990307e-15, 3.990079e-15, 3.990454e-15, 3.990267e-15, 
    3.990239e-15, 3.990001e-15, 3.98985e-15, 3.989472e-15, 3.989167e-15, 
    3.98893e-15, 3.988986e-15, 3.989247e-15, 3.989726e-15, 3.990186e-15, 
    3.990084e-15, 3.990426e-15, 3.989537e-15, 3.989905e-15, 3.98976e-15, 
    3.99014e-15, 3.989317e-15, 3.989993e-15, 3.989142e-15, 3.989218e-15, 
    3.989454e-15, 3.989925e-15, 3.990041e-15, 3.990151e-15, 3.990085e-15, 
    3.98974e-15, 3.989687e-15, 3.98945e-15, 3.98938e-15, 3.989202e-15, 
    3.989051e-15, 3.989187e-15, 3.989328e-15, 3.989743e-15, 3.990113e-15, 
    3.990521e-15, 3.990624e-15, 3.991082e-15, 3.990698e-15, 3.99132e-15, 
    3.990775e-15, 3.991729e-15, 3.990044e-15, 3.990775e-15, 3.989467e-15, 
    3.989609e-15, 3.989858e-15, 3.990448e-15, 3.990138e-15, 3.990505e-15, 
    3.989685e-15, 3.989252e-15, 3.98915e-15, 3.988943e-15, 3.989155e-15, 
    3.989138e-15, 3.98934e-15, 3.989275e-15, 3.989757e-15, 3.989499e-15, 
    3.990236e-15, 3.990504e-15, 3.991273e-15, 3.991741e-15, 3.992231e-15, 
    3.992444e-15, 3.992509e-15, 3.992536e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  9.826105, 9.873506, 9.864278, 9.902594, 9.881325, 9.906432, 9.835701, 
    9.875393, 9.850041, 9.830362, 9.977216, 9.904304, 10.05267, 10.00652, 
    10.1225, 10.0455, 10.13807, 10.12027, 10.17388, 10.1585, 10.22728, 
    10.18098, 10.26303, 10.21621, 10.22353, 10.17946, 9.918943, 9.968123, 
    9.916037, 9.923038, 9.919894, 9.881767, 9.862592, 9.822483, 9.829756, 
    9.859215, 9.926188, 9.903418, 9.96085, 9.959551, 10.02358, 9.99476, 
    10.10163, 10.07127, 10.15915, 10.137, 10.15811, 10.1517, 10.15819, 
    10.12573, 10.13963, 10.11109, 10.00018, 10.03286, 9.935034, 9.876332, 
    9.83744, 9.809905, 9.813795, 9.821215, 9.859387, 9.895354, 9.922818, 
    9.941216, 9.959364, 10.01444, 10.0432, 10.10778, 10.0961, 10.11589, 
    10.1348, 10.16662, 10.16138, 10.17541, 10.11536, 10.15525, 10.08945, 
    10.10742, 9.964327, 9.909556, 9.886354, 9.866053, 9.816787, 9.850794, 
    9.83738, 9.869306, 9.889627, 9.879572, 9.94172, 9.917532, 10.0449, 
    9.990187, 10.1326, 10.0985, 10.14078, 10.11919, 10.1562, 10.12289, 
    10.18063, 10.19324, 10.18462, 10.21772, 10.12104, 10.15811, 9.879292, 
    9.880932, 9.88857, 9.855022, 9.852971, 9.822285, 9.849584, 9.861225, 
    9.890804, 9.90833, 9.925007, 9.961731, 10.00285, 10.0598, 10.1007, 
    10.12818, 10.11133, 10.12621, 10.10957, 10.10178, 10.18851, 10.13976, 
    10.21296, 10.2089, 10.17574, 10.20936, 9.882083, 9.872649, 9.83995, 
    9.865535, 9.818946, 9.845011, 9.860019, 9.918042, 9.930812, 9.94267, 
    9.966108, 9.996241, 10.0487, 10.09423, 10.1359, 10.13285, 10.13392, 
    10.14325, 10.12016, 10.14704, 10.15156, 10.13975, 10.20835, 10.18873, 
    10.20881, 10.19603, 9.875714, 9.891592, 9.883011, 9.899152, 9.887781, 
    9.938412, 9.953623, 10.02482, 9.995648, 10.04191, 10.00038, 10.00781, 
    10.04343, 10.00265, 10.09173, 10.03141, 10.14361, 10.08321, 10.1474, 
    10.13572, 10.15506, 10.1724, 10.19424, 10.23462, 10.22526, 10.25907, 
    9.915288, 9.935937, 9.934113, 9.955744, 9.971761, 10.00652, 10.0617, 
    10.04098, 10.07904, 10.08669, 10.02887, 10.06435, 9.949767, 9.968356, 
    9.957282, 9.916919, 10.04576, 9.97975, 10.10138, 10.06576, 10.16993, 
    10.11805, 10.22011, 10.26394, 10.30526, 10.35371, 9.947212, 9.933169, 
    9.958317, 9.993182, 10.02541, 10.06793, 10.07229, 10.08027, 10.10095, 
    10.11837, 10.0828, 10.12273, 9.972681, 10.05145, 9.927868, 9.965163, 
    9.991123, 9.979725, 10.03861, 10.05239, 10.10852, 10.07948, 10.25312, 
    10.17608, 10.39067, 10.33044, 9.928267, 9.947161, 10.01309, 9.98169, 
    10.07077, 10.09265, 10.11045, 10.13325, 10.1357, 10.14922, 10.12708, 
    10.14835, 10.06802, 10.10387, 10.00554, 10.02953, 10.01855, 10.0064, 
    10.04367, 10.08336, 10.0842, 10.09694, 10.13293, 10.07113, 10.2631, 
    10.1443, 9.96779, 10.0043, 10.00951, 9.995357, 10.09046, 10.05604, 
    10.14889, 10.12375, 10.16497, 10.14447, 10.14146, 10.11518, 10.09883, 
    10.05762, 10.02416, 9.997408, 10.00366, 10.03294, 10.08579, 10.13593, 
    10.12494, 10.16183, 10.06433, 10.10515, 10.08937, 10.13056, 10.04043, 
    10.11717, 10.02087, 10.02929, 10.05536, 10.10793, 10.11957, 10.13202, 
    10.12434, 10.08713, 10.08104, 10.05472, 10.04747, 10.02746, 10.01085, 
    10.02603, 10.04193, 10.08714, 10.128, 10.17265, 10.18359, 10.23597, 
    10.19333, 10.26377, 10.20389, 10.30766, 10.12162, 10.20211, 10.05655, 
    10.07216, 10.10046, 10.16553, 10.13036, 10.17149, 10.0808, 10.03395, 
    10.02184, 9.999043, 10.02235, 10.02047, 10.04258, 10.03547, 10.08864, 
    10.06006, 10.14139, 10.17116, 10.25553, 10.30746, 10.36046, 10.38392, 
    10.39106, 10.39405 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  2.95167e-09, 2.915764e-09, 2.922662e-09, 2.894297e-09, 2.909949e-09, 
    2.891494e-09, 2.944304e-09, 2.91436e-09, 2.93339e-09, 2.948393e-09, 
    2.841078e-09, 2.893047e-09, 2.789385e-09, 2.820859e-09, 2.743332e-09, 
    2.794228e-09, 2.733332e-09, 2.744772e-09, 2.710681e-09, 2.720346e-09, 
    2.677801e-09, 2.706247e-09, 2.656354e-09, 2.684532e-09, 2.680077e-09, 
    2.707197e-09, 2.882407e-09, 2.847427e-09, 2.884512e-09, 2.879453e-09, 
    2.88172e-09, 2.909624e-09, 2.923933e-09, 2.954458e-09, 2.948859e-09, 
    2.926467e-09, 2.877185e-09, 2.89369e-09, 2.852518e-09, 2.853432e-09, 
    2.809163e-09, 2.828921e-09, 2.756884e-09, 2.776917e-09, 2.719941e-09, 
    2.73401e-09, 2.720598e-09, 2.724649e-09, 2.720545e-09, 2.741249e-09, 
    2.732333e-09, 2.750719e-09, 2.825195e-09, 2.802817e-09, 2.870836e-09, 
    2.913667e-09, 2.942975e-09, 2.964209e-09, 2.961185e-09, 2.95544e-09, 
    2.926337e-09, 2.899597e-09, 2.879608e-09, 2.866419e-09, 2.853564e-09, 
    2.815468e-09, 2.795788e-09, 2.752874e-09, 2.760505e-09, 2.747607e-09, 
    2.735419e-09, 2.715236e-09, 2.718535e-09, 2.709727e-09, 2.747947e-09, 
    2.722406e-09, 2.764874e-09, 2.753105e-09, 2.85009e-09, 2.889215e-09, 
    2.906236e-09, 2.921333e-09, 2.958864e-09, 2.932822e-09, 2.943022e-09, 
    2.918896e-09, 2.903811e-09, 2.911248e-09, 2.866061e-09, 2.883428e-09, 
    2.794632e-09, 2.832075e-09, 2.736834e-09, 2.758935e-09, 2.731599e-09, 
    2.745469e-09, 2.721803e-09, 2.74308e-09, 2.706467e-09, 2.698644e-09, 
    2.703984e-09, 2.683608e-09, 2.744271e-09, 2.720597e-09, 2.911457e-09, 
    2.910241e-09, 2.90459e-09, 2.929627e-09, 2.931176e-09, 2.954612e-09, 
    2.933736e-09, 2.924955e-09, 2.902942e-09, 2.890108e-09, 2.878032e-09, 
    2.851899e-09, 2.82337e-09, 2.784587e-09, 2.75749e-09, 2.739669e-09, 
    2.750565e-09, 2.74094e-09, 2.751704e-09, 2.756784e-09, 2.701569e-09, 
    2.73225e-09, 2.686517e-09, 2.689001e-09, 2.709518e-09, 2.688721e-09, 
    2.909388e-09, 2.916398e-09, 2.94106e-09, 2.921718e-09, 2.957191e-09, 
    2.937208e-09, 2.925864e-09, 2.883062e-09, 2.873858e-09, 2.865385e-09, 
    2.848825e-09, 2.827901e-09, 2.792059e-09, 2.761732e-09, 2.734714e-09, 
    2.736673e-09, 2.735983e-09, 2.730025e-09, 2.744839e-09, 2.727611e-09, 
    2.724743e-09, 2.732254e-09, 2.689334e-09, 2.701435e-09, 2.689054e-09, 
    2.696916e-09, 2.914115e-09, 2.902363e-09, 2.9087e-09, 2.896812e-09, 
    2.905175e-09, 2.868424e-09, 2.857621e-09, 2.808321e-09, 2.82831e-09, 
    2.796655e-09, 2.825056e-09, 2.819974e-09, 2.795634e-09, 2.823504e-09, 
    2.763382e-09, 2.803807e-09, 2.729794e-09, 2.769003e-09, 2.72738e-09, 
    2.73483e-09, 2.722522e-09, 2.711607e-09, 2.698021e-09, 2.673363e-09, 
    2.679027e-09, 2.658707e-09, 2.885053e-09, 2.870191e-09, 2.871492e-09, 
    2.856117e-09, 2.84487e-09, 2.820852e-09, 2.783311e-09, 2.797289e-09, 
    2.771753e-09, 2.766693e-09, 2.805539e-09, 2.781536e-09, 2.860346e-09, 
    2.847255e-09, 2.855033e-09, 2.883874e-09, 2.794052e-09, 2.839307e-09, 
    2.757047e-09, 2.780594e-09, 2.713156e-09, 2.746207e-09, 2.682156e-09, 
    2.655819e-09, 2.631584e-09, 2.603895e-09, 2.862157e-09, 2.872168e-09, 
    2.854301e-09, 2.830011e-09, 2.807908e-09, 2.779144e-09, 2.776241e-09, 
    2.770941e-09, 2.757327e-09, 2.746e-09, 2.76927e-09, 2.743178e-09, 
    2.844238e-09, 2.790204e-09, 2.875974e-09, 2.849494e-09, 2.831429e-09, 
    2.839321e-09, 2.798898e-09, 2.789567e-09, 2.752389e-09, 2.771462e-09, 
    2.662262e-09, 2.709312e-09, 2.583267e-09, 2.617102e-09, 2.875685e-09, 
    2.862191e-09, 2.816373e-09, 2.837955e-09, 2.777249e-09, 2.762771e-09, 
    2.751132e-09, 2.736418e-09, 2.734842e-09, 2.726223e-09, 2.74038e-09, 
    2.726779e-09, 2.779083e-09, 2.755421e-09, 2.821524e-09, 2.805091e-09, 
    2.812623e-09, 2.820939e-09, 2.795459e-09, 2.7689e-09, 2.76834e-09, 
    2.759953e-09, 2.736631e-09, 2.777009e-09, 2.656323e-09, 2.729361e-09, 
    2.847647e-09, 2.822377e-09, 2.818813e-09, 2.828509e-09, 2.764214e-09, 
    2.787109e-09, 2.726432e-09, 2.742524e-09, 2.716273e-09, 2.729244e-09, 
    2.731164e-09, 2.748066e-09, 2.758713e-09, 2.78605e-09, 2.808768e-09, 
    2.827098e-09, 2.822811e-09, 2.802763e-09, 2.767295e-09, 2.734698e-09, 
    2.741761e-09, 2.718248e-09, 2.781548e-09, 2.754586e-09, 2.764933e-09, 
    2.738144e-09, 2.797663e-09, 2.746784e-09, 2.811025e-09, 2.805252e-09, 
    2.787568e-09, 2.752778e-09, 2.745222e-09, 2.737203e-09, 2.742145e-09, 
    2.766408e-09, 2.770433e-09, 2.787996e-09, 2.79289e-09, 2.806507e-09, 
    2.817898e-09, 2.807485e-09, 2.796647e-09, 2.766399e-09, 2.739789e-09, 
    2.711452e-09, 2.704622e-09, 2.67255e-09, 2.698587e-09, 2.655928e-09, 
    2.692089e-09, 2.630202e-09, 2.743906e-09, 2.693175e-09, 2.786771e-09, 
    2.776321e-09, 2.757651e-09, 2.715925e-09, 2.738268e-09, 2.712181e-09, 
    2.770591e-09, 2.802076e-09, 2.810363e-09, 2.825975e-09, 2.810008e-09, 
    2.811299e-09, 2.796201e-09, 2.801032e-09, 2.765408e-09, 2.78441e-09, 
    2.731212e-09, 2.712385e-09, 2.660819e-09, 2.630317e-09, 2.600095e-09, 
    2.587006e-09, 2.583052e-09, 2.581404e-09 ;

 W_SCALAR =
  0.6251332, 0.6267919, 0.6264696, 0.6278064, 0.6270649, 0.6279401, 
    0.6254695, 0.6268578, 0.6259717, 0.6252825, 0.6303971, 0.627866, 
    0.6330203, 0.63141, 0.635451, 0.6327699, 0.6359908, 0.6353735, 0.63723, 
    0.6366984, 0.6390704, 0.6374753, 0.6402978, 0.6386895, 0.6389413, 
    0.6374227, 0.6283756, 0.6300823, 0.6282744, 0.6285179, 0.6284087, 
    0.6270803, 0.6264105, 0.6250061, 0.6252612, 0.6262925, 0.6286274, 
    0.6278352, 0.6298306, 0.6297855, 0.6320036, 0.631004, 0.6347262, 
    0.6336693, 0.6367207, 0.635954, 0.6366847, 0.6364631, 0.6366876, 
    0.635563, 0.636045, 0.6350549, 0.6311913, 0.6323281, 0.6289349, 
    0.6268905, 0.6255305, 0.6245646, 0.6247013, 0.6249616, 0.6262986, 
    0.6275542, 0.6285104, 0.6291496, 0.6297791, 0.6316831, 0.6326894, 
    0.6349398, 0.6345338, 0.6352214, 0.6358777, 0.636979, 0.6367977, 
    0.6372827, 0.6352032, 0.6365857, 0.6343026, 0.6349275, 0.6299508, 
    0.628049, 0.6272402, 0.6265315, 0.6248063, 0.625998, 0.6255283, 
    0.6266453, 0.6273546, 0.6270038, 0.6291671, 0.6283265, 0.632749, 
    0.6308459, 0.6358012, 0.6346171, 0.6360848, 0.6353361, 0.6366187, 
    0.6354644, 0.6374632, 0.637898, 0.6376008, 0.6387417, 0.6354004, 
    0.6366847, 0.626994, 0.6270512, 0.6273177, 0.6261459, 0.6260741, 
    0.6249992, 0.6259557, 0.6263629, 0.6273956, 0.6280063, 0.6285864, 
    0.6298611, 0.6312833, 0.6332693, 0.634694, 0.6356481, 0.6350631, 
    0.6355796, 0.6350022, 0.6347315, 0.6377351, 0.6360494, 0.6385776, 
    0.6384379, 0.6372943, 0.6384536, 0.6270913, 0.6267621, 0.6256183, 
    0.6265135, 0.624882, 0.6257956, 0.6263206, 0.6283442, 0.6287882, 0.6292, 
    0.6300128, 0.6310552, 0.6328818, 0.6344689, 0.6359159, 0.6358099, 
    0.6358472, 0.6361703, 0.6353699, 0.6363016, 0.636458, 0.6360492, 
    0.6384192, 0.6377425, 0.6384349, 0.6379943, 0.6268691, 0.627423, 
    0.6271238, 0.6276866, 0.6272901, 0.6290521, 0.6295799, 0.6320466, 
    0.6310347, 0.6326447, 0.6311983, 0.6314548, 0.6326974, 0.6312765, 
    0.6343815, 0.6322775, 0.6361828, 0.6340849, 0.6363142, 0.6359096, 
    0.6365793, 0.637179, 0.6379327, 0.6393225, 0.6390008, 0.6401621, 
    0.6282484, 0.6289662, 0.6289029, 0.6296536, 0.6302085, 0.6314103, 
    0.6333356, 0.6326119, 0.6339401, 0.6342066, 0.6321886, 0.6334281, 
    0.6294463, 0.6300905, 0.6297069, 0.6283051, 0.6327789, 0.6304849, 
    0.6347175, 0.6334772, 0.6370935, 0.6352965, 0.6388237, 0.6403288, 
    0.6417429, 0.643394, 0.6293576, 0.6288701, 0.6297428, 0.6309494, 
    0.6320676, 0.6335529, 0.6337047, 0.6339828, 0.6347026, 0.6353076, 
    0.6340708, 0.6354591, 0.6302401, 0.6329778, 0.6286859, 0.6299799, 
    0.6308783, 0.6304842, 0.6325291, 0.6330107, 0.6349657, 0.6339554, 
    0.6399575, 0.6373057, 0.6446492, 0.6426017, 0.6286998, 0.6293559, 
    0.631637, 0.6305522, 0.633652, 0.6344138, 0.6350328, 0.6358237, 0.635909, 
    0.6363773, 0.6356097, 0.6363469, 0.6335561, 0.634804, 0.6313763, 
    0.6322116, 0.6318274, 0.6314059, 0.6327062, 0.6340903, 0.6341197, 
    0.6345632, 0.6358125, 0.6336645, 0.6402997, 0.6362066, 0.630071, 
    0.6313334, 0.6315134, 0.6310247, 0.6343375, 0.6331382, 0.6363658, 
    0.6354943, 0.6369219, 0.6362127, 0.6361084, 0.6351968, 0.634629, 
    0.6331932, 0.6320238, 0.6310955, 0.6313114, 0.6323308, 0.6341749, 
    0.6359168, 0.6355354, 0.6368135, 0.6334274, 0.6348485, 0.6342995, 
    0.6357304, 0.6325927, 0.6352658, 0.6319087, 0.6322033, 0.6331143, 
    0.634945, 0.6353493, 0.6357813, 0.6355147, 0.6342216, 0.6340095, 
    0.6330922, 0.6328388, 0.6321391, 0.6315597, 0.6320892, 0.6326451, 
    0.6342221, 0.6356417, 0.6371875, 0.6375654, 0.639369, 0.6379012, 
    0.6403226, 0.6382647, 0.6418245, 0.6354202, 0.6382037, 0.6331557, 
    0.6337005, 0.6346855, 0.6369412, 0.6357237, 0.6371473, 0.6340013, 
    0.6323661, 0.6319425, 0.631152, 0.6319605, 0.6318948, 0.632668, 
    0.6324195, 0.6342744, 0.6332784, 0.6361058, 0.637136, 0.6400405, 
    0.6418176, 0.6436235, 0.64442, 0.6446623, 0.6447636,
  0.5461334, 0.5481776, 0.5477803, 0.549428, 0.5485141, 0.5495928, 0.5465479, 
    0.5482588, 0.5471667, 0.5463174, 0.5526217, 0.5495014, 0.5558565, 
    0.5538707, 0.5588548, 0.5555478, 0.5595208, 0.5587592, 0.5610498, 
    0.5603939, 0.5633209, 0.5613524, 0.5648358, 0.5628509, 0.5631616, 
    0.5612875, 0.5501296, 0.5522336, 0.5500049, 0.5503051, 0.5501704, 
    0.548533, 0.5477076, 0.5459769, 0.5462912, 0.5475622, 0.5504401, 
    0.5494635, 0.5519233, 0.5518678, 0.5546027, 0.5533701, 0.5579606, 
    0.556657, 0.5604212, 0.5594754, 0.5603769, 0.5601035, 0.5603804, 
    0.558993, 0.5595876, 0.5583661, 0.553601, 0.5550029, 0.550819, 0.5482991, 
    0.546623, 0.5454329, 0.5456012, 0.545922, 0.5475696, 0.5491171, 
    0.5502957, 0.5510837, 0.5518598, 0.5542075, 0.5554484, 0.5582242, 
    0.5577234, 0.5585716, 0.5593812, 0.56074, 0.5605164, 0.5611148, 
    0.5585491, 0.5602548, 0.5574381, 0.5582089, 0.5520715, 0.549727, 
    0.5487302, 0.5478567, 0.5457306, 0.5471991, 0.5466204, 0.5479969, 
    0.5488711, 0.5484387, 0.5511053, 0.550069, 0.555522, 0.5531752, 
    0.5592868, 0.5578262, 0.5596367, 0.558713, 0.5602955, 0.5588713, 
    0.5613374, 0.561874, 0.5615073, 0.5629152, 0.5587924, 0.5603769, 
    0.5484266, 0.5484971, 0.5488256, 0.5473815, 0.547293, 0.5459684, 
    0.547147, 0.5476488, 0.5489217, 0.5496743, 0.5503895, 0.5519609, 
    0.5537145, 0.5561636, 0.5579209, 0.5590979, 0.5583763, 0.5590134, 
    0.5583012, 0.5579672, 0.561673, 0.5595931, 0.5627128, 0.5625402, 
    0.5611291, 0.5625597, 0.5485467, 0.5481408, 0.5467313, 0.5478345, 
    0.545824, 0.5469497, 0.5475968, 0.5500909, 0.5506383, 0.5511459, 
    0.5521479, 0.5534332, 0.5556858, 0.5576433, 0.5594283, 0.5592976, 
    0.5593436, 0.5597422, 0.5587547, 0.5599043, 0.5600972, 0.5595928, 
    0.5625172, 0.5616822, 0.5625366, 0.5619929, 0.5482727, 0.5489555, 
    0.5485866, 0.5492803, 0.5487916, 0.5509636, 0.5516143, 0.5546558, 
    0.553408, 0.5553933, 0.5536097, 0.5539259, 0.5554583, 0.553706, 
    0.5575355, 0.5549404, 0.5597577, 0.5571697, 0.5599198, 0.5594206, 
    0.5602469, 0.5609868, 0.5619169, 0.5636321, 0.563235, 0.5646683, 
    0.5499728, 0.5508577, 0.5507796, 0.5517051, 0.5523893, 0.5538711, 
    0.5562454, 0.5553529, 0.556991, 0.5573197, 0.5548308, 0.5563595, 
    0.5514495, 0.5522438, 0.5517708, 0.5500427, 0.5555588, 0.5527301, 
    0.55795, 0.5564201, 0.5608813, 0.5586642, 0.5630165, 0.5648741, 
    0.5666198, 0.5686585, 0.5513402, 0.5507392, 0.5518151, 0.5533028, 
    0.5546817, 0.5565135, 0.5567007, 0.5570437, 0.5579316, 0.5586779, 
    0.5571523, 0.5588648, 0.5524282, 0.5558041, 0.5505121, 0.5521074, 
    0.553215, 0.5527291, 0.5552508, 0.5558447, 0.5582561, 0.5570099, 
    0.5644159, 0.5611432, 0.5702085, 0.5676802, 0.5505292, 0.5513381, 
    0.5541506, 0.5528129, 0.5566356, 0.5575754, 0.5583389, 0.5593146, 
    0.5594198, 0.5599976, 0.5590507, 0.5599601, 0.5565174, 0.5580567, 
    0.5538292, 0.5548592, 0.5543854, 0.5538656, 0.5554692, 0.5571763, 
    0.5572125, 0.5577596, 0.5593007, 0.5566511, 0.5648383, 0.559787, 
    0.5522197, 0.5537763, 0.5539982, 0.5533955, 0.5574812, 0.5560019, 
    0.5599835, 0.5589082, 0.5606696, 0.5597946, 0.5596658, 0.5585412, 
    0.5578408, 0.5560698, 0.5546275, 0.5534829, 0.5537491, 0.5550062, 
    0.5572806, 0.5594294, 0.5589589, 0.5605358, 0.5563587, 0.5581115, 
    0.5574344, 0.5591996, 0.5553293, 0.5586263, 0.5544856, 0.554849, 
    0.5559725, 0.5582306, 0.5587294, 0.5592623, 0.5589334, 0.5573383, 
    0.5570767, 0.5559452, 0.5556328, 0.5547699, 0.5540553, 0.5547082, 
    0.5553938, 0.5573388, 0.5590901, 0.5609973, 0.5614637, 0.5636894, 
    0.5618781, 0.5648664, 0.5623266, 0.5667205, 0.5588168, 0.5622514, 
    0.5560235, 0.5566955, 0.5579104, 0.5606934, 0.5591912, 0.5609477, 
    0.5570664, 0.5550497, 0.5545273, 0.5535526, 0.5545495, 0.5544685, 
    0.555422, 0.5551156, 0.5574034, 0.5561749, 0.5596626, 0.5609338, 
    0.5645183, 0.5667121, 0.568942, 0.5699255, 0.5702248, 0.5703499,
  0.5139211, 0.516171, 0.5157337, 0.5175475, 0.5165414, 0.517729, 0.5143773, 
    0.5162604, 0.5150583, 0.5141236, 0.5210646, 0.5176284, 0.5246286, 
    0.5224405, 0.5279334, 0.5242883, 0.5286677, 0.527828, 0.5303538, 
    0.5296305, 0.532859, 0.5306876, 0.5345306, 0.5323405, 0.5326833, 
    0.530616, 0.5183201, 0.5206372, 0.5181828, 0.5185133, 0.518365, 
    0.5165623, 0.5156536, 0.5137489, 0.5140947, 0.5154936, 0.5186619, 
    0.5175866, 0.5202954, 0.5202342, 0.523247, 0.521889, 0.5269477, 
    0.5255108, 0.5296607, 0.5286177, 0.5296118, 0.5293103, 0.5296156, 
    0.5280858, 0.5287414, 0.5273947, 0.5221434, 0.5236879, 0.5190792, 
    0.5163048, 0.5144599, 0.5131503, 0.5133355, 0.5136885, 0.5155017, 
    0.5172054, 0.518503, 0.5193707, 0.5202254, 0.5228116, 0.5241789, 
    0.5272383, 0.5266862, 0.5276212, 0.5285139, 0.5300122, 0.5297656, 
    0.5304255, 0.5275964, 0.5294771, 0.5263717, 0.5272214, 0.5204586, 
    0.5178767, 0.5167793, 0.5158178, 0.5134779, 0.515094, 0.514457, 
    0.5159721, 0.5169345, 0.5164585, 0.5193945, 0.5182534, 0.5242599, 
    0.5216743, 0.5284098, 0.5267995, 0.5287956, 0.5277772, 0.529522, 
    0.5279517, 0.5306711, 0.5312629, 0.5308585, 0.5324115, 0.5278647, 
    0.5296118, 0.5164452, 0.5165228, 0.5168844, 0.5152947, 0.5151973, 
    0.5137395, 0.5150366, 0.5155889, 0.5169901, 0.5178188, 0.5186062, 
    0.5203368, 0.5222684, 0.524967, 0.5269039, 0.5282016, 0.5274059, 
    0.5281084, 0.5273231, 0.5269549, 0.5310413, 0.5287476, 0.5321881, 
    0.5319979, 0.5304413, 0.5320193, 0.5165773, 0.5161306, 0.5145791, 
    0.5157933, 0.5135806, 0.5148195, 0.5155317, 0.5182775, 0.5188802, 
    0.5194392, 0.5205427, 0.5219585, 0.5244404, 0.5265979, 0.5285658, 
    0.5284216, 0.5284724, 0.5289119, 0.5278232, 0.5290906, 0.5293033, 
    0.5287472, 0.5319723, 0.5310513, 0.5319938, 0.5313941, 0.5162758, 
    0.5170274, 0.5166213, 0.5173849, 0.516847, 0.5192384, 0.519955, 
    0.5233055, 0.5219307, 0.5241181, 0.5221529, 0.5225013, 0.5241898, 
    0.5222591, 0.5264791, 0.5236191, 0.528929, 0.5260759, 0.5291077, 
    0.5285573, 0.5294684, 0.5302843, 0.5313102, 0.5332024, 0.5327643, 
    0.5343457, 0.5181475, 0.5191218, 0.5190359, 0.520055, 0.5208086, 
    0.5224409, 0.5250572, 0.5240736, 0.5258789, 0.5262412, 0.5234984, 
    0.5251829, 0.5197735, 0.5206484, 0.5201274, 0.5182244, 0.5243005, 
    0.521184, 0.5269359, 0.5252497, 0.5301681, 0.5277233, 0.5325232, 
    0.5345728, 0.5364995, 0.5387502, 0.5196532, 0.5189914, 0.5201762, 
    0.5218149, 0.523334, 0.5253526, 0.5255589, 0.525937, 0.5269157, 
    0.5277384, 0.5260566, 0.5279446, 0.5208515, 0.5245708, 0.5187413, 
    0.5204982, 0.5217182, 0.5211829, 0.5239611, 0.5246156, 0.5272735, 
    0.5258997, 0.5340672, 0.5304568, 0.540462, 0.5376701, 0.5187601, 
    0.5196508, 0.5227489, 0.5212753, 0.5254872, 0.5265231, 0.5273647, 
    0.5284404, 0.5285564, 0.5291935, 0.5281494, 0.5291522, 0.5253569, 
    0.5270536, 0.5223948, 0.5235295, 0.5230075, 0.5224349, 0.5242018, 
    0.5260832, 0.5261231, 0.5267261, 0.5284251, 0.5255042, 0.5345333, 
    0.5289613, 0.5206218, 0.5223365, 0.522581, 0.521917, 0.5264192, 
    0.5247888, 0.529178, 0.5279924, 0.5299346, 0.5289696, 0.5288277, 
    0.5275878, 0.5268155, 0.5248637, 0.5232744, 0.5220133, 0.5223066, 
    0.5236916, 0.5261981, 0.528567, 0.5280483, 0.529787, 0.525182, 0.5271141, 
    0.5263676, 0.5283136, 0.5240476, 0.5276815, 0.523118, 0.5235183, 
    0.5247564, 0.5272453, 0.5277952, 0.5283827, 0.5280201, 0.5262617, 
    0.5259734, 0.5247263, 0.524382, 0.5234312, 0.5226439, 0.5233632, 
    0.5241186, 0.5262623, 0.5281929, 0.530296, 0.5308103, 0.5332656, 
    0.5312674, 0.5345643, 0.5317621, 0.5366107, 0.5278916, 0.5316792, 
    0.5248126, 0.5255532, 0.5268924, 0.5299608, 0.5283044, 0.5302413, 
    0.5259621, 0.5237395, 0.5231639, 0.52209, 0.5231884, 0.5230991, 
    0.5241497, 0.5238121, 0.5263335, 0.5249794, 0.5288242, 0.5302259, 
    0.5341802, 0.5366014, 0.5390632, 0.5401495, 0.5404799, 0.5406181,
  0.50713, 0.5095204, 0.5090557, 0.5109833, 0.509914, 0.5111762, 0.5076146, 
    0.5096154, 0.5083381, 0.5073451, 0.5147234, 0.5110693, 0.5185162, 
    0.5161872, 0.5220361, 0.518154, 0.5228186, 0.5219238, 0.5246158, 
    0.5238447, 0.5272872, 0.5249716, 0.5290707, 0.5267342, 0.5270998, 
    0.5248953, 0.5118046, 0.5142686, 0.5116586, 0.51201, 0.5118523, 
    0.5099362, 0.5089706, 0.5069472, 0.5073145, 0.5088005, 0.512168, 
    0.5110249, 0.513905, 0.51384, 0.5170455, 0.5156004, 0.520986, 0.5194556, 
    0.5238768, 0.5227652, 0.5238246, 0.5235034, 0.5238289, 0.5221984, 
    0.5228971, 0.5214622, 0.5158711, 0.5175148, 0.5126117, 0.5096625, 
    0.5077024, 0.5063114, 0.5065081, 0.506883, 0.5088092, 0.5106196, 
    0.5119991, 0.5129217, 0.5138307, 0.5165821, 0.5180374, 0.5212955, 
    0.5207074, 0.5217035, 0.5226546, 0.5242515, 0.5239887, 0.5246922, 
    0.521677, 0.5236811, 0.5203725, 0.5212776, 0.5140787, 0.5113333, 
    0.5101668, 0.509145, 0.5066593, 0.508376, 0.5076993, 0.5093089, 
    0.5103317, 0.5098258, 0.512947, 0.5117337, 0.5181237, 0.5153719, 
    0.5225437, 0.5208281, 0.5229548, 0.5218696, 0.523729, 0.5220556, 
    0.524954, 0.525585, 0.5251538, 0.5268098, 0.5219628, 0.5238248, 
    0.5098117, 0.5098942, 0.5102785, 0.5085892, 0.5084858, 0.5069371, 
    0.508315, 0.5089018, 0.5103909, 0.5112717, 0.5121088, 0.5139492, 
    0.5160041, 0.5188765, 0.5209394, 0.5223218, 0.5214741, 0.5222225, 
    0.5213858, 0.5209936, 0.5253486, 0.5229036, 0.5265716, 0.5263687, 
    0.524709, 0.5263916, 0.5099521, 0.5094773, 0.507829, 0.509119, 0.5067685, 
    0.5080844, 0.508841, 0.5117593, 0.5124001, 0.5129945, 0.5141682, 
    0.5156744, 0.5183159, 0.5206133, 0.5227099, 0.5225563, 0.5226104, 
    0.5230787, 0.5219187, 0.5232692, 0.5234959, 0.5229032, 0.5263416, 
    0.5253594, 0.5263644, 0.5257249, 0.5096316, 0.5104305, 0.5099989, 
    0.5108105, 0.5102388, 0.512781, 0.5135431, 0.5171077, 0.5156448, 
    0.5179728, 0.5158812, 0.5162519, 0.5180491, 0.5159942, 0.5204868, 
    0.5174416, 0.523097, 0.5200573, 0.5232874, 0.5227008, 0.5236719, 
    0.5245416, 0.5256354, 0.5276535, 0.5271862, 0.5288734, 0.5116211, 
    0.512657, 0.5125656, 0.5136495, 0.514451, 0.5161877, 0.5189726, 
    0.5179254, 0.5198476, 0.5202335, 0.5173131, 0.5191064, 0.5133501, 
    0.5142806, 0.5137264, 0.5117029, 0.518167, 0.5148503, 0.5209734, 
    0.5191775, 0.5244176, 0.5218123, 0.526929, 0.5291157, 0.5311723, 
    0.533576, 0.5132221, 0.5125183, 0.5137783, 0.5155215, 0.5171381, 
    0.5192871, 0.5195069, 0.5199094, 0.5209519, 0.5218283, 0.5200368, 
    0.5220479, 0.5144966, 0.5184547, 0.5122524, 0.5141208, 0.5154187, 
    0.5148492, 0.5178057, 0.5185024, 0.521333, 0.5198697, 0.5285762, 
    0.5247256, 0.535405, 0.5324223, 0.5122724, 0.5132196, 0.5165154, 
    0.5149474, 0.5194305, 0.5205336, 0.5214301, 0.5225763, 0.5226999, 
    0.5233789, 0.5222663, 0.5233349, 0.5192917, 0.5210987, 0.5161386, 
    0.5173463, 0.5167906, 0.5161813, 0.5180618, 0.5200651, 0.5201076, 
    0.5207499, 0.52256, 0.5194486, 0.5290736, 0.5231314, 0.5142523, 
    0.5160766, 0.5163367, 0.5156302, 0.5204231, 0.5186868, 0.5233623, 
    0.5220989, 0.5241688, 0.5231403, 0.522989, 0.5216678, 0.5208452, 
    0.5187665, 0.5170746, 0.5157326, 0.5160447, 0.5175188, 0.5201876, 
    0.5227112, 0.5221585, 0.5240115, 0.5191055, 0.5211632, 0.520368, 
    0.5224411, 0.5178976, 0.5217677, 0.5169082, 0.5173343, 0.5186523, 
    0.5213029, 0.5218888, 0.5225148, 0.5221285, 0.5202553, 0.5199482, 
    0.5186203, 0.5182537, 0.5172415, 0.5164036, 0.5171692, 0.5179733, 
    0.5202559, 0.5223125, 0.524554, 0.5251024, 0.527721, 0.5255898, 
    0.5291067, 0.5261173, 0.5312911, 0.5219915, 0.5260288, 0.5187122, 
    0.5195007, 0.520927, 0.5241967, 0.5224314, 0.5244957, 0.5199361, 
    0.5175697, 0.516957, 0.5158143, 0.5169832, 0.5168881, 0.5180064, 
    0.517647, 0.5203317, 0.5188897, 0.5229853, 0.5244793, 0.5286967, 
    0.5312811, 0.5339104, 0.535071, 0.5354242, 0.5355718,
  0.5311532, 0.5336223, 0.5331421, 0.5351346, 0.5340291, 0.5353341, 
    0.5316536, 0.5337204, 0.5324008, 0.5313753, 0.5390045, 0.5352235, 
    0.5429347, 0.5405207, 0.5465874, 0.5425591, 0.5474001, 0.5464708, 
    0.5492676, 0.5484662, 0.5520464, 0.5496376, 0.5539031, 0.5514708, 
    0.5518513, 0.5495582, 0.5359839, 0.5385336, 0.5358329, 0.5361964, 
    0.5360332, 0.5340521, 0.5330542, 0.5309644, 0.5313436, 0.5328785, 
    0.5363598, 0.5351776, 0.5381573, 0.53809, 0.5414101, 0.5399128, 
    0.5454971, 0.5439091, 0.5484996, 0.5473447, 0.5484455, 0.5481116, 
    0.5484498, 0.546756, 0.5474817, 0.5459915, 0.5401932, 0.5418965, 
    0.5368188, 0.5337692, 0.5317442, 0.5303081, 0.5305111, 0.5308982, 
    0.5328875, 0.5347585, 0.536185, 0.5371396, 0.5380803, 0.5409299, 
    0.5424383, 0.5458184, 0.545208, 0.5462421, 0.5472298, 0.5488891, 
    0.5486159, 0.5493472, 0.5462146, 0.5482963, 0.5448604, 0.5457999, 
    0.538337, 0.5354964, 0.5342904, 0.5332345, 0.5306672, 0.53244, 0.5317411, 
    0.5334038, 0.5344608, 0.533938, 0.5371657, 0.5359106, 0.5425277, 
    0.5396761, 0.5471146, 0.5453333, 0.5475416, 0.5464146, 0.548346, 
    0.5466077, 0.5496193, 0.5502754, 0.549827, 0.5515496, 0.5465114, 
    0.5484455, 0.5339234, 0.5340087, 0.5344059, 0.5326602, 0.5325534, 
    0.530954, 0.532377, 0.5329832, 0.5345221, 0.5354328, 0.5362986, 
    0.5382029, 0.540331, 0.5433084, 0.5454487, 0.5468841, 0.5460038, 
    0.546781, 0.5459123, 0.5455051, 0.5500296, 0.5474885, 0.5513018, 
    0.5510906, 0.5493646, 0.5511144, 0.5340685, 0.5335779, 0.531875, 
    0.5332076, 0.5307799, 0.5321387, 0.5329203, 0.535937, 0.5365999, 
    0.5372149, 0.5384297, 0.5399894, 0.542727, 0.5451103, 0.5472872, 
    0.5471277, 0.5471839, 0.5476704, 0.5464655, 0.5478683, 0.5481038, 
    0.547488, 0.5510623, 0.5500408, 0.5510861, 0.5504209, 0.5337373, 
    0.534563, 0.5341168, 0.5349559, 0.5343648, 0.536994, 0.5377826, 
    0.5414746, 0.5399587, 0.5423713, 0.5402037, 0.5405877, 0.5424504, 
    0.5403207, 0.5449791, 0.5418206, 0.5476893, 0.5445334, 0.5478872, 
    0.5472778, 0.5482867, 0.5491906, 0.5503279, 0.5524275, 0.5519412, 
    0.5536976, 0.5357941, 0.5368657, 0.5367711, 0.5378927, 0.5387225, 
    0.5405212, 0.543408, 0.5423222, 0.5443158, 0.5447161, 0.5416874, 
    0.5435469, 0.5375829, 0.538546, 0.5379724, 0.5358787, 0.5425726, 
    0.5391359, 0.5454841, 0.5436206, 0.5490617, 0.546355, 0.5516735, 0.55395, 
    0.5560928, 0.5585996, 0.5374504, 0.5367222, 0.5380261, 0.539831, 
    0.5415061, 0.5437343, 0.5439622, 0.5443799, 0.5454617, 0.5463716, 
    0.5445122, 0.5465997, 0.5387697, 0.5428709, 0.536447, 0.5383806, 
    0.5397246, 0.5391347, 0.542198, 0.5429204, 0.5458574, 0.5443388, 
    0.5533881, 0.5493818, 0.5605088, 0.5573961, 0.5364679, 0.5374479, 
    0.5408608, 0.5392365, 0.543883, 0.5450276, 0.5459582, 0.5471485, 
    0.5472769, 0.5479822, 0.5468264, 0.5479365, 0.543739, 0.5456142, 
    0.5404703, 0.5417218, 0.541146, 0.5405145, 0.5424636, 0.5445414, 
    0.5445856, 0.5452521, 0.5471315, 0.5439018, 0.553906, 0.5477251, 
    0.5385168, 0.540406, 0.5406756, 0.5399437, 0.5449129, 0.5431117, 
    0.547965, 0.5466527, 0.5488031, 0.5477344, 0.5475771, 0.546205, 0.545351, 
    0.5431943, 0.5414402, 0.5400498, 0.540373, 0.5419006, 0.5446685, 
    0.5472886, 0.5467145, 0.5486396, 0.5435459, 0.5456811, 0.5448558, 
    0.5470081, 0.5422934, 0.5463087, 0.5412678, 0.5417094, 0.5430759, 
    0.5458262, 0.5464345, 0.5470846, 0.5466834, 0.5447388, 0.5444201, 
    0.5430426, 0.5426625, 0.5416133, 0.5407449, 0.5415384, 0.5423718, 
    0.5447394, 0.5468745, 0.5492035, 0.5497736, 0.5524977, 0.5502804, 
    0.5539405, 0.5508291, 0.5562165, 0.5465411, 0.5507371, 0.543138, 
    0.5439559, 0.545436, 0.5488321, 0.546998, 0.5491429, 0.5444076, 
    0.5419534, 0.5413184, 0.5401344, 0.5413455, 0.541247, 0.5424061, 
    0.5420336, 0.5448181, 0.5433221, 0.5475733, 0.5491259, 0.5535136, 
    0.5562061, 0.5589485, 0.56016, 0.5605288, 0.5606831,
  0.535265, 0.5381082, 0.5375549, 0.5398521, 0.5385771, 0.5400822, 0.5358407, 
    0.5382213, 0.536701, 0.5355206, 0.544323, 0.5399546, 0.5488767, 
    0.5460782, 0.5531207, 0.5484409, 0.5540666, 0.5529851, 0.5562425, 
    0.5553083, 0.5594857, 0.5566739, 0.5616568, 0.5588133, 0.5592578, 
    0.5565813, 0.5408322, 0.5437784, 0.5406579, 0.5410775, 0.5408891, 
    0.5386035, 0.5374536, 0.5350478, 0.5354841, 0.5372512, 0.5412662, 
    0.5399016, 0.5433432, 0.5432654, 0.5471087, 0.5453743, 0.5518528, 
    0.5500077, 0.5553473, 0.5540021, 0.5552841, 0.5548952, 0.5552892, 
    0.553317, 0.5541616, 0.5524276, 0.5456989, 0.5476725, 0.5417963, 
    0.5382774, 0.5359451, 0.534293, 0.5345265, 0.5349716, 0.5372615, 
    0.5394182, 0.5410644, 0.5421669, 0.5432542, 0.5465522, 0.5483008, 
    0.5522264, 0.5515167, 0.552719, 0.5538684, 0.5558012, 0.5554827, 
    0.5563352, 0.552687, 0.5551104, 0.5511127, 0.5522047, 0.543551, 
    0.5402696, 0.5388784, 0.5376613, 0.5347059, 0.5367461, 0.5359415, 
    0.5378564, 0.5390749, 0.5384721, 0.5421971, 0.5407476, 0.5484046, 
    0.5451003, 0.5537342, 0.5516623, 0.5542314, 0.5529197, 0.5551683, 
    0.5531443, 0.5566525, 0.5574179, 0.5568948, 0.5589053, 0.5530323, 
    0.5552842, 0.5384552, 0.5385535, 0.5390115, 0.5369997, 0.5368767, 
    0.5350358, 0.5366736, 0.5373718, 0.5391455, 0.5401961, 0.5411955, 
    0.543396, 0.5458585, 0.5493103, 0.5517965, 0.553466, 0.552442, 0.553346, 
    0.5523354, 0.551862, 0.5571311, 0.5541695, 0.5586159, 0.5583694, 
    0.5563555, 0.5583972, 0.5386226, 0.538057, 0.5360956, 0.5376303, 
    0.5348356, 0.5363992, 0.5372993, 0.540778, 0.5415435, 0.542254, 
    0.5436582, 0.545463, 0.5486357, 0.5514032, 0.5539352, 0.5537495, 
    0.5538149, 0.5543814, 0.5529789, 0.5546118, 0.5548862, 0.5541691, 
    0.5583364, 0.5571442, 0.5583642, 0.5575877, 0.5382407, 0.5391927, 
    0.5386782, 0.5396459, 0.5389642, 0.5419987, 0.54291, 0.5471834, 
    0.5454274, 0.548223, 0.545711, 0.5461558, 0.5483148, 0.5458466, 
    0.5512506, 0.5475845, 0.5544034, 0.5507327, 0.5546339, 0.5539243, 
    0.5550992, 0.5561526, 0.5574791, 0.5599312, 0.5593628, 0.5614164, 
    0.5406131, 0.5418504, 0.5417413, 0.5430373, 0.5439968, 0.5460787, 
    0.549426, 0.5481661, 0.5504799, 0.550945, 0.5474301, 0.5495871, 
    0.5426791, 0.5437927, 0.5431294, 0.5407107, 0.5484566, 0.5444751, 
    0.5518376, 0.5496728, 0.5560024, 0.5528504, 0.5590501, 0.5617115, 
    0.5642214, 0.5671629, 0.5425261, 0.5416847, 0.5431915, 0.5452796, 
    0.5472199, 0.5498047, 0.5500694, 0.5505545, 0.5518116, 0.5528697, 
    0.5507081, 0.5531351, 0.5440515, 0.5488027, 0.541367, 0.5436014, 
    0.5451564, 0.5444738, 0.5480222, 0.5488601, 0.5522715, 0.5505067, 
    0.5610543, 0.5563756, 0.5694073, 0.5657498, 0.541391, 0.5425231, 
    0.5464721, 0.5445915, 0.5499774, 0.551307, 0.5523889, 0.5537737, 
    0.5539231, 0.5547445, 0.5533989, 0.5546913, 0.5498102, 0.5519888, 
    0.5460199, 0.54747, 0.5468026, 0.5460711, 0.5483302, 0.5507421, 
    0.5507933, 0.5515679, 0.553754, 0.5499992, 0.5616602, 0.554445, 
    0.5437589, 0.5459454, 0.5462576, 0.54541, 0.5511737, 0.549082, 0.5547245, 
    0.5531967, 0.5557009, 0.5544558, 0.5542728, 0.5526759, 0.5516829, 
    0.5491779, 0.5471436, 0.5455329, 0.5459072, 0.5476773, 0.5508897, 
    0.5539368, 0.5532687, 0.5555104, 0.549586, 0.5520666, 0.5511073, 
    0.5536103, 0.5481327, 0.5527965, 0.5469437, 0.5474557, 0.5490406, 
    0.5522353, 0.5529429, 0.5536994, 0.5532324, 0.5509713, 0.5506012, 
    0.5490019, 0.5485609, 0.5473441, 0.5463379, 0.5472573, 0.5482237, 
    0.5509722, 0.5534548, 0.5561677, 0.5568324, 0.5600132, 0.5574237, 
    0.5617006, 0.558064, 0.5643664, 0.5530668, 0.5579566, 0.5491126, 
    0.550062, 0.5517816, 0.5557347, 0.5535985, 0.556097, 0.5505866, 
    0.5477386, 0.5470024, 0.5456308, 0.5470338, 0.5469196, 0.5482635, 
    0.5478315, 0.5510635, 0.5493262, 0.5542683, 0.5560772, 0.5612011, 
    0.5643542, 0.5675728, 0.568997, 0.5694308, 0.5696123,
  0.5840983, 0.5875093, 0.5868445, 0.589608, 0.5880732, 0.5898854, 0.584788, 
    0.5876453, 0.5858195, 0.5844043, 0.5950121, 0.5897316, 0.6005515, 
    0.5971429, 0.6057478, 0.6000199, 0.6069103, 0.6055813, 0.6095911, 
    0.6084391, 0.6136036, 0.6101237, 0.6163011, 0.6127701, 0.613321, 
    0.6100094, 0.5907898, 0.5943519, 0.5905796, 0.5910859, 0.5908585, 
    0.588105, 0.5867228, 0.5838382, 0.5843607, 0.5864798, 0.5913137, 
    0.5896677, 0.5938249, 0.5937306, 0.5983964, 0.5962877, 0.6041918, 
    0.6019331, 0.6084871, 0.6068311, 0.6084093, 0.6079302, 0.6084155, 
    0.6059889, 0.6070272, 0.6048968, 0.596682, 0.5990831, 0.5919539, 
    0.5877128, 0.5849131, 0.5829352, 0.5832143, 0.583747, 0.5864922, 
    0.5890854, 0.5910701, 0.5924017, 0.5937171, 0.5977193, 0.599849, 0.60465, 
    0.60378, 0.6052545, 0.6066666, 0.6090466, 0.6086541, 0.6097055, 
    0.6052153, 0.6081952, 0.6032851, 0.6046234, 0.5940765, 0.5901113, 
    0.5884356, 0.5869722, 0.5834292, 0.5858736, 0.5849087, 0.5872067, 
    0.5886721, 0.5879468, 0.5924382, 0.5906877, 0.5999755, 0.595955, 
    0.6065017, 0.6039584, 0.6071131, 0.6055008, 0.6082666, 0.6057768, 
    0.6100972, 0.611043, 0.6103966, 0.6128841, 0.6056391, 0.6084094, 
    0.5879266, 0.5880448, 0.5885958, 0.5861779, 0.5860302, 0.583824, 
    0.5857866, 0.5866246, 0.5887571, 0.5900226, 0.5912283, 0.5938888, 
    0.5968758, 0.601081, 0.6041229, 0.606172, 0.6049144, 0.6060246, 
    0.6047838, 0.6042032, 0.6106886, 0.6070369, 0.6125255, 0.6122202, 
    0.6097306, 0.6122546, 0.5881278, 0.5874478, 0.5850935, 0.586935, 
    0.5835842, 0.5854575, 0.5865376, 0.5907245, 0.5916485, 0.592507, 
    0.5942064, 0.5963954, 0.6002575, 0.6036409, 0.6067488, 0.6065204, 
    0.6066008, 0.6072976, 0.6055735, 0.6075812, 0.607919, 0.6070364, 
    0.6121793, 0.6107047, 0.6122137, 0.611253, 0.5876687, 0.5888139, 
    0.5881948, 0.5893596, 0.5885388, 0.5921984, 0.5933005, 0.5984874, 
    0.5963523, 0.5997542, 0.5966967, 0.5972373, 0.599866, 0.5968614, 
    0.6034541, 0.5989759, 0.6073247, 0.60282, 0.6076084, 0.6067353, 
    0.6081815, 0.6094803, 0.6111187, 0.6141564, 0.6134512, 0.616002, 
    0.5905255, 0.5920193, 0.5918874, 0.5934545, 0.5946166, 0.5971436, 
    0.6012223, 0.5996847, 0.6025106, 0.6030799, 0.5987878, 0.6014192, 
    0.5930212, 0.5943693, 0.5935661, 0.5906433, 0.6000389, 0.5951965, 
    0.6041734, 0.6015237, 0.6092949, 0.6054158, 0.6130636, 0.6163694, 
    0.6194996, 0.6231846, 0.5928361, 0.5918191, 0.5936412, 0.5961727, 
    0.5985318, 0.601685, 0.6020085, 0.6026018, 0.6041414, 0.6054395, 
    0.6027898, 0.6057654, 0.5946829, 0.6004613, 0.5914353, 0.5941375, 
    0.5960231, 0.5951949, 0.5995092, 0.6005313, 0.6047055, 0.6025434, 
    0.6155517, 0.6097554, 0.6260084, 0.6214122, 0.5914643, 0.5928324, 
    0.5976219, 0.5953377, 0.601896, 0.6035231, 0.6048494, 0.6065502, 
    0.6067339, 0.6077446, 0.6060895, 0.6076791, 0.6016917, 0.6043587, 
    0.597072, 0.5988364, 0.5980239, 0.5971342, 0.5998847, 0.6028314, 
    0.6028942, 0.6038428, 0.6065259, 0.6019228, 0.6163054, 0.6073759, 
    0.5943283, 0.5969815, 0.597361, 0.5963311, 0.6033598, 0.6008022, 
    0.6077199, 0.605841, 0.608923, 0.6073893, 0.607164, 0.6052015, 0.6039836, 
    0.6009192, 0.598439, 0.5964803, 0.5969351, 0.5990889, 0.6030121, 
    0.6067508, 0.6059296, 0.6086882, 0.6014177, 0.6044541, 0.6032786, 
    0.6063493, 0.599644, 0.6053496, 0.5981957, 0.598819, 0.6007515, 0.604661, 
    0.6055293, 0.6064588, 0.605885, 0.603112, 0.602659, 0.6007044, 0.6001662, 
    0.5986832, 0.5974587, 0.5985774, 0.5997549, 0.6031131, 0.6061582, 
    0.6094989, 0.6103196, 0.6142582, 0.6110502, 0.6163557, 0.6118423, 
    0.6196809, 0.6056816, 0.6117094, 0.6008395, 0.6019995, 0.6041046, 
    0.6089647, 0.6063348, 0.6094117, 0.6026412, 0.5991636, 0.5982671, 
    0.5965992, 0.5983052, 0.5981663, 0.5998035, 0.5992768, 0.6032249, 
    0.6011004, 0.6071585, 0.6093872, 0.6157342, 0.6196657, 0.6236995, 
    0.6254914, 0.6260381, 0.6262668,
  0.6622252, 0.667787, 0.6666976, 0.671243, 0.6687129, 0.6717016, 0.6633443, 
    0.6680101, 0.6650232, 0.6627214, 0.6802661, 0.6714472, 0.6897115, 
    0.6838751, 0.6987643, 0.6887959, 0.7008166, 0.6984711, 0.7055877, 
    0.7035307, 0.7128337, 0.7065421, 0.7177787, 0.711318, 0.7123192, 
    0.706337, 0.6732006, 0.679154, 0.6728517, 0.6736924, 0.6733148, 
    0.6687651, 0.6664985, 0.6618038, 0.6626507, 0.6661011, 0.6740713, 
    0.6713416, 0.6782681, 0.6781098, 0.6860123, 0.682423, 0.6960332, 
    0.6920996, 0.7036162, 0.7006762, 0.7034776, 0.7026251, 0.7034886, 
    0.699189, 0.7010233, 0.6972685, 0.6830921, 0.6871875, 0.6751375, 
    0.6681209, 0.6635476, 0.6603438, 0.6607947, 0.6616563, 0.6661214, 
    0.6703799, 0.6736662, 0.6758848, 0.6780871, 0.6848565, 0.6885021, 
    0.6968355, 0.6953132, 0.6978964, 0.7003853, 0.7046142, 0.7039137, 
    0.7057924, 0.6978276, 0.7030964, 0.6944497, 0.696789, 0.6786907, 
    0.6720755, 0.6693091, 0.6669068, 0.6611419, 0.6651114, 0.6635405, 
    0.6672909, 0.6696985, 0.6685053, 0.6759458, 0.6730312, 0.6887196, 
    0.6818596, 0.7000939, 0.6956249, 0.7011755, 0.6983296, 0.7032234, 
    0.6988153, 0.7064946, 0.7081949, 0.707032, 0.7115249, 0.698573, 
    0.7034777, 0.6684719, 0.6686662, 0.6695728, 0.665608, 0.665367, 
    0.6617808, 0.6649696, 0.6663378, 0.6698385, 0.6719288, 0.6739293, 
    0.6783754, 0.6834213, 0.6906251, 0.6959125, 0.6995119, 0.6972994, 
    0.6992519, 0.6970701, 0.6960531, 0.7075568, 0.7010406, 0.7108743, 
    0.710321, 0.7058374, 0.7103833, 0.6688027, 0.6676859, 0.6638409, 
    0.6668459, 0.6613927, 0.6644334, 0.6661956, 0.6730922, 0.6746284, 
    0.6760606, 0.6789091, 0.6826057, 0.6892048, 0.6950704, 0.7005307, 
    0.7001271, 0.7002692, 0.7015024, 0.6984575, 0.7020053, 0.7026053, 
    0.7010396, 0.710247, 0.7075859, 0.7103093, 0.7085733, 0.6680484, 
    0.6699321, 0.6689128, 0.6708325, 0.669479, 0.6755454, 0.6773885, 
    0.6861679, 0.6825326, 0.6883391, 0.683117, 0.6840357, 0.6885313, 
    0.6833967, 0.6947443, 0.6870039, 0.7015504, 0.6936398, 0.7020535, 
    0.7005069, 0.703072, 0.7053893, 0.7083312, 0.7138421, 0.7125562, 
    0.7172273, 0.672762, 0.6752465, 0.6750266, 0.6776467, 0.6795995, 
    0.6838763, 0.6908692, 0.6882198, 0.6931019, 0.6940922, 0.6866818, 
    0.6912096, 0.6769206, 0.6791832, 0.6778337, 0.6729575, 0.6888288, 
    0.6805774, 0.6960008, 0.6913906, 0.7050578, 0.69818, 0.711851, 0.7179045, 
    0.723722, 0.7306815, 0.6766108, 0.6749128, 0.6779597, 0.6822283, 
    0.6862439, 0.6916698, 0.6922305, 0.6932604, 0.695945, 0.6982218, 
    0.6935872, 0.6987953, 0.6797112, 0.6895559, 0.6742736, 0.6787934, 
    0.6819748, 0.6805746, 0.6879184, 0.6896765, 0.6969328, 0.6931588, 
    0.7163987, 0.7058818, 0.7360995, 0.7273188, 0.6743218, 0.6766047, 
    0.6846906, 0.6808157, 0.6920354, 0.6948649, 0.6971852, 0.7001796, 
    0.7005044, 0.7022955, 0.6993665, 0.702179, 0.6916814, 0.6963253, 
    0.6837546, 0.6867649, 0.685376, 0.6838605, 0.6885636, 0.6936597, 
    0.6937689, 0.6954229, 0.7001367, 0.6920817, 0.7177866, 0.7016412, 
    0.6791143, 0.6836007, 0.6842464, 0.6824967, 0.69458, 0.6901437, 
    0.7022516, 0.6989285, 0.7043935, 0.7016649, 0.7012656, 0.6978035, 
    0.6956691, 0.6903458, 0.6860851, 0.6827497, 0.6835219, 0.6871975, 
    0.6939742, 0.7005342, 0.6990845, 0.7039745, 0.6912072, 0.6964923, 
    0.6944383, 0.6998249, 0.6881499, 0.6980637, 0.6856694, 0.686735, 
    0.6900563, 0.6968548, 0.6983797, 0.7000182, 0.6990059, 0.6941482, 
    0.6933598, 0.689975, 0.6890477, 0.6865026, 0.6844125, 0.6863218, 
    0.6883404, 0.69415, 0.6994877, 0.7054225, 0.7068936, 0.7140281, 
    0.7082078, 0.7178793, 0.7096372, 0.7240615, 0.6986477, 0.709397, 
    0.6902081, 0.6922148, 0.6958807, 0.7044679, 0.6997993, 0.7052665, 
    0.6933289, 0.6873255, 0.6857913, 0.6829515, 0.6858565, 0.6856192, 
    0.6884239, 0.6875196, 0.6943448, 0.6906587, 0.7012558, 0.7052227, 
    0.7167343, 0.7240329, 0.731664, 0.7351019, 0.7361569, 0.7365991,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.535556e-11, 3.551315e-11, 3.548243e-11, 3.560961e-11, 3.553903e-11, 
    3.562224e-11, 3.538733e-11, 3.551913e-11, 3.543493e-11, 3.536944e-11, 
    3.585634e-11, 3.561499e-11, 3.610765e-11, 3.595332e-11, 3.634116e-11, 
    3.60835e-11, 3.639314e-11, 3.633368e-11, 3.651264e-11, 3.646129e-11, 
    3.669025e-11, 3.653622e-11, 3.680911e-11, 3.665342e-11, 3.667769e-11, 
    3.653094e-11, 3.566385e-11, 3.582654e-11, 3.565413e-11, 3.567733e-11, 
    3.566689e-11, 3.55403e-11, 3.547653e-11, 3.53432e-11, 3.536735e-11, 
    3.546526e-11, 3.568748e-11, 3.561197e-11, 3.580226e-11, 3.579797e-11, 
    3.601002e-11, 3.591435e-11, 3.627134e-11, 3.616973e-11, 3.646339e-11, 
    3.638941e-11, 3.645983e-11, 3.643841e-11, 3.645999e-11, 3.635162e-11, 
    3.639796e-11, 3.630264e-11, 3.593271e-11, 3.604151e-11, 3.571702e-11, 
    3.552212e-11, 3.539293e-11, 3.530133e-11, 3.53142e-11, 3.533888e-11, 
    3.546576e-11, 3.558518e-11, 3.567627e-11, 3.573718e-11, 3.579724e-11, 
    3.597917e-11, 3.607563e-11, 3.629177e-11, 3.625276e-11, 3.63188e-11, 
    3.638202e-11, 3.648812e-11, 3.647064e-11, 3.651735e-11, 3.631688e-11, 
    3.645004e-11, 3.62302e-11, 3.629028e-11, 3.581378e-11, 3.56325e-11, 
    3.555537e-11, 3.548798e-11, 3.532412e-11, 3.543722e-11, 3.539257e-11, 
    3.549868e-11, 3.556613e-11, 3.553271e-11, 3.573881e-11, 3.565857e-11, 
    3.608128e-11, 3.589905e-11, 3.637469e-11, 3.626068e-11, 3.640191e-11, 
    3.632982e-11, 3.645328e-11, 3.63421e-11, 3.65347e-11, 3.657668e-11, 
    3.65479e-11, 3.665819e-11, 3.633569e-11, 3.645942e-11, 3.553199e-11, 
    3.553744e-11, 3.556276e-11, 3.545121e-11, 3.544439e-11, 3.53423e-11, 
    3.543305e-11, 3.547173e-11, 3.556996e-11, 3.562802e-11, 3.568327e-11, 
    3.580492e-11, 3.594081e-11, 3.613111e-11, 3.626802e-11, 3.63598e-11, 
    3.630347e-11, 3.635313e-11, 3.629753e-11, 3.627144e-11, 3.656082e-11, 
    3.639823e-11, 3.664221e-11, 3.662871e-11, 3.651815e-11, 3.663012e-11, 
    3.554118e-11, 3.550981e-11, 3.540109e-11, 3.54861e-11, 3.533112e-11, 
    3.54178e-11, 3.54676e-11, 3.566015e-11, 3.57025e-11, 3.574178e-11, 
    3.581935e-11, 3.591894e-11, 3.60939e-11, 3.624626e-11, 3.638555e-11, 
    3.637528e-11, 3.637886e-11, 3.640991e-11, 3.633281e-11, 3.642249e-11, 
    3.643749e-11, 3.639813e-11, 3.662679e-11, 3.656142e-11, 3.662827e-11, 
    3.658564e-11, 3.551996e-11, 3.557259e-11, 3.554406e-11, 3.559762e-11, 
    3.555979e-11, 3.572766e-11, 3.577797e-11, 3.601385e-11, 3.591697e-11, 
    3.607116e-11, 3.593257e-11, 3.59571e-11, 3.607598e-11, 3.593996e-11, 
    3.62377e-11, 3.603563e-11, 3.641108e-11, 3.620899e-11, 3.642366e-11, 
    3.638463e-11, 3.644913e-11, 3.650696e-11, 3.657967e-11, 3.671403e-11, 
    3.668283e-11, 3.67953e-11, 3.565116e-11, 3.57195e-11, 3.57135e-11, 
    3.578508e-11, 3.583802e-11, 3.5953e-11, 3.613749e-11, 3.606802e-11, 
    3.619546e-11, 3.622106e-11, 3.602732e-11, 3.614617e-11, 3.576493e-11, 
    3.582635e-11, 3.578975e-11, 3.565595e-11, 3.608364e-11, 3.58639e-11, 
    3.626981e-11, 3.615057e-11, 3.649859e-11, 3.632537e-11, 3.666567e-11, 
    3.681131e-11, 3.694861e-11, 3.710898e-11, 3.575685e-11, 3.571029e-11, 
    3.579353e-11, 3.590879e-11, 3.601583e-11, 3.61583e-11, 3.617285e-11, 
    3.619949e-11, 3.626865e-11, 3.632686e-11, 3.62078e-11, 3.634134e-11, 
    3.58405e-11, 3.610273e-11, 3.569217e-11, 3.581563e-11, 3.590147e-11, 
    3.586382e-11, 3.605959e-11, 3.610572e-11, 3.629344e-11, 3.619637e-11, 
    3.677521e-11, 3.651883e-11, 3.723129e-11, 3.703185e-11, 3.569399e-11, 
    3.575654e-11, 3.597452e-11, 3.587075e-11, 3.616772e-11, 3.624092e-11, 
    3.630039e-11, 3.63765e-11, 3.638466e-11, 3.642978e-11, 3.635577e-11, 
    3.64268e-11, 3.615818e-11, 3.627814e-11, 3.59492e-11, 3.60291e-11, 
    3.599231e-11, 3.595189e-11, 3.607643e-11, 3.620923e-11, 3.621208e-11, 
    3.625461e-11, 3.637457e-11, 3.616821e-11, 3.680807e-11, 3.641244e-11, 
    3.582479e-11, 3.594536e-11, 3.596261e-11, 3.591587e-11, 3.623346e-11, 
    3.611829e-11, 3.642868e-11, 3.634467e-11, 3.648221e-11, 3.641383e-11, 
    3.640368e-11, 3.631592e-11, 3.626119e-11, 3.612325e-11, 3.601102e-11, 
    3.59222e-11, 3.594277e-11, 3.604038e-11, 3.621725e-11, 3.63849e-11, 
    3.63481e-11, 3.647126e-11, 3.614537e-11, 3.62819e-11, 3.622901e-11, 
    3.636674e-11, 3.6066e-11, 3.632258e-11, 3.600042e-11, 3.602859e-11, 
    3.611589e-11, 3.629171e-11, 3.633064e-11, 3.63722e-11, 3.634648e-11, 
    3.622205e-11, 3.620165e-11, 3.611352e-11, 3.608913e-11, 3.60221e-11, 
    3.596651e-11, 3.601722e-11, 3.607038e-11, 3.622182e-11, 3.635832e-11, 
    3.650729e-11, 3.654379e-11, 3.671791e-11, 3.657601e-11, 3.681007e-11, 
    3.661086e-11, 3.695583e-11, 3.633744e-11, 3.660592e-11, 3.611989e-11, 
    3.617213e-11, 3.626669e-11, 3.648388e-11, 3.636657e-11, 3.650375e-11, 
    3.620083e-11, 3.604378e-11, 3.600321e-11, 3.592753e-11, 3.600486e-11, 
    3.599858e-11, 3.607264e-11, 3.604876e-11, 3.622674e-11, 3.61311e-11, 
    3.64029e-11, 3.650222e-11, 3.678303e-11, 3.695535e-11, 3.713106e-11, 
    3.72086e-11, 3.723222e-11, 3.724205e-11,
  1.796106e-11, 1.809839e-11, 1.807167e-11, 1.818266e-11, 1.812107e-11, 
    1.819378e-11, 1.798888e-11, 1.810384e-11, 1.803043e-11, 1.797343e-11, 
    1.839876e-11, 1.818762e-11, 1.861919e-11, 1.848379e-11, 1.882469e-11, 
    1.859808e-11, 1.887051e-11, 1.881817e-11, 1.897595e-11, 1.89307e-11, 
    1.9133e-11, 1.899685e-11, 1.923823e-11, 1.910047e-11, 1.912198e-11, 
    1.899236e-11, 1.823006e-11, 1.837241e-11, 1.822163e-11, 1.82419e-11, 
    1.823281e-11, 1.812233e-11, 1.806674e-11, 1.79506e-11, 1.797167e-11, 
    1.805699e-11, 1.825102e-11, 1.818509e-11, 1.83515e-11, 1.834773e-11, 
    1.853366e-11, 1.844974e-11, 1.876333e-11, 1.8674e-11, 1.893259e-11, 
    1.886743e-11, 1.892952e-11, 1.891069e-11, 1.892977e-11, 1.883423e-11, 
    1.887514e-11, 1.879117e-11, 1.846544e-11, 1.856093e-11, 1.827667e-11, 
    1.810652e-11, 1.799392e-11, 1.791416e-11, 1.792543e-11, 1.794691e-11, 
    1.805749e-11, 1.816172e-11, 1.82413e-11, 1.829461e-11, 1.834719e-11, 
    1.850664e-11, 1.859132e-11, 1.878139e-11, 1.874706e-11, 1.880526e-11, 
    1.886095e-11, 1.895456e-11, 1.893915e-11, 1.898042e-11, 1.880374e-11, 
    1.892109e-11, 1.872751e-11, 1.878038e-11, 1.83614e-11, 1.820287e-11, 
    1.813556e-11, 1.80768e-11, 1.793409e-11, 1.803259e-11, 1.799373e-11, 
    1.808625e-11, 1.814513e-11, 1.811601e-11, 1.829607e-11, 1.822598e-11, 
    1.859634e-11, 1.843646e-11, 1.885445e-11, 1.875411e-11, 1.887853e-11, 
    1.881501e-11, 1.89239e-11, 1.882589e-11, 1.89958e-11, 1.903287e-11, 
    1.900754e-11, 1.910495e-11, 1.882046e-11, 1.892951e-11, 1.811518e-11, 
    1.811993e-11, 1.814207e-11, 1.804484e-11, 1.80389e-11, 1.795002e-11, 
    1.802911e-11, 1.806282e-11, 1.814855e-11, 1.819931e-11, 1.824763e-11, 
    1.835404e-11, 1.847314e-11, 1.864021e-11, 1.876061e-11, 1.884147e-11, 
    1.879188e-11, 1.883566e-11, 1.878671e-11, 1.876379e-11, 1.901897e-11, 
    1.887552e-11, 1.909093e-11, 1.907899e-11, 1.89814e-11, 1.908033e-11, 
    1.812327e-11, 1.809595e-11, 1.800119e-11, 1.807533e-11, 1.794035e-11, 
    1.801585e-11, 1.80593e-11, 1.822742e-11, 1.826446e-11, 1.829881e-11, 
    1.836673e-11, 1.845403e-11, 1.860756e-11, 1.874154e-11, 1.88642e-11, 
    1.88552e-11, 1.885837e-11, 1.888579e-11, 1.881787e-11, 1.889696e-11, 
    1.891023e-11, 1.887551e-11, 1.907739e-11, 1.901963e-11, 1.907874e-11, 
    1.904112e-11, 1.810483e-11, 1.815082e-11, 1.812596e-11, 1.817271e-11, 
    1.813976e-11, 1.828643e-11, 1.833049e-11, 1.853724e-11, 1.84523e-11, 
    1.858757e-11, 1.846603e-11, 1.848754e-11, 1.859195e-11, 1.84726e-11, 
    1.873413e-11, 1.855663e-11, 1.888686e-11, 1.870902e-11, 1.889802e-11, 
    1.886366e-11, 1.892058e-11, 1.897159e-11, 1.903586e-11, 1.915463e-11, 
    1.91271e-11, 1.92266e-11, 1.821948e-11, 1.827928e-11, 1.827403e-11, 
    1.83367e-11, 1.838309e-11, 1.848383e-11, 1.864582e-11, 1.858485e-11, 
    1.869687e-11, 1.871938e-11, 1.854923e-11, 1.865361e-11, 1.831936e-11, 
    1.837318e-11, 1.834114e-11, 1.822418e-11, 1.859887e-11, 1.84062e-11, 
    1.876259e-11, 1.865778e-11, 1.896431e-11, 1.881161e-11, 1.911196e-11, 
    1.924084e-11, 1.936253e-11, 1.950499e-11, 1.831197e-11, 1.82713e-11, 
    1.834416e-11, 1.844512e-11, 1.853904e-11, 1.866416e-11, 1.867699e-11, 
    1.870046e-11, 1.876135e-11, 1.881259e-11, 1.870787e-11, 1.882544e-11, 
    1.838564e-11, 1.861564e-11, 1.825591e-11, 1.836392e-11, 1.843917e-11, 
    1.840617e-11, 1.857789e-11, 1.861845e-11, 1.878359e-11, 1.869816e-11, 
    1.920899e-11, 1.898234e-11, 1.961379e-11, 1.943654e-11, 1.825709e-11, 
    1.831184e-11, 1.850284e-11, 1.841187e-11, 1.867253e-11, 1.87369e-11, 
    1.878931e-11, 1.885635e-11, 1.886361e-11, 1.890338e-11, 1.883822e-11, 
    1.890081e-11, 1.866443e-11, 1.876992e-11, 1.848099e-11, 1.855114e-11, 
    1.851887e-11, 1.848347e-11, 1.85928e-11, 1.870951e-11, 1.871204e-11, 
    1.874952e-11, 1.885524e-11, 1.867359e-11, 1.923825e-11, 1.888874e-11, 
    1.83716e-11, 1.847733e-11, 1.849248e-11, 1.845148e-11, 1.873044e-11, 
    1.862918e-11, 1.890241e-11, 1.882842e-11, 1.894972e-11, 1.888941e-11, 
    1.888054e-11, 1.88032e-11, 1.875511e-11, 1.863381e-11, 1.853535e-11, 
    1.845743e-11, 1.847554e-11, 1.856117e-11, 1.871667e-11, 1.886425e-11, 
    1.883188e-11, 1.894049e-11, 1.865359e-11, 1.877367e-11, 1.872721e-11, 
    1.884845e-11, 1.858323e-11, 1.88089e-11, 1.85257e-11, 1.855047e-11, 
    1.862717e-11, 1.878181e-11, 1.881613e-11, 1.885275e-11, 1.883015e-11, 
    1.872063e-11, 1.870272e-11, 1.862531e-11, 1.860394e-11, 1.854508e-11, 
    1.849638e-11, 1.854086e-11, 1.858762e-11, 1.872069e-11, 1.88409e-11, 
    1.897231e-11, 1.900453e-11, 1.915852e-11, 1.903309e-11, 1.92402e-11, 
    1.906401e-11, 1.936943e-11, 1.882205e-11, 1.905889e-11, 1.863067e-11, 
    1.867663e-11, 1.875985e-11, 1.895129e-11, 1.884788e-11, 1.896886e-11, 
    1.870202e-11, 1.856411e-11, 1.852853e-11, 1.846216e-11, 1.853005e-11, 
    1.852453e-11, 1.858957e-11, 1.856866e-11, 1.872511e-11, 1.864101e-11, 
    1.888031e-11, 1.896791e-11, 1.921616e-11, 1.936892e-11, 1.952493e-11, 
    1.959393e-11, 1.961495e-11, 1.962374e-11,
  1.683516e-11, 1.69854e-11, 1.695616e-11, 1.707766e-11, 1.701022e-11, 
    1.708985e-11, 1.686558e-11, 1.699137e-11, 1.691102e-11, 1.684867e-11, 
    1.731454e-11, 1.70831e-11, 1.755646e-11, 1.740779e-11, 1.778232e-11, 
    1.753328e-11, 1.783273e-11, 1.777514e-11, 1.794877e-11, 1.789895e-11, 
    1.812179e-11, 1.797178e-11, 1.823779e-11, 1.808592e-11, 1.810964e-11, 
    1.796684e-11, 1.712958e-11, 1.728564e-11, 1.712035e-11, 1.714256e-11, 
    1.71326e-11, 1.701161e-11, 1.695076e-11, 1.682371e-11, 1.684675e-11, 
    1.694009e-11, 1.715255e-11, 1.708031e-11, 1.726267e-11, 1.725854e-11, 
    1.746252e-11, 1.737042e-11, 1.771483e-11, 1.761665e-11, 1.790103e-11, 
    1.782932e-11, 1.789766e-11, 1.787693e-11, 1.789793e-11, 1.779281e-11, 
    1.783781e-11, 1.774545e-11, 1.738765e-11, 1.749247e-11, 1.718065e-11, 
    1.699431e-11, 1.687108e-11, 1.678386e-11, 1.679618e-11, 1.681967e-11, 
    1.694063e-11, 1.705472e-11, 1.714189e-11, 1.720031e-11, 1.725795e-11, 
    1.74329e-11, 1.752584e-11, 1.773471e-11, 1.769695e-11, 1.776095e-11, 
    1.78222e-11, 1.792522e-11, 1.790825e-11, 1.795369e-11, 1.775927e-11, 
    1.788838e-11, 1.767545e-11, 1.773358e-11, 1.727357e-11, 1.709979e-11, 
    1.702611e-11, 1.696177e-11, 1.680565e-11, 1.691339e-11, 1.687088e-11, 
    1.697211e-11, 1.703656e-11, 1.700467e-11, 1.72019e-11, 1.712511e-11, 
    1.753136e-11, 1.735586e-11, 1.781505e-11, 1.77047e-11, 1.784154e-11, 
    1.777166e-11, 1.789147e-11, 1.778363e-11, 1.797063e-11, 1.801145e-11, 
    1.798355e-11, 1.809085e-11, 1.777766e-11, 1.789765e-11, 1.700378e-11, 
    1.700897e-11, 1.70332e-11, 1.69268e-11, 1.69203e-11, 1.682307e-11, 
    1.690958e-11, 1.694647e-11, 1.70403e-11, 1.70959e-11, 1.714883e-11, 
    1.726545e-11, 1.739611e-11, 1.757953e-11, 1.771184e-11, 1.780077e-11, 
    1.774622e-11, 1.779437e-11, 1.774055e-11, 1.771534e-11, 1.799614e-11, 
    1.783823e-11, 1.80754e-11, 1.806225e-11, 1.795477e-11, 1.806373e-11, 
    1.701262e-11, 1.698272e-11, 1.687904e-11, 1.696015e-11, 1.68125e-11, 
    1.689507e-11, 1.694263e-11, 1.712669e-11, 1.716727e-11, 1.720491e-11, 
    1.727937e-11, 1.737513e-11, 1.754367e-11, 1.769089e-11, 1.782577e-11, 
    1.781587e-11, 1.781935e-11, 1.784953e-11, 1.777481e-11, 1.786181e-11, 
    1.787643e-11, 1.783822e-11, 1.806048e-11, 1.799686e-11, 1.806197e-11, 
    1.802053e-11, 1.699244e-11, 1.704279e-11, 1.701557e-11, 1.706677e-11, 
    1.703069e-11, 1.719136e-11, 1.723966e-11, 1.746646e-11, 1.737324e-11, 
    1.752172e-11, 1.73883e-11, 1.741191e-11, 1.752655e-11, 1.739551e-11, 
    1.768275e-11, 1.748776e-11, 1.785071e-11, 1.765516e-11, 1.786299e-11, 
    1.782518e-11, 1.78878e-11, 1.794396e-11, 1.801473e-11, 1.814561e-11, 
    1.811527e-11, 1.822496e-11, 1.711798e-11, 1.718351e-11, 1.717775e-11, 
    1.724644e-11, 1.729732e-11, 1.740783e-11, 1.75857e-11, 1.751872e-11, 
    1.764178e-11, 1.766652e-11, 1.747961e-11, 1.759426e-11, 1.722744e-11, 
    1.728647e-11, 1.725132e-11, 1.712314e-11, 1.753413e-11, 1.732267e-11, 
    1.771403e-11, 1.759883e-11, 1.793595e-11, 1.776794e-11, 1.809858e-11, 
    1.824069e-11, 1.837493e-11, 1.853227e-11, 1.721934e-11, 1.717476e-11, 
    1.725462e-11, 1.736537e-11, 1.746843e-11, 1.760584e-11, 1.761994e-11, 
    1.764574e-11, 1.771266e-11, 1.7769e-11, 1.765389e-11, 1.778314e-11, 
    1.730015e-11, 1.755254e-11, 1.715791e-11, 1.727631e-11, 1.735884e-11, 
    1.732263e-11, 1.751108e-11, 1.755562e-11, 1.773712e-11, 1.76432e-11, 
    1.820556e-11, 1.795582e-11, 1.86525e-11, 1.845666e-11, 1.715919e-11, 
    1.721919e-11, 1.74287e-11, 1.732888e-11, 1.761504e-11, 1.768579e-11, 
    1.77434e-11, 1.781714e-11, 1.782512e-11, 1.786888e-11, 1.779719e-11, 
    1.786605e-11, 1.760614e-11, 1.772209e-11, 1.740471e-11, 1.748172e-11, 
    1.744628e-11, 1.740743e-11, 1.752745e-11, 1.765569e-11, 1.765846e-11, 
    1.769966e-11, 1.781597e-11, 1.761621e-11, 1.823786e-11, 1.785282e-11, 
    1.728472e-11, 1.740071e-11, 1.741732e-11, 1.737233e-11, 1.767869e-11, 
    1.756741e-11, 1.786782e-11, 1.778642e-11, 1.791988e-11, 1.785351e-11, 
    1.784375e-11, 1.775868e-11, 1.77058e-11, 1.75725e-11, 1.746438e-11, 
    1.737885e-11, 1.739873e-11, 1.749273e-11, 1.766356e-11, 1.782583e-11, 
    1.779023e-11, 1.790972e-11, 1.759422e-11, 1.772621e-11, 1.767514e-11, 
    1.780845e-11, 1.751694e-11, 1.776499e-11, 1.745378e-11, 1.748097e-11, 
    1.756521e-11, 1.773517e-11, 1.777289e-11, 1.781318e-11, 1.778832e-11, 
    1.766791e-11, 1.764822e-11, 1.756316e-11, 1.75397e-11, 1.747505e-11, 
    1.74216e-11, 1.747043e-11, 1.752177e-11, 1.766796e-11, 1.780015e-11, 
    1.794476e-11, 1.798024e-11, 1.814993e-11, 1.801172e-11, 1.824002e-11, 
    1.80458e-11, 1.838258e-11, 1.777944e-11, 1.804014e-11, 1.756905e-11, 
    1.761955e-11, 1.771102e-11, 1.792163e-11, 1.780782e-11, 1.794097e-11, 
    1.764745e-11, 1.749597e-11, 1.745689e-11, 1.738405e-11, 1.745856e-11, 
    1.745249e-11, 1.752391e-11, 1.750095e-11, 1.767283e-11, 1.758041e-11, 
    1.78435e-11, 1.793992e-11, 1.821345e-11, 1.838199e-11, 1.855427e-11, 
    1.863054e-11, 1.865378e-11, 1.86635e-11,
  1.718953e-11, 1.735434e-11, 1.732224e-11, 1.745561e-11, 1.738157e-11, 
    1.746898e-11, 1.722288e-11, 1.736089e-11, 1.727273e-11, 1.720434e-11, 
    1.771586e-11, 1.746157e-11, 1.798196e-11, 1.781836e-11, 1.823073e-11, 
    1.795645e-11, 1.828629e-11, 1.82228e-11, 1.841423e-11, 1.835929e-11, 
    1.860521e-11, 1.843962e-11, 1.873332e-11, 1.85656e-11, 1.859178e-11, 
    1.843417e-11, 1.751261e-11, 1.76841e-11, 1.750247e-11, 1.752687e-11, 
    1.751592e-11, 1.738309e-11, 1.731634e-11, 1.717697e-11, 1.720223e-11, 
    1.730462e-11, 1.753784e-11, 1.745851e-11, 1.765881e-11, 1.765428e-11, 
    1.787857e-11, 1.777727e-11, 1.815635e-11, 1.804821e-11, 1.836158e-11, 
    1.828252e-11, 1.835787e-11, 1.833501e-11, 1.835816e-11, 1.824228e-11, 
    1.829189e-11, 1.819008e-11, 1.779622e-11, 1.791153e-11, 1.75687e-11, 
    1.736413e-11, 1.722892e-11, 1.713329e-11, 1.714679e-11, 1.717255e-11, 
    1.730522e-11, 1.743041e-11, 1.752612e-11, 1.759029e-11, 1.765363e-11, 
    1.784601e-11, 1.794826e-11, 1.817825e-11, 1.813665e-11, 1.820716e-11, 
    1.827467e-11, 1.838826e-11, 1.836955e-11, 1.841968e-11, 1.820531e-11, 
    1.834764e-11, 1.811297e-11, 1.8177e-11, 1.767084e-11, 1.747989e-11, 
    1.739902e-11, 1.732841e-11, 1.715718e-11, 1.727533e-11, 1.722871e-11, 
    1.733974e-11, 1.741047e-11, 1.737547e-11, 1.759204e-11, 1.750769e-11, 
    1.795433e-11, 1.776127e-11, 1.826679e-11, 1.814519e-11, 1.829599e-11, 
    1.821897e-11, 1.835105e-11, 1.823215e-11, 1.843835e-11, 1.84834e-11, 
    1.845261e-11, 1.857103e-11, 1.822557e-11, 1.835786e-11, 1.737449e-11, 
    1.73802e-11, 1.740679e-11, 1.729003e-11, 1.72829e-11, 1.717628e-11, 
    1.727114e-11, 1.731161e-11, 1.741458e-11, 1.747562e-11, 1.753375e-11, 
    1.766188e-11, 1.780553e-11, 1.800736e-11, 1.815306e-11, 1.825104e-11, 
    1.819093e-11, 1.824399e-11, 1.818468e-11, 1.815691e-11, 1.846651e-11, 
    1.829235e-11, 1.855398e-11, 1.853945e-11, 1.842087e-11, 1.854109e-11, 
    1.73842e-11, 1.735138e-11, 1.723765e-11, 1.732662e-11, 1.716468e-11, 
    1.725523e-11, 1.730741e-11, 1.750944e-11, 1.7554e-11, 1.759535e-11, 
    1.767717e-11, 1.778245e-11, 1.796787e-11, 1.812998e-11, 1.82786e-11, 
    1.826769e-11, 1.827153e-11, 1.83048e-11, 1.822244e-11, 1.831834e-11, 
    1.833446e-11, 1.829233e-11, 1.853751e-11, 1.84673e-11, 1.853915e-11, 
    1.849342e-11, 1.736205e-11, 1.741731e-11, 1.738744e-11, 1.744364e-11, 
    1.740403e-11, 1.758047e-11, 1.763354e-11, 1.788292e-11, 1.778037e-11, 
    1.794372e-11, 1.779693e-11, 1.78229e-11, 1.794906e-11, 1.780485e-11, 
    1.812102e-11, 1.790636e-11, 1.830609e-11, 1.809065e-11, 1.831964e-11, 
    1.827796e-11, 1.8347e-11, 1.840894e-11, 1.848702e-11, 1.86315e-11, 
    1.8598e-11, 1.871915e-11, 1.749987e-11, 1.757185e-11, 1.756551e-11, 
    1.764098e-11, 1.76969e-11, 1.781841e-11, 1.801414e-11, 1.794041e-11, 
    1.807588e-11, 1.810314e-11, 1.789737e-11, 1.802357e-11, 1.762011e-11, 
    1.768498e-11, 1.764634e-11, 1.750554e-11, 1.795738e-11, 1.772479e-11, 
    1.815547e-11, 1.802859e-11, 1.84001e-11, 1.821487e-11, 1.857956e-11, 
    1.873654e-11, 1.888489e-11, 1.905896e-11, 1.76112e-11, 1.756222e-11, 
    1.764997e-11, 1.777173e-11, 1.788508e-11, 1.803632e-11, 1.805183e-11, 
    1.808024e-11, 1.815395e-11, 1.821603e-11, 1.808923e-11, 1.823161e-11, 
    1.770004e-11, 1.797764e-11, 1.754372e-11, 1.767383e-11, 1.776454e-11, 
    1.772472e-11, 1.7932e-11, 1.798102e-11, 1.818091e-11, 1.807745e-11, 
    1.869773e-11, 1.842203e-11, 1.919204e-11, 1.897529e-11, 1.754512e-11, 
    1.761103e-11, 1.784137e-11, 1.773159e-11, 1.804644e-11, 1.812435e-11, 
    1.818782e-11, 1.82691e-11, 1.827789e-11, 1.832614e-11, 1.82471e-11, 
    1.832301e-11, 1.803664e-11, 1.816434e-11, 1.781497e-11, 1.78997e-11, 
    1.78607e-11, 1.781796e-11, 1.795001e-11, 1.809122e-11, 1.809425e-11, 
    1.813964e-11, 1.826785e-11, 1.804772e-11, 1.873345e-11, 1.830847e-11, 
    1.768304e-11, 1.781059e-11, 1.782885e-11, 1.777936e-11, 1.811653e-11, 
    1.7994e-11, 1.832496e-11, 1.823523e-11, 1.838237e-11, 1.830918e-11, 
    1.829842e-11, 1.820466e-11, 1.814639e-11, 1.799961e-11, 1.788062e-11, 
    1.778654e-11, 1.780839e-11, 1.791181e-11, 1.809988e-11, 1.827868e-11, 
    1.823944e-11, 1.837117e-11, 1.802352e-11, 1.81689e-11, 1.811264e-11, 
    1.825951e-11, 1.793846e-11, 1.821165e-11, 1.786895e-11, 1.789887e-11, 
    1.799158e-11, 1.817877e-11, 1.822032e-11, 1.826473e-11, 1.823732e-11, 
    1.810466e-11, 1.808298e-11, 1.798932e-11, 1.79635e-11, 1.789235e-11, 
    1.783355e-11, 1.788727e-11, 1.794377e-11, 1.810472e-11, 1.825037e-11, 
    1.840982e-11, 1.844895e-11, 1.863629e-11, 1.848371e-11, 1.873583e-11, 
    1.852136e-11, 1.889339e-11, 1.822756e-11, 1.851508e-11, 1.79958e-11, 
    1.80514e-11, 1.815216e-11, 1.838433e-11, 1.825882e-11, 1.840565e-11, 
    1.808213e-11, 1.791538e-11, 1.787237e-11, 1.779225e-11, 1.787421e-11, 
    1.786753e-11, 1.794612e-11, 1.792085e-11, 1.811008e-11, 1.800831e-11, 
    1.829815e-11, 1.840449e-11, 1.870643e-11, 1.889272e-11, 1.908329e-11, 
    1.916771e-11, 1.919345e-11, 1.920421e-11,
  1.871146e-11, 1.888764e-11, 1.885332e-11, 1.899597e-11, 1.891676e-11, 
    1.901028e-11, 1.87471e-11, 1.889466e-11, 1.880038e-11, 1.872728e-11, 
    1.927461e-11, 1.900235e-11, 1.955982e-11, 1.938441e-11, 1.982681e-11, 
    1.953247e-11, 1.988647e-11, 1.981828e-11, 2.002394e-11, 1.996489e-11, 
    2.022933e-11, 2.005123e-11, 2.036721e-11, 2.018671e-11, 2.021488e-11, 
    2.004537e-11, 1.905696e-11, 1.92406e-11, 1.904611e-11, 1.907222e-11, 
    1.90605e-11, 1.89184e-11, 1.884702e-11, 1.869803e-11, 1.872503e-11, 
    1.883448e-11, 1.908397e-11, 1.899906e-11, 1.921347e-11, 1.920862e-11, 
    1.944895e-11, 1.934037e-11, 1.974693e-11, 1.963088e-11, 1.996735e-11, 
    1.988242e-11, 1.996336e-11, 1.99388e-11, 1.996368e-11, 1.98392e-11, 
    1.989248e-11, 1.978314e-11, 1.936068e-11, 1.948428e-11, 1.9117e-11, 
    1.889813e-11, 1.875356e-11, 1.865137e-11, 1.866579e-11, 1.869332e-11, 
    1.883512e-11, 1.896901e-11, 1.907142e-11, 1.91401e-11, 1.920792e-11, 
    1.941406e-11, 1.952368e-11, 1.977045e-11, 1.972578e-11, 1.980149e-11, 
    1.987398e-11, 1.999603e-11, 1.997591e-11, 2.002979e-11, 1.979949e-11, 
    1.995238e-11, 1.970036e-11, 1.97691e-11, 1.92264e-11, 1.902195e-11, 
    1.893545e-11, 1.885991e-11, 1.867689e-11, 1.880317e-11, 1.875333e-11, 
    1.887203e-11, 1.894768e-11, 1.891024e-11, 1.914198e-11, 1.905169e-11, 
    1.953019e-11, 1.932323e-11, 1.986552e-11, 1.973495e-11, 1.989689e-11, 
    1.981416e-11, 1.995604e-11, 1.982832e-11, 2.004987e-11, 2.009831e-11, 
    2.00652e-11, 2.019255e-11, 1.982125e-11, 1.996336e-11, 1.890919e-11, 
    1.891529e-11, 1.894374e-11, 1.881889e-11, 1.881126e-11, 1.86973e-11, 
    1.879868e-11, 1.884196e-11, 1.895207e-11, 1.901738e-11, 1.907958e-11, 
    1.921676e-11, 1.937066e-11, 1.958705e-11, 1.974339e-11, 1.98486e-11, 
    1.978405e-11, 1.984103e-11, 1.977734e-11, 1.974753e-11, 2.008015e-11, 
    1.989298e-11, 2.01742e-11, 2.015858e-11, 2.003108e-11, 2.016034e-11, 
    1.891958e-11, 1.888447e-11, 1.876288e-11, 1.8858e-11, 1.868491e-11, 
    1.878168e-11, 1.883746e-11, 1.905358e-11, 1.910125e-11, 1.914552e-11, 
    1.923314e-11, 1.934592e-11, 1.95447e-11, 1.971863e-11, 1.98782e-11, 
    1.986648e-11, 1.987061e-11, 1.990635e-11, 1.981789e-11, 1.99209e-11, 
    1.993822e-11, 1.989295e-11, 2.015649e-11, 2.008099e-11, 2.015825e-11, 
    2.010907e-11, 1.889588e-11, 1.8955e-11, 1.892304e-11, 1.898316e-11, 
    1.89408e-11, 1.91296e-11, 1.918643e-11, 1.945362e-11, 1.93437e-11, 
    1.951881e-11, 1.936144e-11, 1.938927e-11, 1.952454e-11, 1.936992e-11, 
    1.970902e-11, 1.947876e-11, 1.990774e-11, 1.967644e-11, 1.992229e-11, 
    1.987751e-11, 1.995168e-11, 2.001825e-11, 2.010219e-11, 2.025761e-11, 
    2.022156e-11, 2.035194e-11, 1.904332e-11, 1.912037e-11, 1.911358e-11, 
    1.919438e-11, 1.925427e-11, 1.938445e-11, 1.959432e-11, 1.951525e-11, 
    1.966056e-11, 1.968981e-11, 1.94691e-11, 1.960444e-11, 1.917204e-11, 
    1.924152e-11, 1.920013e-11, 1.90494e-11, 1.953346e-11, 1.928415e-11, 
    1.974598e-11, 1.960983e-11, 2.000875e-11, 1.980978e-11, 2.020173e-11, 
    2.037068e-11, 2.053044e-11, 2.07181e-11, 1.916249e-11, 1.911006e-11, 
    1.920401e-11, 1.933444e-11, 1.945592e-11, 1.961812e-11, 1.963476e-11, 
    1.966525e-11, 1.974435e-11, 1.981101e-11, 1.96749e-11, 1.982773e-11, 
    1.925766e-11, 1.955518e-11, 1.909026e-11, 1.922957e-11, 1.932674e-11, 
    1.928407e-11, 1.950622e-11, 1.95588e-11, 1.977331e-11, 1.966225e-11, 
    2.032891e-11, 2.003234e-11, 2.086166e-11, 2.062789e-11, 1.909175e-11, 
    1.916231e-11, 1.940907e-11, 1.929143e-11, 1.962897e-11, 1.971259e-11, 
    1.978071e-11, 1.9868e-11, 1.987744e-11, 1.992928e-11, 1.984437e-11, 
    1.992592e-11, 1.961846e-11, 1.975551e-11, 1.938077e-11, 1.947159e-11, 
    1.942978e-11, 1.938398e-11, 1.952554e-11, 1.967703e-11, 1.968027e-11, 
    1.9729e-11, 1.986671e-11, 1.963035e-11, 2.036738e-11, 1.991033e-11, 
    1.923943e-11, 1.937609e-11, 1.939565e-11, 1.934261e-11, 1.970419e-11, 
    1.957273e-11, 1.992801e-11, 1.983162e-11, 1.99897e-11, 1.991105e-11, 
    1.98995e-11, 1.979879e-11, 1.973624e-11, 1.957874e-11, 1.945114e-11, 
    1.93503e-11, 1.937372e-11, 1.948458e-11, 1.968632e-11, 1.987829e-11, 
    1.983615e-11, 1.997766e-11, 1.960438e-11, 1.97604e-11, 1.970002e-11, 
    1.98577e-11, 1.951315e-11, 1.980634e-11, 1.943862e-11, 1.94707e-11, 
    1.957012e-11, 1.977101e-11, 1.981562e-11, 1.986331e-11, 1.983387e-11, 
    1.969146e-11, 1.966818e-11, 1.95677e-11, 1.954001e-11, 1.946371e-11, 
    1.940068e-11, 1.945827e-11, 1.951886e-11, 1.969152e-11, 1.984789e-11, 
    2.00192e-11, 2.006126e-11, 2.026279e-11, 2.009866e-11, 2.036995e-11, 
    2.013918e-11, 2.053964e-11, 1.982341e-11, 2.013239e-11, 1.957465e-11, 
    1.963429e-11, 1.974245e-11, 1.999181e-11, 1.985696e-11, 2.001472e-11, 
    1.966727e-11, 1.948842e-11, 1.944229e-11, 1.935642e-11, 1.944426e-11, 
    1.943711e-11, 1.952136e-11, 1.949426e-11, 1.969726e-11, 1.958807e-11, 
    1.989921e-11, 2.001348e-11, 2.033825e-11, 2.053889e-11, 2.074432e-11, 
    2.083541e-11, 2.086318e-11, 2.087479e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
