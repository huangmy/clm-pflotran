netcdf ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-01-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "timestep fractional area burned for crop" ;
		BAF_CROP:units = "proportion" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "timestep fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned in this timestep" ;
		LFC2:units = "per timestep" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "timestep fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/timestep" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 08/14/14 18:42:38" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "bandre" ;
		:version = "clm4_5_67" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c130821.nc" ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-01-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 10102 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "08/14/14" ;

 time_written =
  "18:42:38" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  4.490659e-14, 4.502776e-14, 4.500422e-14, 4.510186e-14, 4.504772e-14, 
    4.511163e-14, 4.493118e-14, 4.503255e-14, 4.496786e-14, 4.491752e-14, 
    4.529107e-14, 4.510622e-14, 4.548291e-14, 4.536523e-14, 4.566065e-14, 
    4.546458e-14, 4.570015e-14, 4.565504e-14, 4.579087e-14, 4.575198e-14, 
    4.592545e-14, 4.580882e-14, 4.601533e-14, 4.589763e-14, 4.591603e-14, 
    4.580496e-14, 4.514348e-14, 4.526806e-14, 4.513609e-14, 4.515386e-14, 
    4.51459e-14, 4.504883e-14, 4.499986e-14, 4.489735e-14, 4.491597e-14, 
    4.499127e-14, 4.516186e-14, 4.510401e-14, 4.524983e-14, 4.524654e-14, 
    4.540864e-14, 4.533558e-14, 4.560769e-14, 4.553044e-14, 4.57536e-14, 
    4.569751e-14, 4.575096e-14, 4.573476e-14, 4.575117e-14, 4.56689e-14, 
    4.570415e-14, 4.563174e-14, 4.534926e-14, 4.543234e-14, 4.518434e-14, 
    4.503489e-14, 4.493562e-14, 4.48651e-14, 4.487507e-14, 4.489407e-14, 
    4.499171e-14, 4.508348e-14, 4.515334e-14, 4.520005e-14, 4.524606e-14, 
    4.538511e-14, 4.545872e-14, 4.562329e-14, 4.559364e-14, 4.564389e-14, 
    4.569193e-14, 4.577248e-14, 4.575923e-14, 4.57947e-14, 4.564259e-14, 
    4.57437e-14, 4.557676e-14, 4.562242e-14, 4.525843e-14, 4.511962e-14, 
    4.506046e-14, 4.500874e-14, 4.488274e-14, 4.496976e-14, 4.493546e-14, 
    4.501708e-14, 4.506889e-14, 4.504327e-14, 4.520133e-14, 4.51399e-14, 
    4.546308e-14, 4.532399e-14, 4.568633e-14, 4.559973e-14, 4.570708e-14, 
    4.565232e-14, 4.574612e-14, 4.56617e-14, 4.580791e-14, 4.583971e-14, 
    4.581798e-14, 4.590147e-14, 4.565702e-14, 4.575095e-14, 4.504255e-14, 
    4.504672e-14, 4.50662e-14, 4.498056e-14, 4.497533e-14, 4.489683e-14, 
    4.496669e-14, 4.499642e-14, 4.50719e-14, 4.51165e-14, 4.515889e-14, 
    4.525204e-14, 4.535595e-14, 4.550115e-14, 4.560534e-14, 4.567514e-14, 
    4.563236e-14, 4.567013e-14, 4.56279e-14, 4.56081e-14, 4.582779e-14, 
    4.570447e-14, 4.588947e-14, 4.587924e-14, 4.579554e-14, 4.58804e-14, 
    4.504966e-14, 4.502562e-14, 4.494205e-14, 4.500745e-14, 4.488828e-14, 
    4.495499e-14, 4.499331e-14, 4.514116e-14, 4.517365e-14, 4.520372e-14, 
    4.526313e-14, 4.533932e-14, 4.547282e-14, 4.558886e-14, 4.569473e-14, 
    4.568698e-14, 4.56897e-14, 4.571333e-14, 4.565478e-14, 4.572294e-14, 
    4.573436e-14, 4.570447e-14, 4.587787e-14, 4.582837e-14, 4.587902e-14, 
    4.58468e-14, 4.503343e-14, 4.50739e-14, 4.505203e-14, 4.509313e-14, 
    4.506417e-14, 4.519288e-14, 4.523144e-14, 4.541174e-14, 4.533781e-14, 
    4.545548e-14, 4.534978e-14, 4.536851e-14, 4.545926e-14, 4.53555e-14, 
    4.558244e-14, 4.542859e-14, 4.571425e-14, 4.556073e-14, 4.572385e-14, 
    4.569427e-14, 4.574327e-14, 4.578711e-14, 4.584228e-14, 4.594395e-14, 
    4.592042e-14, 4.600542e-14, 4.51342e-14, 4.518662e-14, 4.518203e-14, 
    4.523688e-14, 4.527743e-14, 4.536528e-14, 4.550603e-14, 4.545313e-14, 
    4.555025e-14, 4.556973e-14, 4.542219e-14, 4.551277e-14, 4.522171e-14, 
    4.526876e-14, 4.524076e-14, 4.513832e-14, 4.546528e-14, 4.529759e-14, 
    4.560706e-14, 4.551639e-14, 4.578086e-14, 4.564937e-14, 4.590746e-14, 
    4.601754e-14, 4.612116e-14, 4.624198e-14, 4.521525e-14, 4.517964e-14, 
    4.524341e-14, 4.533154e-14, 4.541332e-14, 4.552192e-14, 4.553304e-14, 
    4.555336e-14, 4.560599e-14, 4.565023e-14, 4.555976e-14, 4.566132e-14, 
    4.527962e-14, 4.547984e-14, 4.516615e-14, 4.526067e-14, 4.532636e-14, 
    4.529757e-14, 4.544709e-14, 4.548229e-14, 4.562519e-14, 4.555137e-14, 
    4.599036e-14, 4.579634e-14, 4.633398e-14, 4.618398e-14, 4.516718e-14, 
    4.521514e-14, 4.538182e-14, 4.530255e-14, 4.552917e-14, 4.558485e-14, 
    4.563014e-14, 4.568796e-14, 4.569422e-14, 4.572846e-14, 4.567234e-14, 
    4.572626e-14, 4.552215e-14, 4.56134e-14, 4.536281e-14, 4.542384e-14, 
    4.539578e-14, 4.536497e-14, 4.546003e-14, 4.556118e-14, 4.556338e-14, 
    4.559576e-14, 4.568695e-14, 4.553009e-14, 4.60153e-14, 4.571581e-14, 
    4.52674e-14, 4.53596e-14, 4.537281e-14, 4.53371e-14, 4.557929e-14, 
    4.549159e-14, 4.572763e-14, 4.566389e-14, 4.576832e-14, 4.571644e-14, 
    4.57088e-14, 4.564213e-14, 4.560059e-14, 4.549561e-14, 4.541011e-14, 
    4.534228e-14, 4.535806e-14, 4.543255e-14, 4.556737e-14, 4.569476e-14, 
    4.566686e-14, 4.576039e-14, 4.551275e-14, 4.561662e-14, 4.557649e-14, 
    4.568115e-14, 4.545171e-14, 4.5647e-14, 4.540172e-14, 4.542326e-14, 
    4.548985e-14, 4.562364e-14, 4.565328e-14, 4.568485e-14, 4.566539e-14, 
    4.55708e-14, 4.555531e-14, 4.548824e-14, 4.54697e-14, 4.541857e-14, 
    4.537621e-14, 4.54149e-14, 4.545552e-14, 4.557085e-14, 4.567464e-14, 
    4.578773e-14, 4.581541e-14, 4.594725e-14, 4.583988e-14, 4.601695e-14, 
    4.586634e-14, 4.612697e-14, 4.565836e-14, 4.586199e-14, 4.549289e-14, 
    4.553273e-14, 4.560467e-14, 4.576966e-14, 4.568066e-14, 4.578475e-14, 
    4.555471e-14, 4.54351e-14, 4.540418e-14, 4.53464e-14, 4.540551e-14, 
    4.54007e-14, 4.545723e-14, 4.543907e-14, 4.557468e-14, 4.550186e-14, 
    4.570859e-14, 4.578394e-14, 4.59965e-14, 4.612657e-14, 4.625888e-14, 
    4.631722e-14, 4.633497e-14, 4.634239e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -1.89636e-14, -1.898576e-14, -1.898144e-14, -1.899932e-14, -1.898938e-14, 
    -1.90011e-14, -1.896806e-14, -1.898667e-14, -1.897478e-14, -1.896555e-14, 
    -1.903401e-14, -1.900011e-14, -1.906878e-14, -1.904732e-14, 
    -1.910104e-14, -1.906548e-14, -1.910818e-14, -1.909995e-14, 
    -1.912453e-14, -1.911749e-14, -1.914899e-14, -1.912777e-14, 
    -1.916516e-14, -1.914389e-14, -1.914725e-14, -1.912708e-14, 
    -1.900688e-14, -1.902982e-14, -1.900553e-14, -1.900881e-14, 
    -1.900732e-14, -1.898961e-14, -1.898072e-14, -1.896185e-14, 
    -1.896527e-14, -1.89791e-14, -1.901027e-14, -1.899966e-14, -1.902626e-14, 
    -1.902566e-14, -1.905521e-14, -1.90419e-14, -1.909136e-14, -1.907731e-14, 
    -1.911778e-14, -1.910763e-14, -1.911732e-14, -1.911437e-14, 
    -1.911735e-14, -1.910246e-14, -1.910885e-14, -1.909571e-14, -1.90444e-14, 
    -1.905954e-14, -1.901435e-14, -1.898717e-14, -1.896889e-14, 
    -1.895595e-14, -1.895778e-14, -1.896129e-14, -1.897918e-14, 
    -1.899591e-14, -1.900866e-14, -1.901719e-14, -1.902557e-14, 
    -1.905107e-14, -1.906438e-14, -1.909423e-14, -1.90888e-14, -1.909796e-14, 
    -1.910662e-14, -1.912122e-14, -1.911881e-14, -1.912525e-14, 
    -1.909767e-14, -1.911603e-14, -1.908571e-14, -1.909402e-14, 
    -1.902808e-14, -1.900251e-14, -1.899182e-14, -1.898228e-14, -1.89592e-14, 
    -1.897516e-14, -1.896887e-14, -1.898377e-14, -1.899325e-14, 
    -1.898855e-14, -1.901742e-14, -1.900621e-14, -1.906517e-14, 
    -1.903983e-14, -1.910561e-14, -1.908991e-14, -1.910936e-14, 
    -1.909943e-14, -1.911646e-14, -1.910113e-14, -1.912763e-14, 
    -1.913341e-14, -1.912946e-14, -1.914454e-14, -1.910029e-14, 
    -1.911734e-14, -1.898843e-14, -1.89892e-14, -1.899275e-14, -1.897714e-14, 
    -1.897617e-14, -1.896177e-14, -1.897456e-14, -1.898002e-14, 
    -1.899378e-14, -1.900195e-14, -1.900969e-14, -1.902669e-14, 
    -1.904566e-14, -1.907205e-14, -1.909093e-14, -1.910357e-14, -1.90958e-14, 
    -1.910266e-14, -1.9095e-14, -1.90914e-14, -1.913126e-14, -1.910892e-14, 
    -1.914237e-14, -1.914052e-14, -1.912541e-14, -1.914072e-14, 
    -1.898973e-14, -1.898532e-14, -1.897006e-14, -1.8982e-14, -1.89602e-14, 
    -1.897244e-14, -1.897949e-14, -1.90065e-14, -1.901237e-14, -1.901788e-14, 
    -1.902869e-14, -1.904258e-14, -1.90669e-14, -1.908796e-14, -1.910711e-14, 
    -1.910571e-14, -1.910621e-14, -1.91105e-14, -1.909989e-14, -1.911224e-14, 
    -1.911433e-14, -1.910889e-14, -1.914027e-14, -1.913131e-14, 
    -1.914048e-14, -1.913464e-14, -1.898675e-14, -1.899416e-14, 
    -1.899016e-14, -1.899769e-14, -1.89924e-14, -1.901595e-14, -1.9023e-14, 
    -1.905583e-14, -1.904232e-14, -1.906376e-14, -1.904448e-14, 
    -1.904791e-14, -1.906455e-14, -1.904551e-14, -1.908685e-14, 
    -1.905893e-14, -1.911067e-14, -1.908296e-14, -1.911241e-14, 
    -1.910703e-14, -1.911591e-14, -1.912387e-14, -1.913383e-14, 
    -1.915226e-14, -1.914799e-14, -1.916333e-14, -1.900517e-14, 
    -1.901478e-14, -1.901389e-14, -1.902391e-14, -1.903132e-14, 
    -1.904729e-14, -1.907291e-14, -1.906327e-14, -1.90809e-14, -1.908446e-14, 
    -1.905763e-14, -1.907415e-14, -1.902117e-14, -1.90298e-14, -1.902463e-14, 
    -1.900595e-14, -1.906555e-14, -1.903505e-14, -1.909125e-14, 
    -1.907478e-14, -1.912274e-14, -1.909897e-14, -1.914564e-14, 
    -1.916563e-14, -1.918419e-14, -1.920605e-14, -1.901997e-14, 
    -1.901345e-14, -1.902509e-14, -1.904123e-14, -1.905605e-14, 
    -1.907579e-14, -1.907778e-14, -1.908149e-14, -1.909102e-14, 
    -1.909905e-14, -1.90827e-14, -1.910106e-14, -1.903189e-14, -1.906817e-14, 
    -1.901103e-14, -1.902834e-14, -1.904026e-14, -1.903499e-14, 
    -1.906216e-14, -1.906856e-14, -1.909456e-14, -1.908111e-14, 
    -1.916074e-14, -1.912561e-14, -1.922252e-14, -1.919559e-14, 
    -1.901119e-14, -1.901993e-14, -1.905035e-14, -1.903589e-14, 
    -1.907708e-14, -1.908721e-14, -1.90954e-14, -1.910593e-14, -1.910703e-14, 
    -1.911325e-14, -1.910306e-14, -1.911283e-14, -1.907583e-14, 
    -1.909238e-14, -1.904683e-14, -1.905797e-14, -1.905283e-14, 
    -1.904722e-14, -1.906452e-14, -1.908297e-14, -1.908329e-14, 
    -1.908922e-14, -1.9106e-14, -1.907725e-14, -1.916539e-14, -1.911119e-14, 
    -1.902946e-14, -1.904635e-14, -1.904868e-14, -1.904215e-14, -1.90862e-14, 
    -1.907028e-14, -1.911309e-14, -1.910153e-14, -1.912045e-14, 
    -1.911106e-14, -1.910968e-14, -1.909758e-14, -1.909006e-14, 
    -1.907102e-14, -1.905547e-14, -1.904309e-14, -1.904597e-14, 
    -1.905956e-14, -1.908408e-14, -1.910716e-14, -1.910212e-14, 
    -1.911901e-14, -1.90741e-14, -1.9093e-14, -1.908572e-14, -1.910467e-14, 
    -1.906303e-14, -1.909871e-14, -1.905391e-14, -1.905783e-14, 
    -1.906996e-14, -1.909433e-14, -1.909961e-14, -1.910536e-14, -1.91018e-14, 
    -1.908469e-14, -1.908185e-14, -1.906965e-14, -1.906631e-14, 
    -1.905697e-14, -1.904927e-14, -1.905633e-14, -1.906375e-14, 
    -1.908467e-14, -1.910352e-14, -1.912399e-14, -1.912897e-14, 
    -1.915298e-14, -1.913353e-14, -1.91657e-14, -1.91385e-14, -1.918545e-14, 
    -1.910067e-14, -1.913756e-14, -1.907049e-14, -1.907772e-14, 
    -1.909087e-14, -1.912079e-14, -1.910458e-14, -1.912351e-14, 
    -1.908173e-14, -1.906007e-14, -1.905436e-14, -1.904386e-14, -1.90546e-14, 
    -1.905373e-14, -1.9064e-14, -1.90607e-14, -1.908536e-14, -1.907212e-14, 
    -1.910966e-14, -1.912334e-14, -1.916175e-14, -1.918525e-14, 
    -1.920898e-14, -1.921948e-14, -1.922266e-14, -1.9224e-14 ;

 CH4_SURF_DIFF_UNSAT =
  1.517012e-11, 1.516283e-11, 1.516434e-11, 1.515781e-11, 1.516153e-11, 
    1.515711e-11, 1.516874e-11, 1.516251e-11, 1.516658e-11, 1.516952e-11, 
    1.514272e-11, 1.51575e-11, 1.504166e-11, 1.504085e-11, 1.503779e-11, 
    1.504169e-11, 1.503605e-11, 1.503803e-11, 1.503076e-11, 1.503326e-11, 
    1.501937e-11, 1.502949e-11, 1.500936e-11, 1.502209e-11, 1.502031e-11, 
    1.502977e-11, 1.515479e-11, 1.514473e-11, 1.515534e-11, 1.515401e-11, 
    1.515461e-11, 1.516145e-11, 1.516459e-11, 1.517064e-11, 1.516961e-11, 
    1.516514e-11, 1.51534e-11, 1.515767e-11, 1.514636e-11, 1.514664e-11, 
    1.504145e-11, 1.504025e-11, 1.503963e-11, 1.504127e-11, 1.503316e-11, 
    1.503619e-11, 1.503331e-11, 1.503426e-11, 1.50333e-11, 1.503747e-11, 
    1.503586e-11, 1.503888e-11, 1.504054e-11, 1.504163e-11, 1.515167e-11, 
    1.516234e-11, 1.516848e-11, 1.517238e-11, 1.517185e-11, 1.517081e-11, 
    1.516511e-11, 1.515911e-11, 1.515406e-11, 1.515044e-11, 1.514668e-11, 
    1.504113e-11, 1.50417e-11, 1.503915e-11, 1.504003e-11, 1.503844e-11, 
    1.503646e-11, 1.503198e-11, 1.503282e-11, 1.503048e-11, 1.50385e-11, 
    1.503373e-11, 1.504044e-11, 1.503919e-11, 1.514555e-11, 1.515655e-11, 
    1.516065e-11, 1.516405e-11, 1.517143e-11, 1.516646e-11, 1.516848e-11, 
    1.516353e-11, 1.516011e-11, 1.516183e-11, 1.515034e-11, 1.515506e-11, 
    1.50417e-11, 1.503996e-11, 1.503671e-11, 1.503986e-11, 1.503572e-11, 
    1.503814e-11, 1.50336e-11, 1.503777e-11, 1.502955e-11, 1.502711e-11, 
    1.50288e-11, 1.502174e-11, 1.503796e-11, 1.503331e-11, 1.516188e-11, 
    1.51616e-11, 1.51603e-11, 1.51658e-11, 1.516612e-11, 1.517067e-11, 
    1.516665e-11, 1.516483e-11, 1.515991e-11, 1.515678e-11, 1.515364e-11, 
    1.514617e-11, 1.504067e-11, 1.504156e-11, 1.50397e-11, 1.503721e-11, 
    1.503887e-11, 1.503743e-11, 1.503901e-11, 1.503963e-11, 1.502805e-11, 
    1.503584e-11, 1.502285e-11, 1.502378e-11, 1.503042e-11, 1.502368e-11, 
    1.516141e-11, 1.516299e-11, 1.516811e-11, 1.516415e-11, 1.517114e-11, 
    1.516734e-11, 1.516501e-11, 1.515495e-11, 1.515251e-11, 1.515014e-11, 
    1.514522e-11, 1.504033e-11, 1.50417e-11, 1.504014e-11, 1.503633e-11, 
    1.503669e-11, 1.503656e-11, 1.503541e-11, 1.503805e-11, 1.50349e-11, 
    1.503427e-11, 1.503585e-11, 1.50239e-11, 1.502802e-11, 1.50238e-11, 
    1.502656e-11, 1.516248e-11, 1.515977e-11, 1.516125e-11, 1.515843e-11, 
    1.516043e-11, 1.515099e-11, 1.514786e-11, 1.504147e-11, 1.50403e-11, 
    1.504171e-11, 1.504056e-11, 1.504091e-11, 1.504168e-11, 1.504068e-11, 
    1.504028e-11, 1.504159e-11, 1.503536e-11, 1.504074e-11, 1.503485e-11, 
    1.503635e-11, 1.503377e-11, 1.503101e-11, 1.502692e-11, 1.501749e-11, 
    1.50199e-11, 1.501058e-11, 1.515549e-11, 1.515149e-11, 1.515186e-11, 
    1.514744e-11, 1.514398e-11, 1.504086e-11, 1.504153e-11, 1.504172e-11, 
    1.504097e-11, 1.504059e-11, 1.504158e-11, 1.504146e-11, 1.514868e-11, 
    1.514471e-11, 1.514711e-11, 1.515517e-11, 1.50417e-11, 1.514218e-11, 
    1.503965e-11, 1.504143e-11, 1.503143e-11, 1.503823e-11, 1.502116e-11, 
    1.500907e-11, 1.499495e-11, 1.497481e-11, 1.514922e-11, 1.515205e-11, 
    1.51469e-11, 1.504014e-11, 1.50415e-11, 1.504137e-11, 1.504123e-11, 
    1.504091e-11, 1.503969e-11, 1.503822e-11, 1.504078e-11, 1.503779e-11, 
    1.514374e-11, 1.504168e-11, 1.515308e-11, 1.51454e-11, 1.504002e-11, 
    1.51422e-11, 1.504171e-11, 1.504168e-11, 1.503909e-11, 1.504095e-11, 
    1.501232e-11, 1.503035e-11, 1.495682e-11, 1.498497e-11, 1.515301e-11, 
    1.514923e-11, 1.504111e-11, 1.514176e-11, 1.504129e-11, 1.504024e-11, 
    1.503894e-11, 1.503663e-11, 1.503635e-11, 1.50346e-11, 1.503733e-11, 
    1.503473e-11, 1.504137e-11, 1.503947e-11, 1.504082e-11, 1.504158e-11, 
    1.504132e-11, 1.504086e-11, 1.504173e-11, 1.504075e-11, 1.504072e-11, 
    1.503996e-11, 1.503661e-11, 1.504128e-11, 1.50093e-11, 1.503521e-11, 
    1.514486e-11, 1.504073e-11, 1.504098e-11, 1.504029e-11, 1.504038e-11, 
    1.504163e-11, 1.503465e-11, 1.503769e-11, 1.503225e-11, 1.503525e-11, 
    1.503564e-11, 1.503852e-11, 1.503984e-11, 1.504161e-11, 1.504147e-11, 
    1.504041e-11, 1.504073e-11, 1.504163e-11, 1.504062e-11, 1.503632e-11, 
    1.503755e-11, 1.503275e-11, 1.504147e-11, 1.503936e-11, 1.504043e-11, 
    1.503695e-11, 1.504171e-11, 1.503828e-11, 1.504139e-11, 1.504159e-11, 
    1.504164e-11, 1.503913e-11, 1.50381e-11, 1.503677e-11, 1.503763e-11, 
    1.504056e-11, 1.504087e-11, 1.504166e-11, 1.504171e-11, 1.504155e-11, 
    1.504104e-11, 1.504152e-11, 1.504171e-11, 1.504056e-11, 1.503722e-11, 
    1.503096e-11, 1.5029e-11, 1.50171e-11, 1.502707e-11, 1.500909e-11, 
    1.502482e-11, 1.499401e-11, 1.503787e-11, 1.502524e-11, 1.504163e-11, 
    1.504124e-11, 1.503971e-11, 1.503213e-11, 1.503697e-11, 1.503115e-11, 
    1.504088e-11, 1.504164e-11, 1.504142e-11, 1.504049e-11, 1.504143e-11, 
    1.504138e-11, 1.504172e-11, 1.504168e-11, 1.504048e-11, 1.504157e-11, 
    1.503564e-11, 1.503121e-11, 1.501163e-11, 1.499411e-11, 1.497172e-11, 
    1.496029e-11, 1.495663e-11, 1.495507e-11 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931945e-23, 1.931947e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.93194e-23, 1.931941e-23, 1.931939e-23, 1.93194e-23, 1.93194e-23, 
    1.931941e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931945e-23, 1.931944e-23, 1.931946e-23, 
    1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931945e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.931941e-23, 1.93194e-23, 1.931942e-23, 1.931941e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.93194e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931941e-23, 1.931942e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931941e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931944e-23, 1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.93194e-23, 
    1.93194e-23, 1.931939e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931943e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.93194e-23, 
    1.931939e-23, 1.931938e-23, 1.931937e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931945e-23, 1.931944e-23, 1.931946e-23, 1.931945e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 
    1.931939e-23, 1.931941e-23, 1.931936e-23, 1.931938e-23, 1.931946e-23, 
    1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931939e-23, 1.931942e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 
    1.931944e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 
    1.931942e-23, 1.931944e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931941e-23, 1.931941e-23, 1.93194e-23, 1.931941e-23, 1.931939e-23, 
    1.93194e-23, 1.931938e-23, 1.931942e-23, 1.93194e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 
    1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931941e-23, 1.931939e-23, 1.931938e-23, 1.931937e-23, 
    1.931937e-23, 1.931936e-23, 1.931936e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.975377e-24, 1.975379e-24, 1.975374e-24, 1.975376e-24, 1.975372e-24, 
    1.975375e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975371e-24, 
    1.975369e-24, 1.975371e-24, 1.975368e-24, 1.97537e-24, 1.975369e-24, 
    1.975371e-24, 1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975378e-24, 
    1.975378e-24, 1.975379e-24, 1.97538e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 1.975377e-24, 
    1.975375e-24, 1.975376e-24, 1.975373e-24, 1.975374e-24, 1.975371e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 1.975378e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975377e-24, 
    1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975373e-24, 
    1.975371e-24, 1.975373e-24, 1.975373e-24, 1.975377e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975375e-24, 1.975376e-24, 1.975372e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 1.97537e-24, 
    1.975371e-24, 1.97537e-24, 1.975372e-24, 1.975371e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 1.975372e-24, 
    1.975373e-24, 1.975372e-24, 1.975373e-24, 1.975373e-24, 1.97537e-24, 
    1.975372e-24, 1.97537e-24, 1.97537e-24, 1.975371e-24, 1.97537e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975371e-24, 1.975372e-24, 1.97537e-24, 1.97537e-24, 1.97537e-24, 
    1.97537e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975375e-24, 1.975376e-24, 
    1.975375e-24, 1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975376e-24, 
    1.975373e-24, 1.975375e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.97537e-24, 1.975369e-24, 
    1.975369e-24, 1.975368e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975375e-24, 1.975374e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 
    1.975373e-24, 1.975374e-24, 1.975371e-24, 1.975372e-24, 1.975369e-24, 
    1.975368e-24, 1.975367e-24, 1.975365e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975377e-24, 1.975374e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975374e-24, 
    1.975368e-24, 1.975371e-24, 1.975365e-24, 1.975366e-24, 1.975378e-24, 
    1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975374e-24, 1.975373e-24, 
    1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975372e-24, 1.975374e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975368e-24, 1.975372e-24, 
    1.975377e-24, 1.975376e-24, 1.975376e-24, 1.975376e-24, 1.975373e-24, 
    1.975374e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975373e-24, 1.975374e-24, 1.975375e-24, 
    1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975374e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975375e-24, 1.975373e-24, 1.975375e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975373e-24, 1.975374e-24, 1.975374e-24, 1.975375e-24, 1.975375e-24, 
    1.975376e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975371e-24, 1.975371e-24, 1.975369e-24, 1.97537e-24, 1.975368e-24, 
    1.97537e-24, 1.975367e-24, 1.975372e-24, 1.97537e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 
    1.975374e-24, 1.975375e-24, 1.975375e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975374e-24, 
    1.975372e-24, 1.975371e-24, 1.975368e-24, 1.975367e-24, 1.975365e-24, 
    1.975365e-24, 1.975365e-24, 1.975364e-24 ;

 CONC_CH4_SAT =
  8.462784e-08, 8.473351e-08, 8.471293e-08, 8.479815e-08, 8.47508e-08, 
    8.480664e-08, 8.464917e-08, 8.47378e-08, 8.468118e-08, 8.463721e-08, 
    8.496334e-08, 8.480192e-08, 8.512928e-08, 8.502701e-08, 8.528312e-08, 
    8.511353e-08, 8.531718e-08, 8.527798e-08, 8.539523e-08, 8.536166e-08, 
    8.551176e-08, 8.541071e-08, 8.558894e-08, 8.548752e-08, 8.55035e-08, 
    8.540741e-08, 8.483422e-08, 8.494335e-08, 8.48278e-08, 8.484336e-08, 
    8.483633e-08, 8.475187e-08, 8.470941e-08, 8.461958e-08, 8.463585e-08, 
    8.470172e-08, 8.485036e-08, 8.47998e-08, 8.492663e-08, 8.492376e-08, 
    8.506463e-08, 8.500118e-08, 8.523705e-08, 8.517009e-08, 8.536306e-08, 
    8.531465e-08, 8.536083e-08, 8.534681e-08, 8.536101e-08, 8.528998e-08, 
    8.532044e-08, 8.525781e-08, 8.501312e-08, 8.508526e-08, 8.486983e-08, 
    8.474011e-08, 8.46531e-08, 8.459145e-08, 8.460017e-08, 8.461684e-08, 
    8.470212e-08, 8.478192e-08, 8.484272e-08, 8.488337e-08, 8.492335e-08, 
    8.504475e-08, 8.510831e-08, 8.525069e-08, 8.522483e-08, 8.526847e-08, 
    8.530983e-08, 8.537944e-08, 8.536796e-08, 8.539865e-08, 8.526717e-08, 
    8.535468e-08, 8.521013e-08, 8.524975e-08, 8.493505e-08, 8.481341e-08, 
    8.476232e-08, 8.471692e-08, 8.46069e-08, 8.468295e-08, 8.4653e-08, 
    8.472404e-08, 8.476923e-08, 8.474685e-08, 8.488448e-08, 8.483106e-08, 
    8.511208e-08, 8.499127e-08, 8.5305e-08, 8.523012e-08, 8.53229e-08, 
    8.527554e-08, 8.535672e-08, 8.528367e-08, 8.541e-08, 8.543755e-08, 
    8.541875e-08, 8.549066e-08, 8.527964e-08, 8.536091e-08, 8.474626e-08, 
    8.474992e-08, 8.476685e-08, 8.469239e-08, 8.468778e-08, 8.461917e-08, 
    8.468015e-08, 8.470616e-08, 8.477178e-08, 8.48107e-08, 8.484761e-08, 
    8.492864e-08, 8.501907e-08, 8.514493e-08, 8.523499e-08, 8.529528e-08, 
    8.525826e-08, 8.529095e-08, 8.525444e-08, 8.523728e-08, 8.542729e-08, 
    8.532078e-08, 8.548032e-08, 8.547148e-08, 8.539941e-08, 8.547248e-08, 
    8.475247e-08, 8.473145e-08, 8.465868e-08, 8.471564e-08, 8.461168e-08, 
    8.467001e-08, 8.470357e-08, 8.483236e-08, 8.48604e-08, 8.488664e-08, 
    8.493823e-08, 8.500444e-08, 8.512036e-08, 8.522083e-08, 8.531219e-08, 
    8.530549e-08, 8.530786e-08, 8.532833e-08, 8.527772e-08, 8.533663e-08, 
    8.534658e-08, 8.532066e-08, 8.54703e-08, 8.54276e-08, 8.54713e-08, 
    8.544348e-08, 8.473827e-08, 8.477357e-08, 8.475451e-08, 8.47904e-08, 
    8.476519e-08, 8.487742e-08, 8.491101e-08, 8.506756e-08, 8.500318e-08, 
    8.510537e-08, 8.50135e-08, 8.502985e-08, 8.510905e-08, 8.501842e-08, 
    8.521545e-08, 8.508229e-08, 8.532913e-08, 8.519686e-08, 8.533742e-08, 
    8.53118e-08, 8.535412e-08, 8.539208e-08, 8.543962e-08, 8.552744e-08, 
    8.550708e-08, 8.558028e-08, 8.482608e-08, 8.487186e-08, 8.486767e-08, 
    8.491541e-08, 8.495072e-08, 8.502693e-08, 8.514904e-08, 8.510312e-08, 
    8.518722e-08, 8.520414e-08, 8.507625e-08, 8.515497e-08, 8.490234e-08, 
    8.494343e-08, 8.491886e-08, 8.482979e-08, 8.511392e-08, 8.496846e-08, 
    8.52365e-08, 8.515797e-08, 8.538669e-08, 8.527327e-08, 8.549591e-08, 
    8.559111e-08, 8.567977e-08, 8.578395e-08, 8.489665e-08, 8.486558e-08, 
    8.492104e-08, 8.499792e-08, 8.506868e-08, 8.51628e-08, 8.517232e-08, 
    8.518997e-08, 8.523546e-08, 8.527375e-08, 8.519571e-08, 8.528333e-08, 
    8.495327e-08, 8.512645e-08, 8.485398e-08, 8.493645e-08, 8.499332e-08, 
    8.496822e-08, 8.509782e-08, 8.512836e-08, 8.525229e-08, 8.518818e-08, 
    8.556778e-08, 8.540031e-08, 8.586255e-08, 8.573405e-08, 8.485477e-08, 
    8.489646e-08, 8.504146e-08, 8.497252e-08, 8.516898e-08, 8.521727e-08, 
    8.525635e-08, 8.53065e-08, 8.531179e-08, 8.534145e-08, 8.529285e-08, 
    8.533947e-08, 8.516299e-08, 8.524193e-08, 8.502473e-08, 8.507779e-08, 
    8.505334e-08, 8.502661e-08, 8.510906e-08, 8.519698e-08, 8.51986e-08, 
    8.522679e-08, 8.530658e-08, 8.516977e-08, 8.55898e-08, 8.533137e-08, 
    8.49419e-08, 8.502234e-08, 8.503351e-08, 8.500243e-08, 8.521244e-08, 
    8.513651e-08, 8.534069e-08, 8.528556e-08, 8.537578e-08, 8.5331e-08, 
    8.532441e-08, 8.526674e-08, 8.523087e-08, 8.514004e-08, 8.506591e-08, 
    8.50069e-08, 8.502062e-08, 8.50854e-08, 8.520229e-08, 8.531238e-08, 
    8.528833e-08, 8.536893e-08, 8.515478e-08, 8.524485e-08, 8.521015e-08, 
    8.530053e-08, 8.510195e-08, 8.527188e-08, 8.505849e-08, 8.507719e-08, 
    8.513499e-08, 8.525112e-08, 8.527639e-08, 8.530381e-08, 8.528684e-08, 
    8.520521e-08, 8.51917e-08, 8.513353e-08, 8.511758e-08, 8.50731e-08, 
    8.503636e-08, 8.506999e-08, 8.510533e-08, 8.520514e-08, 8.5295e-08, 
    8.539266e-08, 8.541642e-08, 8.553077e-08, 8.543805e-08, 8.559129e-08, 
    8.546157e-08, 8.568557e-08, 8.528133e-08, 8.545724e-08, 8.513754e-08, 
    8.517204e-08, 8.523465e-08, 8.537732e-08, 8.53001e-08, 8.539028e-08, 
    8.519115e-08, 8.508776e-08, 8.506065e-08, 8.501054e-08, 8.506179e-08, 
    8.505761e-08, 8.510662e-08, 8.509087e-08, 8.520844e-08, 8.514532e-08, 
    8.532432e-08, 8.53895e-08, 8.55727e-08, 8.568473e-08, 8.579803e-08, 
    8.584807e-08, 8.586326e-08, 8.586963e-08,
  2.316417e-10, 2.322397e-10, 2.321232e-10, 2.326058e-10, 2.323377e-10, 
    2.32654e-10, 2.317625e-10, 2.322639e-10, 2.319435e-10, 2.316949e-10, 
    2.335471e-10, 2.326272e-10, 2.344984e-10, 2.339122e-10, 2.353819e-10, 
    2.344079e-10, 2.355778e-10, 2.353526e-10, 2.360272e-10, 2.358339e-10, 
    2.366984e-10, 2.361163e-10, 2.371439e-10, 2.365587e-10, 2.366508e-10, 
    2.360973e-10, 2.328104e-10, 2.334327e-10, 2.32774e-10, 2.328622e-10, 
    2.328223e-10, 2.323436e-10, 2.321031e-10, 2.315952e-10, 2.316872e-10, 
    2.320597e-10, 2.329018e-10, 2.326153e-10, 2.333376e-10, 2.333213e-10, 
    2.341278e-10, 2.337643e-10, 2.351173e-10, 2.347328e-10, 2.35842e-10, 
    2.355635e-10, 2.358291e-10, 2.357484e-10, 2.358302e-10, 2.354215e-10, 
    2.355967e-10, 2.352366e-10, 2.338326e-10, 2.34246e-10, 2.330129e-10, 
    2.322768e-10, 2.317847e-10, 2.314362e-10, 2.314855e-10, 2.315797e-10, 
    2.32062e-10, 2.32514e-10, 2.328586e-10, 2.330903e-10, 2.333189e-10, 
    2.340135e-10, 2.343781e-10, 2.351956e-10, 2.350471e-10, 2.352978e-10, 
    2.355357e-10, 2.359362e-10, 2.358702e-10, 2.360468e-10, 2.352904e-10, 
    2.357936e-10, 2.349628e-10, 2.351903e-10, 2.333852e-10, 2.326924e-10, 
    2.324026e-10, 2.321457e-10, 2.315235e-10, 2.319535e-10, 2.317841e-10, 
    2.321862e-10, 2.324421e-10, 2.323153e-10, 2.330967e-10, 2.327925e-10, 
    2.343997e-10, 2.337075e-10, 2.355079e-10, 2.350775e-10, 2.356109e-10, 
    2.353386e-10, 2.358054e-10, 2.353853e-10, 2.361122e-10, 2.362708e-10, 
    2.361625e-10, 2.36577e-10, 2.353621e-10, 2.358295e-10, 2.32312e-10, 
    2.323327e-10, 2.324286e-10, 2.320069e-10, 2.319809e-10, 2.315929e-10, 
    2.319377e-10, 2.320849e-10, 2.324566e-10, 2.326771e-10, 2.328863e-10, 
    2.333491e-10, 2.338666e-10, 2.345883e-10, 2.351055e-10, 2.35452e-10, 
    2.352393e-10, 2.354271e-10, 2.352173e-10, 2.351187e-10, 2.362116e-10, 
    2.355986e-10, 2.365174e-10, 2.364665e-10, 2.360512e-10, 2.364722e-10, 
    2.323471e-10, 2.322282e-10, 2.318162e-10, 2.321386e-10, 2.315506e-10, 
    2.318803e-10, 2.320701e-10, 2.327997e-10, 2.32959e-10, 2.33109e-10, 
    2.33404e-10, 2.33783e-10, 2.344473e-10, 2.350241e-10, 2.355494e-10, 
    2.355108e-10, 2.355244e-10, 2.356421e-10, 2.353511e-10, 2.356898e-10, 
    2.357471e-10, 2.35598e-10, 2.364597e-10, 2.362136e-10, 2.364654e-10, 
    2.363051e-10, 2.322667e-10, 2.324667e-10, 2.323587e-10, 2.32562e-10, 
    2.324191e-10, 2.330561e-10, 2.332481e-10, 2.341445e-10, 2.337757e-10, 
    2.343613e-10, 2.338349e-10, 2.339285e-10, 2.343821e-10, 2.338631e-10, 
    2.349931e-10, 2.342288e-10, 2.356467e-10, 2.348861e-10, 2.356944e-10, 
    2.355471e-10, 2.357906e-10, 2.36009e-10, 2.362828e-10, 2.367889e-10, 
    2.366716e-10, 2.370939e-10, 2.327643e-10, 2.330244e-10, 2.330006e-10, 
    2.332735e-10, 2.334754e-10, 2.339118e-10, 2.346119e-10, 2.343485e-10, 
    2.348312e-10, 2.349282e-10, 2.341945e-10, 2.346459e-10, 2.331987e-10, 
    2.334336e-10, 2.332932e-10, 2.327852e-10, 2.344103e-10, 2.335768e-10, 
    2.351142e-10, 2.346632e-10, 2.359779e-10, 2.353253e-10, 2.366072e-10, 
    2.371562e-10, 2.376686e-10, 2.38271e-10, 2.331662e-10, 2.329887e-10, 
    2.333057e-10, 2.337455e-10, 2.34151e-10, 2.346909e-10, 2.347456e-10, 
    2.348469e-10, 2.351083e-10, 2.353283e-10, 2.348797e-10, 2.353834e-10, 
    2.334896e-10, 2.344822e-10, 2.329224e-10, 2.333936e-10, 2.337192e-10, 
    2.335756e-10, 2.343182e-10, 2.344934e-10, 2.352048e-10, 2.348367e-10, 
    2.370214e-10, 2.360562e-10, 2.387265e-10, 2.379824e-10, 2.32927e-10, 
    2.331652e-10, 2.33995e-10, 2.336002e-10, 2.347265e-10, 2.350037e-10, 
    2.352283e-10, 2.355164e-10, 2.35547e-10, 2.357175e-10, 2.354381e-10, 
    2.357062e-10, 2.34692e-10, 2.351454e-10, 2.338993e-10, 2.342033e-10, 
    2.340632e-10, 2.3391e-10, 2.343827e-10, 2.34887e-10, 2.348965e-10, 
    2.350583e-10, 2.355163e-10, 2.34731e-10, 2.371482e-10, 2.35659e-10, 
    2.33425e-10, 2.338853e-10, 2.339495e-10, 2.337715e-10, 2.34976e-10, 
    2.3454e-10, 2.357132e-10, 2.353961e-10, 2.359152e-10, 2.356574e-10, 
    2.356196e-10, 2.35288e-10, 2.350818e-10, 2.345603e-10, 2.341352e-10, 
    2.337972e-10, 2.338757e-10, 2.342468e-10, 2.349175e-10, 2.355503e-10, 
    2.354119e-10, 2.358758e-10, 2.346449e-10, 2.351621e-10, 2.349627e-10, 
    2.354822e-10, 2.343418e-10, 2.353169e-10, 2.340927e-10, 2.341999e-10, 
    2.345313e-10, 2.35198e-10, 2.353435e-10, 2.35501e-10, 2.354036e-10, 
    2.349343e-10, 2.348568e-10, 2.34523e-10, 2.344314e-10, 2.341765e-10, 
    2.339659e-10, 2.341586e-10, 2.343612e-10, 2.34934e-10, 2.354504e-10, 
    2.360123e-10, 2.361492e-10, 2.368079e-10, 2.362734e-10, 2.371567e-10, 
    2.364085e-10, 2.377017e-10, 2.353714e-10, 2.363839e-10, 2.34546e-10, 
    2.34744e-10, 2.351034e-10, 2.359238e-10, 2.354797e-10, 2.359984e-10, 
    2.348537e-10, 2.342603e-10, 2.341051e-10, 2.33818e-10, 2.341116e-10, 
    2.340877e-10, 2.343687e-10, 2.342783e-10, 2.34953e-10, 2.345906e-10, 
    2.356189e-10, 2.35994e-10, 2.370501e-10, 2.376971e-10, 2.383528e-10, 
    2.386426e-10, 2.387307e-10, 2.387676e-10,
  1.287514e-13, 1.292006e-13, 1.291131e-13, 1.294758e-13, 1.292743e-13, 
    1.29512e-13, 1.288421e-13, 1.292187e-13, 1.289781e-13, 1.287914e-13, 
    1.30183e-13, 1.294919e-13, 1.308989e-13, 1.304579e-13, 1.315645e-13, 
    1.308307e-13, 1.317148e-13, 1.315426e-13, 1.320633e-13, 1.319135e-13, 
    1.325839e-13, 1.321325e-13, 1.3293e-13, 1.324756e-13, 1.32547e-13, 
    1.321177e-13, 1.296297e-13, 1.300971e-13, 1.296023e-13, 1.296687e-13, 
    1.296387e-13, 1.292787e-13, 1.290978e-13, 1.287165e-13, 1.287856e-13, 
    1.290654e-13, 1.296985e-13, 1.29483e-13, 1.30026e-13, 1.300137e-13, 
    1.306201e-13, 1.303467e-13, 1.313652e-13, 1.310756e-13, 1.319197e-13, 
    1.317038e-13, 1.319097e-13, 1.318472e-13, 1.319105e-13, 1.315946e-13, 
    1.317296e-13, 1.314552e-13, 1.303981e-13, 1.30709e-13, 1.29782e-13, 
    1.292283e-13, 1.288588e-13, 1.285972e-13, 1.286342e-13, 1.287048e-13, 
    1.29067e-13, 1.294069e-13, 1.296661e-13, 1.298402e-13, 1.300119e-13, 
    1.305339e-13, 1.308083e-13, 1.314242e-13, 1.313124e-13, 1.315012e-13, 
    1.316823e-13, 1.319928e-13, 1.319415e-13, 1.320785e-13, 1.314957e-13, 
    1.318821e-13, 1.312488e-13, 1.314203e-13, 1.300613e-13, 1.29541e-13, 
    1.293229e-13, 1.2913e-13, 1.286626e-13, 1.289855e-13, 1.288583e-13, 
    1.291604e-13, 1.293528e-13, 1.292575e-13, 1.298449e-13, 1.296163e-13, 
    1.308246e-13, 1.303039e-13, 1.316608e-13, 1.313353e-13, 1.317406e-13, 
    1.315321e-13, 1.318913e-13, 1.315673e-13, 1.321292e-13, 1.322522e-13, 
    1.321682e-13, 1.324899e-13, 1.315498e-13, 1.3191e-13, 1.29255e-13, 
    1.292705e-13, 1.293427e-13, 1.290256e-13, 1.290061e-13, 1.287148e-13, 
    1.289737e-13, 1.290843e-13, 1.293637e-13, 1.295295e-13, 1.296869e-13, 
    1.300346e-13, 1.304236e-13, 1.309666e-13, 1.313563e-13, 1.316176e-13, 
    1.314572e-13, 1.315988e-13, 1.314406e-13, 1.313663e-13, 1.322063e-13, 
    1.31731e-13, 1.324436e-13, 1.324041e-13, 1.320818e-13, 1.324085e-13, 
    1.292814e-13, 1.29192e-13, 1.288825e-13, 1.291247e-13, 1.28683e-13, 
    1.289306e-13, 1.290731e-13, 1.296216e-13, 1.297416e-13, 1.298542e-13, 
    1.300759e-13, 1.303607e-13, 1.308605e-13, 1.312949e-13, 1.316929e-13, 
    1.316631e-13, 1.316736e-13, 1.317648e-13, 1.315415e-13, 1.318018e-13, 
    1.318461e-13, 1.317306e-13, 1.323988e-13, 1.322079e-13, 1.324033e-13, 
    1.322789e-13, 1.29221e-13, 1.293713e-13, 1.292901e-13, 1.294429e-13, 
    1.293355e-13, 1.298144e-13, 1.299586e-13, 1.306325e-13, 1.303553e-13, 
    1.307958e-13, 1.303998e-13, 1.304701e-13, 1.308113e-13, 1.30421e-13, 
    1.312715e-13, 1.306959e-13, 1.317683e-13, 1.311908e-13, 1.318053e-13, 
    1.316912e-13, 1.318799e-13, 1.320491e-13, 1.322616e-13, 1.326544e-13, 
    1.325633e-13, 1.328913e-13, 1.295951e-13, 1.297906e-13, 1.297728e-13, 
    1.299778e-13, 1.301295e-13, 1.304577e-13, 1.309845e-13, 1.307862e-13, 
    1.311497e-13, 1.312228e-13, 1.306704e-13, 1.3101e-13, 1.299215e-13, 
    1.300979e-13, 1.299925e-13, 1.296108e-13, 1.308326e-13, 1.302056e-13, 
    1.313628e-13, 1.310231e-13, 1.320251e-13, 1.315219e-13, 1.325133e-13, 
    1.329395e-13, 1.333381e-13, 1.338066e-13, 1.298971e-13, 1.297639e-13, 
    1.30002e-13, 1.303324e-13, 1.306376e-13, 1.31044e-13, 1.310853e-13, 
    1.311615e-13, 1.313585e-13, 1.315243e-13, 1.311861e-13, 1.315658e-13, 
    1.301398e-13, 1.308868e-13, 1.29714e-13, 1.300678e-13, 1.303128e-13, 
    1.302048e-13, 1.307635e-13, 1.308953e-13, 1.314311e-13, 1.311538e-13, 
    1.328347e-13, 1.320856e-13, 1.341616e-13, 1.33582e-13, 1.297175e-13, 
    1.298964e-13, 1.305201e-13, 1.302233e-13, 1.310708e-13, 1.312796e-13, 
    1.314489e-13, 1.316674e-13, 1.316911e-13, 1.318232e-13, 1.316071e-13, 
    1.318145e-13, 1.310448e-13, 1.313864e-13, 1.304483e-13, 1.306769e-13, 
    1.305716e-13, 1.304563e-13, 1.308119e-13, 1.311916e-13, 1.311989e-13, 
    1.313207e-13, 1.316668e-13, 1.310742e-13, 1.32933e-13, 1.317774e-13, 
    1.300917e-13, 1.304376e-13, 1.30486e-13, 1.303522e-13, 1.312587e-13, 
    1.309304e-13, 1.318199e-13, 1.315754e-13, 1.319765e-13, 1.317767e-13, 
    1.317473e-13, 1.314939e-13, 1.313385e-13, 1.309456e-13, 1.306256e-13, 
    1.303715e-13, 1.304305e-13, 1.307097e-13, 1.312146e-13, 1.316936e-13, 
    1.315873e-13, 1.319459e-13, 1.310094e-13, 1.313989e-13, 1.312486e-13, 
    1.316409e-13, 1.307811e-13, 1.315153e-13, 1.305938e-13, 1.306744e-13, 
    1.309238e-13, 1.314259e-13, 1.315357e-13, 1.316554e-13, 1.31581e-13, 
    1.312273e-13, 1.31169e-13, 1.309176e-13, 1.308486e-13, 1.306568e-13, 
    1.304984e-13, 1.306433e-13, 1.307957e-13, 1.312271e-13, 1.316163e-13, 
    1.320517e-13, 1.321579e-13, 1.326688e-13, 1.322541e-13, 1.329395e-13, 
    1.323585e-13, 1.333634e-13, 1.315566e-13, 1.323397e-13, 1.309349e-13, 
    1.310841e-13, 1.313546e-13, 1.31983e-13, 1.31639e-13, 1.320409e-13, 
    1.311666e-13, 1.307197e-13, 1.306031e-13, 1.303871e-13, 1.30608e-13, 
    1.3059e-13, 1.308014e-13, 1.307334e-13, 1.312414e-13, 1.309685e-13, 
    1.317468e-13, 1.320375e-13, 1.328572e-13, 1.333601e-13, 1.338705e-13, 
    1.340963e-13, 1.341649e-13, 1.341937e-13,
  1.866922e-17, 1.87439e-17, 1.872935e-17, 1.878968e-17, 1.875617e-17, 
    1.879571e-17, 1.868431e-17, 1.874691e-17, 1.870692e-17, 1.867588e-17, 
    1.890713e-17, 1.879236e-17, 1.90261e-17, 1.895283e-17, 1.913685e-17, 
    1.901476e-17, 1.916251e-17, 1.913321e-17, 1.922275e-17, 1.919686e-17, 
    1.931273e-17, 1.92347e-17, 1.937267e-17, 1.929403e-17, 1.930637e-17, 
    1.923215e-17, 1.881532e-17, 1.889286e-17, 1.881076e-17, 1.882179e-17, 
    1.881682e-17, 1.87569e-17, 1.872679e-17, 1.866345e-17, 1.867492e-17, 
    1.872141e-17, 1.882675e-17, 1.879091e-17, 1.888113e-17, 1.887909e-17, 
    1.897978e-17, 1.893437e-17, 1.910369e-17, 1.905551e-17, 1.919793e-17, 
    1.916063e-17, 1.91962e-17, 1.91854e-17, 1.919634e-17, 1.914187e-17, 
    1.916508e-17, 1.911867e-17, 1.89429e-17, 1.899456e-17, 1.884062e-17, 
    1.874848e-17, 1.868708e-17, 1.864361e-17, 1.864975e-17, 1.866149e-17, 
    1.872168e-17, 1.877823e-17, 1.882138e-17, 1.88503e-17, 1.88788e-17, 
    1.896541e-17, 1.901105e-17, 1.911349e-17, 1.90949e-17, 1.912632e-17, 
    1.915692e-17, 1.921055e-17, 1.92017e-17, 1.922536e-17, 1.912542e-17, 
    1.919143e-17, 1.908434e-17, 1.911286e-17, 1.888692e-17, 1.880056e-17, 
    1.876423e-17, 1.873216e-17, 1.865448e-17, 1.870814e-17, 1.868699e-17, 
    1.873724e-17, 1.876923e-17, 1.875339e-17, 1.885109e-17, 1.881309e-17, 
    1.901376e-17, 1.892725e-17, 1.91532e-17, 1.909871e-17, 1.916699e-17, 
    1.913147e-17, 1.919302e-17, 1.913733e-17, 1.923413e-17, 1.925538e-17, 
    1.924087e-17, 1.929651e-17, 1.913442e-17, 1.919624e-17, 1.875296e-17, 
    1.875555e-17, 1.876755e-17, 1.871481e-17, 1.871156e-17, 1.866315e-17, 
    1.870619e-17, 1.872456e-17, 1.877105e-17, 1.879864e-17, 1.882484e-17, 
    1.888255e-17, 1.894712e-17, 1.903738e-17, 1.910221e-17, 1.914575e-17, 
    1.911901e-17, 1.914259e-17, 1.911625e-17, 1.910389e-17, 1.924745e-17, 
    1.916532e-17, 1.92885e-17, 1.928167e-17, 1.922594e-17, 1.928244e-17, 
    1.875736e-17, 1.874249e-17, 1.869102e-17, 1.87313e-17, 1.865787e-17, 
    1.869901e-17, 1.87227e-17, 1.881396e-17, 1.883394e-17, 1.885261e-17, 
    1.888941e-17, 1.89367e-17, 1.901974e-17, 1.909199e-17, 1.915876e-17, 
    1.91536e-17, 1.915542e-17, 1.917116e-17, 1.913303e-17, 1.917755e-17, 
    1.91852e-17, 1.916527e-17, 1.928076e-17, 1.924774e-17, 1.928153e-17, 
    1.926002e-17, 1.874731e-17, 1.877231e-17, 1.875881e-17, 1.878422e-17, 
    1.876635e-17, 1.884599e-17, 1.886991e-17, 1.898183e-17, 1.893579e-17, 
    1.900897e-17, 1.894319e-17, 1.895486e-17, 1.901151e-17, 1.894672e-17, 
    1.908808e-17, 1.899236e-17, 1.917177e-17, 1.907464e-17, 1.917816e-17, 
    1.915845e-17, 1.919105e-17, 1.922029e-17, 1.925702e-17, 1.932495e-17, 
    1.93092e-17, 1.936597e-17, 1.880956e-17, 1.884206e-17, 1.883912e-17, 
    1.887313e-17, 1.88983e-17, 1.89528e-17, 1.904036e-17, 1.90074e-17, 
    1.906784e-17, 1.908e-17, 1.898815e-17, 1.90446e-17, 1.886378e-17, 
    1.889304e-17, 1.887557e-17, 1.881216e-17, 1.901509e-17, 1.891092e-17, 
    1.91033e-17, 1.904679e-17, 1.921613e-17, 1.912977e-17, 1.930055e-17, 
    1.937428e-17, 1.944338e-17, 1.952459e-17, 1.885974e-17, 1.883764e-17, 
    1.887715e-17, 1.893198e-17, 1.898269e-17, 1.905025e-17, 1.905712e-17, 
    1.906981e-17, 1.910258e-17, 1.913018e-17, 1.907388e-17, 1.913709e-17, 
    1.889997e-17, 1.902411e-17, 1.882935e-17, 1.888805e-17, 1.892872e-17, 
    1.89108e-17, 1.900362e-17, 1.902553e-17, 1.911465e-17, 1.906853e-17, 
    1.935614e-17, 1.922657e-17, 1.958622e-17, 1.948564e-17, 1.882994e-17, 
    1.885963e-17, 1.896317e-17, 1.891388e-17, 1.905472e-17, 1.908945e-17, 
    1.911763e-17, 1.915433e-17, 1.915843e-17, 1.918125e-17, 1.914396e-17, 
    1.917975e-17, 1.905039e-17, 1.910723e-17, 1.895124e-17, 1.898923e-17, 
    1.897173e-17, 1.895259e-17, 1.901168e-17, 1.907479e-17, 1.907602e-17, 
    1.909629e-17, 1.915413e-17, 1.905529e-17, 1.937309e-17, 1.917326e-17, 
    1.889203e-17, 1.894944e-17, 1.89575e-17, 1.893528e-17, 1.908597e-17, 
    1.903136e-17, 1.918068e-17, 1.91387e-17, 1.920774e-17, 1.917322e-17, 
    1.916815e-17, 1.912512e-17, 1.909925e-17, 1.903389e-17, 1.89807e-17, 
    1.893849e-17, 1.89483e-17, 1.899467e-17, 1.907862e-17, 1.915886e-17, 
    1.914065e-17, 1.920246e-17, 1.904451e-17, 1.91093e-17, 1.908429e-17, 
    1.914976e-17, 1.900655e-17, 1.91286e-17, 1.897542e-17, 1.898882e-17, 
    1.903028e-17, 1.911377e-17, 1.913208e-17, 1.915227e-17, 1.913963e-17, 
    1.908073e-17, 1.907104e-17, 1.902924e-17, 1.901776e-17, 1.898589e-17, 
    1.895957e-17, 1.898365e-17, 1.900896e-17, 1.908071e-17, 1.91455e-17, 
    1.922073e-17, 1.92391e-17, 1.93274e-17, 1.925568e-17, 1.937423e-17, 
    1.927367e-17, 1.944768e-17, 1.913551e-17, 1.927048e-17, 1.903213e-17, 
    1.905692e-17, 1.910191e-17, 1.920882e-17, 1.914943e-17, 1.921884e-17, 
    1.907065e-17, 1.899632e-17, 1.897696e-17, 1.894108e-17, 1.897778e-17, 
    1.897479e-17, 1.900993e-17, 1.899863e-17, 1.908309e-17, 1.903771e-17, 
    1.916805e-17, 1.921826e-17, 1.936006e-17, 1.944717e-17, 1.953572e-17, 
    1.95749e-17, 1.958682e-17, 1.959181e-17,
  7.811738e-22, 7.847107e-22, 7.840216e-22, 7.868805e-22, 7.852925e-22, 
    7.871665e-22, 7.818885e-22, 7.848529e-22, 7.829589e-22, 7.814895e-22, 
    7.924481e-22, 7.870076e-22, 7.980991e-22, 7.946196e-22, 8.033665e-22, 
    7.975596e-22, 8.045871e-22, 8.031944e-22, 8.074501e-22, 8.062195e-22, 
    8.117452e-22, 8.080182e-22, 8.14689e-22, 8.108386e-22, 8.114337e-22, 
    8.078967e-22, 7.880969e-22, 7.917711e-22, 7.878805e-22, 7.884035e-22, 
    7.881679e-22, 7.853267e-22, 7.838993e-22, 7.80901e-22, 7.814442e-22, 
    7.83645e-22, 7.886387e-22, 7.869393e-22, 7.91218e-22, 7.911211e-22, 
    7.958995e-22, 7.937436e-22, 8.017896e-22, 7.994984e-22, 8.062708e-22, 
    8.044988e-22, 8.061882e-22, 8.056752e-22, 8.061949e-22, 8.036063e-22, 
    8.047097e-22, 8.025023e-22, 7.94148e-22, 7.96601e-22, 7.892968e-22, 
    7.849263e-22, 7.820192e-22, 7.799621e-22, 7.802528e-22, 7.808079e-22, 
    7.83658e-22, 7.863382e-22, 7.883846e-22, 7.897557e-22, 7.911072e-22, 
    7.952153e-22, 7.973838e-22, 8.022552e-22, 8.013716e-22, 8.028659e-22, 
    8.043224e-22, 8.068698e-22, 8.064497e-22, 8.075737e-22, 8.028239e-22, 
    8.059609e-22, 8.008694e-22, 8.022257e-22, 7.914891e-22, 7.873969e-22, 
    7.856729e-22, 7.841545e-22, 7.804766e-22, 7.830165e-22, 7.820152e-22, 
    7.843954e-22, 7.859114e-22, 7.851609e-22, 7.897931e-22, 7.879912e-22, 
    7.975125e-22, 7.934052e-22, 8.041459e-22, 8.015527e-22, 8.048007e-22, 
    8.031119e-22, 8.060367e-22, 8.033908e-22, 8.07991e-22, 8.090008e-22, 
    8.08311e-22, 8.109572e-22, 8.03252e-22, 8.061896e-22, 7.851405e-22, 
    7.85263e-22, 7.85832e-22, 7.833322e-22, 7.831786e-22, 7.808868e-22, 
    7.829246e-22, 7.837943e-22, 7.859982e-22, 7.873057e-22, 7.885485e-22, 
    7.912849e-22, 7.943481e-22, 7.986356e-22, 8.017194e-22, 8.037919e-22, 
    8.02519e-22, 8.03641e-22, 8.023874e-22, 8.017994e-22, 8.086234e-22, 
    8.047209e-22, 8.105764e-22, 8.102514e-22, 8.07601e-22, 8.10288e-22, 
    7.853487e-22, 7.846445e-22, 7.82206e-22, 7.84114e-22, 7.806372e-22, 
    7.825843e-22, 7.837058e-22, 7.880319e-22, 7.889803e-22, 7.89865e-22, 
    7.916102e-22, 7.93854e-22, 7.977974e-22, 8.012326e-22, 8.044099e-22, 
    8.04165e-22, 8.042513e-22, 8.049988e-22, 8.03186e-22, 8.053023e-22, 
    8.056651e-22, 8.047187e-22, 8.10208e-22, 8.08638e-22, 8.102445e-22, 
    8.092217e-22, 7.84873e-22, 7.860577e-22, 7.854176e-22, 7.866221e-22, 
    7.857746e-22, 7.895505e-22, 7.906844e-22, 7.959957e-22, 7.938106e-22, 
    7.972854e-22, 7.941622e-22, 7.94716e-22, 7.974049e-22, 7.943299e-22, 
    8.010458e-22, 7.964955e-22, 8.050278e-22, 8.004059e-22, 8.053313e-22, 
    8.043954e-22, 8.059437e-22, 8.073329e-22, 8.090793e-22, 8.123461e-22, 
    8.115734e-22, 8.143607e-22, 7.878238e-22, 7.893645e-22, 7.892261e-22, 
    7.908383e-22, 7.92032e-22, 7.946187e-22, 7.987776e-22, 7.972118e-22, 
    8.000844e-22, 8.006626e-22, 7.962971e-22, 7.989789e-22, 7.903946e-22, 
    7.917817e-22, 7.909537e-22, 7.879468e-22, 7.975762e-22, 7.926297e-22, 
    8.017709e-22, 7.990834e-22, 8.071352e-22, 8.030298e-22, 8.111491e-22, 
    8.14767e-22, 8.181651e-22, 8.221589e-22, 7.902032e-22, 7.891557e-22, 
    7.910293e-22, 7.936294e-22, 7.960375e-22, 7.992478e-22, 7.99575e-22, 
    8.001779e-22, 8.01737e-22, 8.030502e-22, 8.003711e-22, 8.033793e-22, 
    7.921088e-22, 7.980049e-22, 7.887624e-22, 7.915444e-22, 7.934749e-22, 
    7.926251e-22, 7.970322e-22, 7.980733e-22, 8.023107e-22, 8.001175e-22, 
    8.138759e-22, 8.076304e-22, 8.251956e-22, 8.202422e-22, 7.887906e-22, 
    7.901984e-22, 7.9511e-22, 7.92771e-22, 7.994608e-22, 8.011122e-22, 
    8.024532e-22, 8.04199e-22, 8.043944e-22, 8.054778e-22, 8.037065e-22, 
    8.054066e-22, 7.992546e-22, 8.019578e-22, 7.945447e-22, 7.96348e-22, 
    7.955173e-22, 7.946086e-22, 7.974151e-22, 8.00414e-22, 8.004737e-22, 
    8.014371e-22, 8.041864e-22, 7.994878e-22, 8.147061e-22, 8.050951e-22, 
    7.917349e-22, 7.944577e-22, 7.948416e-22, 7.937871e-22, 8.009467e-22, 
    7.983501e-22, 8.054508e-22, 8.034557e-22, 8.067368e-22, 8.050965e-22, 
    8.048555e-22, 8.028097e-22, 8.015784e-22, 7.984699e-22, 7.959431e-22, 
    7.939395e-22, 7.944048e-22, 7.966063e-22, 8.005965e-22, 8.044141e-22, 
    8.035478e-22, 8.064857e-22, 7.989751e-22, 8.02056e-22, 8.008661e-22, 
    8.039824e-22, 7.971711e-22, 8.029719e-22, 7.956927e-22, 7.963289e-22, 
    7.982985e-22, 8.022681e-22, 8.031409e-22, 8.041011e-22, 8.035e-22, 
    8.006971e-22, 8.002364e-22, 7.982496e-22, 7.977035e-22, 7.961901e-22, 
    7.9494e-22, 7.960832e-22, 7.972853e-22, 8.006965e-22, 8.037794e-22, 
    8.073534e-22, 8.082274e-22, 8.124644e-22, 8.090134e-22, 8.147617e-22, 
    8.098664e-22, 8.183733e-22, 8.033021e-22, 8.097169e-22, 7.983867e-22, 
    7.995655e-22, 8.017042e-22, 8.067869e-22, 8.039668e-22, 8.07263e-22, 
    8.00218e-22, 7.966844e-22, 7.957659e-22, 7.94062e-22, 7.958048e-22, 
    7.956628e-22, 7.973321e-22, 7.967953e-22, 8.008098e-22, 7.986522e-22, 
    8.048506e-22, 8.072358e-22, 8.1407e-22, 8.183499e-22, 8.227086e-22, 
    8.246382e-22, 8.252254e-22, 8.254712e-22,
  1.00598e-26, 1.011182e-26, 1.010168e-26, 1.014375e-26, 1.012038e-26, 
    1.014797e-26, 1.007031e-26, 1.01139e-26, 1.008605e-26, 1.006445e-26, 
    1.022578e-26, 1.014563e-26, 1.030924e-26, 1.025786e-26, 1.038717e-26, 
    1.030127e-26, 1.040502e-26, 1.038464e-26, 1.044663e-26, 1.042875e-26, 
    1.050919e-26, 1.045489e-26, 1.055257e-26, 1.049591e-26, 1.050461e-26, 
    1.045312e-26, 1.016168e-26, 1.02158e-26, 1.015849e-26, 1.016619e-26, 
    1.016272e-26, 1.012088e-26, 1.009987e-26, 1.00558e-26, 1.006378e-26, 
    1.009614e-26, 1.016965e-26, 1.014463e-26, 1.020768e-26, 1.020625e-26, 
    1.027676e-26, 1.024493e-26, 1.036384e-26, 1.032995e-26, 1.042949e-26, 
    1.040374e-26, 1.042829e-26, 1.042084e-26, 1.042839e-26, 1.039073e-26, 
    1.040681e-26, 1.037439e-26, 1.02509e-26, 1.028711e-26, 1.017935e-26, 
    1.011497e-26, 1.007223e-26, 1.0042e-26, 1.004627e-26, 1.005443e-26, 
    1.009633e-26, 1.013578e-26, 1.016592e-26, 1.018612e-26, 1.020605e-26, 
    1.026663e-26, 1.029867e-26, 1.037072e-26, 1.035766e-26, 1.037977e-26, 
    1.040118e-26, 1.043819e-26, 1.043209e-26, 1.044843e-26, 1.037915e-26, 
    1.042498e-26, 1.035023e-26, 1.03703e-26, 1.021163e-26, 1.015137e-26, 
    1.012596e-26, 1.010363e-26, 1.004956e-26, 1.008689e-26, 1.007217e-26, 
    1.010718e-26, 1.012949e-26, 1.011845e-26, 1.018667e-26, 1.016012e-26, 
    1.030058e-26, 1.023993e-26, 1.039862e-26, 1.036033e-26, 1.040813e-26, 
    1.038342e-26, 1.042608e-26, 1.038755e-26, 1.045449e-26, 1.046917e-26, 
    1.045915e-26, 1.049764e-26, 1.038549e-26, 1.042831e-26, 1.011815e-26, 
    1.011995e-26, 1.012833e-26, 1.009153e-26, 1.008928e-26, 1.005559e-26, 
    1.008555e-26, 1.009833e-26, 1.013077e-26, 1.015002e-26, 1.016833e-26, 
    1.020866e-26, 1.025384e-26, 1.031718e-26, 1.03628e-26, 1.039348e-26, 
    1.037464e-26, 1.039125e-26, 1.037269e-26, 1.036399e-26, 1.046368e-26, 
    1.040697e-26, 1.04921e-26, 1.048737e-26, 1.044882e-26, 1.048791e-26, 
    1.012121e-26, 1.011085e-26, 1.007498e-26, 1.010304e-26, 1.005192e-26, 
    1.008054e-26, 1.009703e-26, 1.016071e-26, 1.01747e-26, 1.018773e-26, 
    1.021346e-26, 1.024656e-26, 1.030479e-26, 1.035559e-26, 1.040246e-26, 
    1.03989e-26, 1.040015e-26, 1.041101e-26, 1.038451e-26, 1.041542e-26, 
    1.042068e-26, 1.040694e-26, 1.048674e-26, 1.046391e-26, 1.048727e-26, 
    1.04724e-26, 1.011421e-26, 1.013165e-26, 1.012223e-26, 1.013995e-26, 
    1.012748e-26, 1.018309e-26, 1.01998e-26, 1.027817e-26, 1.024592e-26, 
    1.029723e-26, 1.025111e-26, 1.025928e-26, 1.029897e-26, 1.025359e-26, 
    1.035282e-26, 1.028554e-26, 1.041143e-26, 1.034335e-26, 1.041584e-26, 
    1.040225e-26, 1.042474e-26, 1.044493e-26, 1.047032e-26, 1.051806e-26, 
    1.050668e-26, 1.054774e-26, 1.015766e-26, 1.018035e-26, 1.017832e-26, 
    1.020208e-26, 1.021968e-26, 1.025785e-26, 1.031929e-26, 1.029615e-26, 
    1.033862e-26, 1.034716e-26, 1.028263e-26, 1.032226e-26, 1.019553e-26, 
    1.021598e-26, 1.020378e-26, 1.015946e-26, 1.030152e-26, 1.022848e-26, 
    1.036356e-26, 1.032381e-26, 1.044205e-26, 1.038219e-26, 1.050043e-26, 
    1.055371e-26, 1.060513e-26, 1.066582e-26, 1.019272e-26, 1.017728e-26, 
    1.02049e-26, 1.024324e-26, 1.02788e-26, 1.032624e-26, 1.033108e-26, 
    1.033999e-26, 1.036307e-26, 1.03825e-26, 1.034284e-26, 1.038738e-26, 
    1.022078e-26, 1.030786e-26, 1.017148e-26, 1.021247e-26, 1.024096e-26, 
    1.022843e-26, 1.02935e-26, 1.030888e-26, 1.037155e-26, 1.03391e-26, 
    1.054057e-26, 1.044924e-26, 1.071205e-26, 1.063667e-26, 1.01719e-26, 
    1.019265e-26, 1.026509e-26, 1.023058e-26, 1.032939e-26, 1.035381e-26, 
    1.037367e-26, 1.039939e-26, 1.040223e-26, 1.041797e-26, 1.039222e-26, 
    1.041693e-26, 1.032634e-26, 1.036633e-26, 1.025676e-26, 1.028338e-26, 
    1.027112e-26, 1.02577e-26, 1.029915e-26, 1.034348e-26, 1.034437e-26, 
    1.035862e-26, 1.039916e-26, 1.032979e-26, 1.055278e-26, 1.041237e-26, 
    1.02153e-26, 1.025546e-26, 1.026114e-26, 1.024558e-26, 1.035137e-26, 
    1.031297e-26, 1.041757e-26, 1.038851e-26, 1.043626e-26, 1.041243e-26, 
    1.040893e-26, 1.037894e-26, 1.036071e-26, 1.031473e-26, 1.02774e-26, 
    1.024783e-26, 1.025469e-26, 1.02872e-26, 1.034618e-26, 1.040251e-26, 
    1.038986e-26, 1.043261e-26, 1.032221e-26, 1.036778e-26, 1.035017e-26, 
    1.039625e-26, 1.029554e-26, 1.03813e-26, 1.027371e-26, 1.02831e-26, 
    1.03122e-26, 1.037091e-26, 1.038385e-26, 1.039796e-26, 1.038916e-26, 
    1.034767e-26, 1.034086e-26, 1.031148e-26, 1.030341e-26, 1.028105e-26, 
    1.02626e-26, 1.027947e-26, 1.029723e-26, 1.034767e-26, 1.039329e-26, 
    1.044522e-26, 1.045793e-26, 1.051978e-26, 1.046934e-26, 1.05536e-26, 
    1.048172e-26, 1.060825e-26, 1.038621e-26, 1.047957e-26, 1.031351e-26, 
    1.033094e-26, 1.036256e-26, 1.043697e-26, 1.039602e-26, 1.04439e-26, 
    1.034059e-26, 1.028834e-26, 1.027479e-26, 1.024963e-26, 1.027536e-26, 
    1.027327e-26, 1.029793e-26, 1.029e-26, 1.034934e-26, 1.031744e-26, 
    1.040885e-26, 1.044351e-26, 1.054345e-26, 1.060792e-26, 1.06742e-26, 
    1.070357e-26, 1.071252e-26, 1.071626e-26,
  4.063717e-32, 4.088939e-32, 4.084022e-32, 4.104447e-32, 4.0931e-32, 
    4.106493e-32, 4.068812e-32, 4.08995e-32, 4.076442e-32, 4.065971e-32, 
    4.144812e-32, 4.105358e-32, 4.186733e-32, 4.16092e-32, 4.225985e-32, 
    4.182718e-32, 4.234887e-32, 4.224713e-32, 4.255546e-32, 4.246665e-32, 
    4.286594e-32, 4.259649e-32, 4.307971e-32, 4.280037e-32, 4.284342e-32, 
    4.25877e-32, 4.113161e-32, 4.139807e-32, 4.111611e-32, 4.115353e-32, 
    4.11367e-32, 4.09334e-32, 4.083138e-32, 4.061782e-32, 4.065649e-32, 
    4.081331e-32, 4.117036e-32, 4.104876e-32, 4.135761e-32, 4.135045e-32, 
    4.170411e-32, 4.154435e-32, 4.214227e-32, 4.197159e-32, 4.247036e-32, 
    4.234261e-32, 4.246438e-32, 4.24274e-32, 4.246486e-32, 4.227789e-32, 
    4.235778e-32, 4.219547e-32, 4.157427e-32, 4.175612e-32, 4.121755e-32, 
    4.090464e-32, 4.069741e-32, 4.0551e-32, 4.057167e-32, 4.061114e-32, 
    4.081423e-32, 4.100576e-32, 4.115225e-32, 4.125051e-32, 4.134943e-32, 
    4.165312e-32, 4.181418e-32, 4.217694e-32, 4.211113e-32, 4.222254e-32, 
    4.232991e-32, 4.251354e-32, 4.248325e-32, 4.256434e-32, 4.221948e-32, 
    4.244793e-32, 4.207372e-32, 4.217483e-32, 4.13772e-32, 4.108151e-32, 
    4.095801e-32, 4.084969e-32, 4.058758e-32, 4.076848e-32, 4.069711e-32, 
    4.086694e-32, 4.097524e-32, 4.092162e-32, 4.12532e-32, 4.112406e-32, 
    4.182375e-32, 4.151923e-32, 4.23172e-32, 4.212462e-32, 4.236437e-32, 
    4.224101e-32, 4.245341e-32, 4.226183e-32, 4.25945e-32, 4.266742e-32, 
    4.261759e-32, 4.280904e-32, 4.225146e-32, 4.246444e-32, 4.092015e-32, 
    4.092889e-32, 4.096958e-32, 4.079099e-32, 4.078005e-32, 4.061679e-32, 
    4.076198e-32, 4.082398e-32, 4.098148e-32, 4.107497e-32, 4.116397e-32, 
    4.13625e-32, 4.158903e-32, 4.190729e-32, 4.213704e-32, 4.229172e-32, 
    4.219675e-32, 4.228053e-32, 4.218691e-32, 4.214306e-32, 4.264013e-32, 
    4.235856e-32, 4.278146e-32, 4.275795e-32, 4.256629e-32, 4.27606e-32, 
    4.093503e-32, 4.088474e-32, 4.071073e-32, 4.084686e-32, 4.059903e-32, 
    4.073768e-32, 4.081762e-32, 4.112689e-32, 4.119494e-32, 4.125831e-32, 
    4.138656e-32, 4.155252e-32, 4.184499e-32, 4.21007e-32, 4.233623e-32, 
    4.23186e-32, 4.232481e-32, 4.237863e-32, 4.224652e-32, 4.24005e-32, 
    4.242662e-32, 4.235846e-32, 4.275481e-32, 4.264127e-32, 4.275745e-32, 
    4.268348e-32, 4.090106e-32, 4.09857e-32, 4.093996e-32, 4.102604e-32, 
    4.096543e-32, 4.123567e-32, 4.131803e-32, 4.171113e-32, 4.154928e-32, 
    4.180693e-32, 4.157535e-32, 4.161634e-32, 4.181562e-32, 4.15878e-32, 
    4.208669e-32, 4.174816e-32, 4.238072e-32, 4.203891e-32, 4.240259e-32, 
    4.233519e-32, 4.244677e-32, 4.254697e-32, 4.267316e-32, 4.290964e-32, 
    4.285365e-32, 4.305592e-32, 4.111208e-32, 4.122239e-32, 4.121256e-32, 
    4.132954e-32, 4.141771e-32, 4.160918e-32, 4.191791e-32, 4.180156e-32, 
    4.201523e-32, 4.205827e-32, 4.173366e-32, 4.193284e-32, 4.129673e-32, 
    4.139909e-32, 4.133803e-32, 4.112084e-32, 4.182851e-32, 4.14618e-32, 
    4.214087e-32, 4.194067e-32, 4.253269e-32, 4.223475e-32, 4.282289e-32, 
    4.308526e-32, 4.334133e-32, 4.36443e-32, 4.128264e-32, 4.120751e-32, 
    4.134367e-32, 4.153578e-32, 4.171435e-32, 4.195288e-32, 4.197729e-32, 
    4.202215e-32, 4.21384e-32, 4.223639e-32, 4.203646e-32, 4.226098e-32, 
    4.142309e-32, 4.186041e-32, 4.117927e-32, 4.138154e-32, 4.152439e-32, 
    4.146156e-32, 4.178825e-32, 4.186559e-32, 4.21811e-32, 4.201769e-32, 
    4.302049e-32, 4.256832e-32, 4.387941e-32, 4.349871e-32, 4.118134e-32, 
    4.128232e-32, 4.164551e-32, 4.147237e-32, 4.196879e-32, 4.209176e-32, 
    4.219184e-32, 4.232098e-32, 4.23351e-32, 4.241314e-32, 4.228542e-32, 
    4.240804e-32, 4.195339e-32, 4.215484e-32, 4.160373e-32, 4.17374e-32, 
    4.167582e-32, 4.160845e-32, 4.181668e-32, 4.203963e-32, 4.204422e-32, 
    4.211595e-32, 4.231965e-32, 4.19708e-32, 4.308055e-32, 4.238517e-32, 
    4.139579e-32, 4.159709e-32, 4.162568e-32, 4.154761e-32, 4.207943e-32, 
    4.188612e-32, 4.24112e-32, 4.226668e-32, 4.250397e-32, 4.238568e-32, 
    4.236831e-32, 4.221844e-32, 4.212653e-32, 4.189501e-32, 4.170733e-32, 
    4.15589e-32, 4.159336e-32, 4.175654e-32, 4.205325e-32, 4.233647e-32, 
    4.227347e-32, 4.248586e-32, 4.193264e-32, 4.216211e-32, 4.207336e-32, 
    4.230543e-32, 4.179851e-32, 4.223012e-32, 4.168883e-32, 4.173602e-32, 
    4.188229e-32, 4.217784e-32, 4.224317e-32, 4.231393e-32, 4.227e-32, 
    4.206077e-32, 4.202649e-32, 4.187868e-32, 4.183804e-32, 4.172573e-32, 
    4.163302e-32, 4.171777e-32, 4.180695e-32, 4.206079e-32, 4.229074e-32, 
    4.254842e-32, 4.26116e-32, 4.291799e-32, 4.266817e-32, 4.308456e-32, 
    4.272955e-32, 4.33567e-32, 4.225496e-32, 4.271899e-32, 4.188889e-32, 
    4.197659e-32, 4.21358e-32, 4.25074e-32, 4.230431e-32, 4.254181e-32, 
    4.202514e-32, 4.176227e-32, 4.169425e-32, 4.156795e-32, 4.169714e-32, 
    4.168661e-32, 4.181052e-32, 4.177066e-32, 4.206923e-32, 4.190863e-32, 
    4.236793e-32, 4.253988e-32, 4.303475e-32, 4.335516e-32, 4.368632e-32, 
    4.383589e-32, 4.388183e-32, 4.390106e-32,
  5.366649e-38, 5.41176e-38, 5.402953e-38, 5.439585e-38, 5.419224e-38, 
    5.443264e-38, 5.375752e-38, 5.413568e-38, 5.389389e-38, 5.37068e-38, 
    5.512514e-38, 5.441223e-38, 5.589091e-38, 5.541893e-38, 5.663037e-38, 
    5.581729e-38, 5.679819e-38, 5.660633e-38, 5.718716e-38, 5.701981e-38, 
    5.777319e-38, 5.726458e-38, 5.817414e-38, 5.765008e-38, 5.773114e-38, 
    5.724797e-38, 5.455261e-38, 5.503409e-38, 5.452471e-38, 5.4592e-38, 
    5.456175e-38, 5.419651e-38, 5.401359e-38, 5.363203e-38, 5.370104e-38, 
    5.398132e-38, 5.462229e-38, 5.440365e-38, 5.496089e-38, 5.49479e-38, 
    5.559227e-38, 5.530071e-38, 5.64074e-38, 5.608453e-38, 5.702678e-38, 
    5.678654e-38, 5.701551e-38, 5.694593e-38, 5.701641e-38, 5.666475e-38, 
    5.6815e-38, 5.650829e-38, 5.535523e-38, 5.568735e-38, 5.470733e-38, 
    5.414479e-38, 5.377408e-38, 5.351285e-38, 5.35497e-38, 5.362006e-38, 
    5.398297e-38, 5.43264e-38, 5.458978e-38, 5.476678e-38, 5.494603e-38, 
    5.549891e-38, 5.579354e-38, 5.647306e-38, 5.634844e-38, 5.65596e-38, 
    5.676269e-38, 5.710809e-38, 5.705104e-38, 5.720385e-38, 5.655387e-38, 
    5.69845e-38, 5.627764e-38, 5.646914e-38, 5.499614e-38, 5.44625e-38, 
    5.424052e-38, 5.404648e-38, 5.357806e-38, 5.390111e-38, 5.377353e-38, 
    5.407744e-38, 5.427161e-38, 5.417545e-38, 5.477163e-38, 5.453903e-38, 
    5.581106e-38, 5.525487e-38, 5.67388e-38, 5.637398e-38, 5.682742e-38, 
    5.659475e-38, 5.699483e-38, 5.66343e-38, 5.726078e-38, 5.739846e-38, 
    5.730435e-38, 5.766658e-38, 5.661458e-38, 5.701558e-38, 5.417279e-38, 
    5.418846e-38, 5.426147e-38, 5.394138e-38, 5.392182e-38, 5.363018e-38, 
    5.388953e-38, 5.400044e-38, 5.428283e-38, 5.445075e-38, 5.461085e-38, 
    5.496976e-38, 5.53821e-38, 5.596422e-38, 5.639752e-38, 5.6691e-38, 
    5.651076e-38, 5.66698e-38, 5.649207e-38, 5.640896e-38, 5.734688e-38, 
    5.681645e-38, 5.761432e-38, 5.75698e-38, 5.720752e-38, 5.757482e-38, 
    5.419946e-38, 5.410934e-38, 5.379791e-38, 5.404146e-38, 5.359851e-38, 
    5.384606e-38, 5.398901e-38, 5.454405e-38, 5.466664e-38, 5.478082e-38, 
    5.50135e-38, 5.53156e-38, 5.585003e-38, 5.632864e-38, 5.677458e-38, 
    5.674147e-38, 5.675313e-38, 5.685419e-38, 5.660519e-38, 5.689532e-38, 
    5.69444e-38, 5.68163e-38, 5.756385e-38, 5.734912e-38, 5.756886e-38, 
    5.74289e-38, 5.413859e-38, 5.429039e-38, 5.420832e-38, 5.436281e-38, 
    5.425398e-38, 5.473993e-38, 5.488887e-38, 5.560501e-38, 5.530968e-38, 
    5.578032e-38, 5.535723e-38, 5.543198e-38, 5.579606e-38, 5.537995e-38, 
    5.630203e-38, 5.567269e-38, 5.685812e-38, 5.621154e-38, 5.689926e-38, 
    5.677263e-38, 5.698239e-38, 5.71711e-38, 5.740938e-38, 5.785512e-38, 
    5.775035e-38, 5.812952e-38, 5.451749e-38, 5.471604e-38, 5.469839e-38, 
    5.490989e-38, 5.50701e-38, 5.541896e-38, 5.598375e-38, 5.577057e-38, 
    5.6167e-38, 5.624837e-38, 5.564635e-38, 5.60113e-38, 5.485027e-38, 
    5.503615e-38, 5.492529e-38, 5.45332e-38, 5.581981e-38, 5.515025e-38, 
    5.640476e-38, 5.602614e-38, 5.714417e-38, 5.658273e-38, 5.769282e-38, 
    5.818447e-38, 5.866195e-38, 5.923491e-38, 5.482473e-38, 5.46893e-38, 
    5.493557e-38, 5.5285e-38, 5.5611e-38, 5.604918e-38, 5.60953e-38, 
    5.618006e-38, 5.640012e-38, 5.658598e-38, 5.620703e-38, 5.663266e-38, 
    5.507964e-38, 5.587828e-38, 5.463839e-38, 5.500423e-38, 5.526427e-38, 
    5.514989e-38, 5.574623e-38, 5.588786e-38, 5.648097e-38, 5.617167e-38, 
    5.80628e-38, 5.721126e-38, 5.969034e-38, 5.895584e-38, 5.464216e-38, 
    5.482418e-38, 5.54852e-38, 5.516957e-38, 5.607924e-38, 5.631174e-38, 
    5.650144e-38, 5.674588e-38, 5.677244e-38, 5.691906e-38, 5.667911e-38, 
    5.69095e-38, 5.605014e-38, 5.643125e-38, 5.540903e-38, 5.565314e-38, 
    5.554064e-38, 5.541764e-38, 5.579826e-38, 5.621302e-38, 5.62218e-38, 
    5.635751e-38, 5.674296e-38, 5.608305e-38, 5.817534e-38, 5.686612e-38, 
    5.50303e-38, 5.539676e-38, 5.544904e-38, 5.530667e-38, 5.628839e-38, 
    5.592547e-38, 5.691545e-38, 5.664351e-38, 5.709009e-38, 5.686747e-38, 
    5.683481e-38, 5.655189e-38, 5.637759e-38, 5.594173e-38, 5.559816e-38, 
    5.532727e-38, 5.539011e-38, 5.568813e-38, 5.62388e-38, 5.677496e-38, 
    5.665631e-38, 5.705597e-38, 5.601099e-38, 5.644498e-38, 5.627686e-38, 
    5.671672e-38, 5.576496e-38, 5.657368e-38, 5.55644e-38, 5.565067e-38, 
    5.591845e-38, 5.647472e-38, 5.659884e-38, 5.673264e-38, 5.66498e-38, 
    5.625305e-38, 5.618825e-38, 5.591186e-38, 5.583734e-38, 5.563186e-38, 
    5.546248e-38, 5.561727e-38, 5.578039e-38, 5.625312e-38, 5.66891e-38, 
    5.717383e-38, 5.729308e-38, 5.787057e-38, 5.739972e-38, 5.818287e-38, 
    5.751551e-38, 5.869029e-38, 5.6621e-38, 5.749578e-38, 5.593059e-38, 
    5.6094e-38, 5.639505e-38, 5.709639e-38, 5.671462e-38, 5.716127e-38, 
    5.61857e-38, 5.569856e-38, 5.55743e-38, 5.534373e-38, 5.557958e-38, 
    5.556035e-38, 5.578699e-38, 5.571404e-38, 5.626911e-38, 5.596677e-38, 
    5.683405e-38, 5.715767e-38, 5.808973e-38, 5.868764e-38, 5.931615e-38, 
    5.960584e-38, 5.969511e-38, 5.973248e-38,
  2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 
    2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 3.082857e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  4.994591e-06, 4.730369e-06, 4.781403e-06, 4.570714e-06, 4.687216e-06, 
    4.549785e-06, 4.940677e-06, 4.719986e-06, 4.860528e-06, 4.970608e-06, 
    4.170714e-06, 4.561377e-06, 3.776003e-06, 4.014818e-06, 3.426535e-06, 
    3.812812e-06, 3.350878e-06, 3.437374e-06, 3.18011e-06, 3.252823e-06, 
    2.934725e-06, 3.146826e-06, 2.776593e-06, 2.984648e-06, 2.951576e-06, 
    3.153961e-06, 4.481774e-06, 4.218712e-06, 4.497538e-06, 4.459654e-06, 
    4.476628e-06, 4.68482e-06, 4.790854e-06, 5.014907e-06, 4.974013e-06, 
    4.809529e-06, 4.442652e-06, 4.566145e-06, 4.256963e-06, 4.263863e-06, 
    3.926113e-06, 4.075866e-06, 3.529176e-06, 3.68122e-06, 3.249771e-06, 
    3.355946e-06, 3.25473e-06, 3.285258e-06, 3.254333e-06, 3.410705e-06, 
    3.343283e-06, 3.482417e-06, 4.047667e-06, 3.87796e-06, 4.394967e-06, 
    4.7149e-06, 4.930949e-06, 5.085899e-06, 5.063918e-06, 5.022094e-06, 
    4.808572e-06, 4.610202e-06, 4.460776e-06, 4.361724e-06, 4.264856e-06, 
    3.974053e-06, 3.824635e-06, 3.498798e-06, 3.556631e-06, 3.458878e-06, 
    3.366596e-06, 3.214374e-06, 3.239189e-06, 3.172973e-06, 3.461412e-06, 
    3.268385e-06, 3.58977e-06, 3.500504e-06, 4.238834e-06, 4.532714e-06, 
    4.659707e-06, 4.771588e-06, 5.047038e-06, 4.856371e-06, 4.931302e-06, 
    4.753529e-06, 4.641583e-06, 4.696843e-06, 4.359026e-06, 4.48941e-06, 
    3.815851e-06, 4.099778e-06, 3.377299e-06, 3.544723e-06, 3.337721e-06, 
    3.442627e-06, 3.263829e-06, 3.424544e-06, 3.148491e-06, 3.089915e-06, 
    3.129887e-06, 2.977739e-06, 3.433564e-06, 3.254745e-06, 4.698403e-06, 
    4.689378e-06, 4.647375e-06, 4.832837e-06, 4.844239e-06, 5.016039e-06, 
    4.863074e-06, 4.798349e-06, 4.635104e-06, 4.539389e-06, 4.448975e-06, 
    4.252315e-06, 4.033869e-06, 3.739528e-06, 3.533761e-06, 3.39873e-06, 
    3.481234e-06, 3.408348e-06, 3.489879e-06, 3.528386e-06, 3.111807e-06, 
    3.342668e-06, 2.999379e-06, 3.017875e-06, 3.171413e-06, 3.015787e-06, 
    4.68304e-06, 4.735034e-06, 4.916895e-06, 4.774406e-06, 5.034842e-06, 
    4.888617e-06, 4.805091e-06, 4.486712e-06, 4.417639e-06, 4.353964e-06, 
    4.22909e-06, 4.06815e-06, 3.796272e-06, 3.565964e-06, 3.361256e-06, 
    3.376063e-06, 3.370848e-06, 3.32584e-06, 3.437868e-06, 3.307614e-06, 
    3.286002e-06, 3.342676e-06, 3.020357e-06, 3.110763e-06, 3.018269e-06, 
    3.076951e-06, 4.718109e-06, 4.630806e-06, 4.677924e-06, 4.589453e-06, 
    4.651743e-06, 4.376869e-06, 4.295534e-06, 3.919777e-06, 4.071253e-06, 
    3.831187e-06, 4.046597e-06, 4.008105e-06, 3.823527e-06, 4.034829e-06, 
    3.578533e-06, 3.885538e-06, 3.324096e-06, 3.621246e-06, 3.305872e-06, 
    3.36213e-06, 3.269215e-06, 3.187087e-06, 3.085219e-06, 2.901804e-06, 
    2.943738e-06, 2.793809e-06, 4.501573e-06, 4.390123e-06, 4.399864e-06, 
    4.284123e-06, 4.199222e-06, 4.014734e-06, 3.729807e-06, 3.835955e-06, 
    3.642004e-06, 3.603594e-06, 3.898582e-06, 3.716347e-06, 4.316029e-06, 
    4.217299e-06, 4.275961e-06, 4.492769e-06, 3.811431e-06, 4.157195e-06, 
    3.530408e-06, 3.70916e-06, 3.198738e-06, 3.448287e-06, 2.966967e-06, 
    2.772731e-06, 2.596611e-06, 2.399739e-06, 4.329652e-06, 4.404938e-06, 
    4.27042e-06, 4.084171e-06, 3.916582e-06, 3.698154e-06, 3.676081e-06, 
    3.635853e-06, 3.532506e-06, 3.446657e-06, 3.623203e-06, 3.425283e-06, 
    4.194585e-06, 3.782188e-06, 4.433547e-06, 4.234219e-06, 4.094888e-06, 
    4.157253e-06, 3.848156e-06, 3.777299e-06, 3.495112e-06, 3.639789e-06, 
    2.820017e-06, 3.169914e-06, 2.256406e-06, 2.493052e-06, 4.431353e-06, 
    4.329895e-06, 3.980828e-06, 4.146913e-06, 3.68374e-06, 3.57383e-06, 
    3.485532e-06, 3.374172e-06, 3.362228e-06, 3.29715e-06, 3.404108e-06, 
    3.301332e-06, 3.697695e-06, 3.518066e-06, 4.019817e-06, 3.895208e-06, 
    3.952332e-06, 4.015387e-06, 3.822046e-06, 3.620402e-06, 3.616093e-06, 
    3.552468e-06, 3.375992e-06, 3.681919e-06, 2.776551e-06, 3.321032e-06, 
    4.220182e-06, 4.026373e-06, 3.999291e-06, 4.072733e-06, 3.584786e-06, 
    3.758654e-06, 3.298722e-06, 3.420337e-06, 3.222162e-06, 3.319938e-06, 
    3.334444e-06, 3.462306e-06, 3.543037e-06, 3.750615e-06, 3.923117e-06, 
    4.062043e-06, 4.029571e-06, 3.877542e-06, 3.608207e-06, 3.361168e-06, 
    3.414606e-06, 3.237022e-06, 3.716395e-06, 3.511765e-06, 3.590274e-06, 
    3.3872e-06, 3.838804e-06, 3.452804e-06, 3.94021e-06, 3.896402e-06, 
    3.762139e-06, 3.498103e-06, 3.440762e-06, 3.380105e-06, 3.417464e-06, 
    3.601467e-06, 3.631997e-06, 3.765367e-06, 3.80257e-06, 3.90592e-06, 
    3.992336e-06, 3.913365e-06, 3.831112e-06, 3.601367e-06, 3.399668e-06, 
    3.185933e-06, 3.134645e-06, 2.895892e-06, 3.089564e-06, 2.773674e-06, 
    3.041174e-06, 2.586839e-06, 3.430918e-06, 3.049147e-06, 3.756058e-06, 
    3.67669e-06, 3.535038e-06, 3.219627e-06, 3.388142e-06, 3.191456e-06, 
    3.633191e-06, 3.872363e-06, 3.935186e-06, 4.053555e-06, 3.932496e-06, 
    3.942287e-06, 3.827683e-06, 3.864362e-06, 3.593842e-06, 3.738132e-06, 
    3.334822e-06, 3.192975e-06, 2.809334e-06, 2.587566e-06, 2.373024e-06, 
    2.282111e-06, 2.254907e-06, 2.243604e-06,
  7.830288e-06, 7.669716e-06, 7.70068e-06, 7.573055e-06, 7.643577e-06, 
    7.560408e-06, 7.79748e-06, 7.663407e-06, 7.748738e-06, 7.815705e-06, 
    7.332205e-06, 7.567415e-06, 6.816401e-06, 6.926776e-06, 6.656883e-06, 
    6.833329e-06, 6.622676e-06, 6.661816e-06, 6.545916e-06, 6.578533e-06, 
    6.436691e-06, 6.531025e-06, 6.367121e-06, 6.45881e-06, 6.444155e-06, 
    6.534213e-06, 7.519364e-06, 7.360983e-06, 7.528875e-06, 7.506006e-06, 
    7.516258e-06, 7.642112e-06, 7.706379e-06, 7.842691e-06, 7.817779e-06, 
    7.717741e-06, 7.495748e-06, 7.57032e-06, 7.384053e-06, 7.388197e-06, 
    6.885664e-06, 6.955164e-06, 6.703507e-06, 6.772931e-06, 6.577162e-06, 
    6.624983e-06, 6.579386e-06, 6.593119e-06, 6.579208e-06, 6.649735e-06, 
    6.619262e-06, 6.682254e-06, 6.942041e-06, 6.8634e-06, 7.467025e-06, 
    7.660287e-06, 7.791553e-06, 7.88597e-06, 7.872562e-06, 7.847054e-06, 
    7.717159e-06, 7.596959e-06, 7.506708e-06, 7.447029e-06, 7.388794e-06, 
    6.90782e-06, 6.838787e-06, 6.68968e-06, 6.716013e-06, 6.671557e-06, 
    6.629793e-06, 6.561266e-06, 6.572406e-06, 6.542713e-06, 6.672721e-06, 
    6.585516e-06, 6.731128e-06, 6.690471e-06, 7.37305e-06, 7.55012e-06, 
    7.62686e-06, 7.694718e-06, 7.862265e-06, 7.746196e-06, 7.791762e-06, 
    7.683782e-06, 7.615947e-06, 7.64942e-06, 7.445405e-06, 7.523977e-06, 
    6.834741e-06, 6.966285e-06, 6.634628e-06, 6.710587e-06, 6.616758e-06, 
    6.664205e-06, 6.583471e-06, 6.65601e-06, 6.531764e-06, 6.505606e-06, 
    6.523446e-06, 6.455761e-06, 6.660095e-06, 6.579386e-06, 7.650359e-06, 
    7.644889e-06, 7.619458e-06, 7.731895e-06, 7.738828e-06, 7.843374e-06, 
    7.750285e-06, 7.710961e-06, 7.612035e-06, 7.55415e-06, 7.499582e-06, 
    7.381251e-06, 6.935615e-06, 6.799653e-06, 6.705596e-06, 6.644324e-06, 
    6.681723e-06, 6.648676e-06, 6.685646e-06, 6.703157e-06, 6.515369e-06, 
    6.61898e-06, 6.465355e-06, 6.473566e-06, 6.542011e-06, 6.472639e-06, 
    7.64105e-06, 7.672569e-06, 7.783007e-06, 7.696448e-06, 7.854837e-06, 
    7.765803e-06, 7.715037e-06, 7.522322e-06, 7.480701e-06, 7.442347e-06, 
    7.367317e-06, 6.951573e-06, 6.825741e-06, 6.720256e-06, 6.627385e-06, 
    6.634075e-06, 6.631718e-06, 6.611397e-06, 6.662044e-06, 6.603183e-06, 
    6.593443e-06, 6.618993e-06, 6.474668e-06, 6.514916e-06, 6.473741e-06, 
    6.499843e-06, 7.662309e-06, 7.609426e-06, 7.637955e-06, 7.584402e-06, 
    7.622087e-06, 7.456107e-06, 7.407175e-06, 6.882711e-06, 6.953012e-06, 
    6.841818e-06, 6.941549e-06, 6.92366e-06, 6.838253e-06, 6.936084e-06, 
    6.725971e-06, 6.866876e-06, 6.61061e-06, 6.745449e-06, 6.602398e-06, 
    6.627779e-06, 6.585903e-06, 6.549034e-06, 6.503524e-06, 6.422171e-06, 
    6.440702e-06, 6.374675e-06, 7.53132e-06, 7.464103e-06, 7.469995e-06, 
    7.400361e-06, 7.349391e-06, 6.926748e-06, 6.7952e-06, 6.844034e-06, 
    6.754985e-06, 6.73743e-06, 6.872945e-06, 6.789017e-06, 7.419522e-06, 
    7.360202e-06, 7.395449e-06, 7.52599e-06, 6.832711e-06, 7.324174e-06, 
    6.704067e-06, 6.785731e-06, 6.554254e-06, 6.666749e-06, 6.450982e-06, 
    6.365412e-06, 6.288766e-06, 6.204174e-06, 7.427725e-06, 7.473052e-06, 
    7.392135e-06, 6.959008e-06, 6.881256e-06, 6.780682e-06, 6.770578e-06, 
    6.752166e-06, 6.705031e-06, 6.66603e-06, 6.746369e-06, 6.656345e-06, 
    7.346528e-06, 6.81926e-06, 7.490274e-06, 7.37035e-06, 6.964007e-06, 
    7.324236e-06, 6.849665e-06, 6.817029e-06, 6.688009e-06, 6.753972e-06, 
    6.386143e-06, 6.541324e-06, 6.143512e-06, 6.244099e-06, 7.488968e-06, 
    7.427881e-06, 6.910998e-06, 7.318046e-06, 6.774086e-06, 6.723848e-06, 
    6.683675e-06, 6.633209e-06, 6.627821e-06, 6.598466e-06, 6.646758e-06, 
    6.600355e-06, 6.780472e-06, 6.698456e-06, 6.929113e-06, 6.871376e-06, 
    6.897813e-06, 6.927055e-06, 6.837627e-06, 6.745086e-06, 6.743141e-06, 
    6.714106e-06, 6.633955e-06, 6.773252e-06, 6.367043e-06, 6.609158e-06, 
    7.361976e-06, 6.932122e-06, 6.919575e-06, 6.953712e-06, 6.728845e-06, 
    6.80845e-06, 6.599177e-06, 6.654104e-06, 6.564765e-06, 6.608738e-06, 
    6.615278e-06, 6.673129e-06, 6.709819e-06, 6.804753e-06, 6.884277e-06, 
    6.948741e-06, 6.933643e-06, 6.86321e-06, 6.73952e-06, 6.627333e-06, 
    6.651493e-06, 6.571436e-06, 6.789053e-06, 6.69558e-06, 6.731338e-06, 
    6.639105e-06, 6.845342e-06, 6.668744e-06, 6.892201e-06, 6.871936e-06, 
    6.810053e-06, 6.689354e-06, 6.663358e-06, 6.63589e-06, 6.652804e-06, 
    6.736447e-06, 6.750401e-06, 6.811542e-06, 6.828645e-06, 6.876338e-06, 
    6.916357e-06, 6.879774e-06, 6.841789e-06, 6.736411e-06, 6.644736e-06, 
    6.548514e-06, 6.525579e-06, 6.419528e-06, 6.505422e-06, 6.365779e-06, 
    6.483829e-06, 6.284486e-06, 6.658853e-06, 6.487418e-06, 6.807266e-06, 
    6.770858e-06, 6.706157e-06, 6.563597e-06, 6.639531e-06, 6.550973e-06, 
    6.750949e-06, 6.860806e-06, 6.889873e-06, 6.944786e-06, 6.888628e-06, 
    6.893161e-06, 6.840226e-06, 6.857142e-06, 6.732977e-06, 6.799031e-06, 
    6.615443e-06, 6.55166e-06, 6.381478e-06, 6.284832e-06, 6.192828e-06, 
    6.154339e-06, 6.14289e-06, 6.13814e-06,
  9.692865e-06, 9.704537e-06, 9.702479e-06, 9.71033e-06, 9.7062e-06, 
    9.711014e-06, 9.695445e-06, 9.704944e-06, 9.699098e-06, 9.694025e-06, 
    9.720122e-06, 9.710638e-06, 1.004604e-05, 1.008932e-05, 9.978725e-06, 
    1.005284e-05, 9.963439e-06, 9.980909e-06, 9.927876e-06, 9.943213e-06, 
    9.873816e-06, 9.920758e-06, 9.836911e-06, 9.885127e-06, 9.877655e-06, 
    9.922287e-06, 9.713113e-06, 9.719332e-06, 9.712644e-06, 9.713754e-06, 
    9.713264e-06, 9.706291e-06, 9.702087e-06, 9.691866e-06, 9.693861e-06, 
    9.701303e-06, 9.714233e-06, 9.710481e-06, 9.718628e-06, 9.718492e-06, 
    1.007349e-05, 1.010007e-05, 9.999055e-06, 1.002831e-05, 9.942575e-06, 
    9.964485e-06, 9.943608e-06, 9.949962e-06, 9.943526e-06, 9.975563e-06, 
    9.961899e-06, 9.989862e-06, 1.009512e-05, 1.006477e-05, 9.715508e-06, 
    9.705142e-06, 9.695901e-06, 9.68827e-06, 9.689401e-06, 9.691509e-06, 
    9.701344e-06, 9.708991e-06, 9.713723e-06, 9.716338e-06, 9.718472e-06, 
    1.008205e-05, 1.005502e-05, 9.993084e-06, 1.000441e-05, 9.985187e-06, 
    9.966652e-06, 9.935135e-06, 9.940357e-06, 9.926348e-06, 9.985701e-06, 
    9.94645e-06, 1.001083e-05, 9.99343e-06, 9.718969e-06, 9.71156e-06, 
    9.707224e-06, 9.702882e-06, 9.690259e-06, 9.699282e-06, 9.695885e-06, 
    9.703615e-06, 9.707882e-06, 9.705836e-06, 9.716404e-06, 9.712888e-06, 
    1.005341e-05, 1.010424e-05, 9.968823e-06, 1.000209e-05, 9.960766e-06, 
    9.981963e-06, 9.945503e-06, 9.978346e-06, 9.921112e-06, 9.908429e-06, 
    9.917104e-06, 9.883584e-06, 9.98015e-06, 9.943607e-06, 9.705776e-06, 
    9.706119e-06, 9.707673e-06, 9.700308e-06, 9.699813e-06, 9.691809e-06, 
    9.698985e-06, 9.701774e-06, 9.708114e-06, 9.711348e-06, 9.714056e-06, 
    9.718717e-06, 1.009268e-05, 1.003926e-05, 9.999952e-06, 9.973158e-06, 
    9.989632e-06, 9.975094e-06, 9.991339e-06, 9.998907e-06, 9.913188e-06, 
    9.96177e-06, 9.888439e-06, 9.892567e-06, 9.926013e-06, 9.892103e-06, 
    9.706358e-06, 9.704352e-06, 9.696553e-06, 9.702766e-06, 9.690873e-06, 
    9.697844e-06, 9.701491e-06, 9.712968e-06, 9.714914e-06, 9.716525e-06, 
    9.719151e-06, 1.009872e-05, 1.00498e-05, 1.000622e-05, 9.965569e-06, 
    9.968576e-06, 9.967518e-06, 9.958329e-06, 9.981009e-06, 9.954581e-06, 
    9.950109e-06, 9.961778e-06, 9.89312e-06, 9.912973e-06, 9.892655e-06, 
    9.905607e-06, 9.705017e-06, 9.708267e-06, 9.706549e-06, 9.709703e-06, 
    9.707514e-06, 9.715965e-06, 9.717842e-06, 1.007233e-05, 1.009926e-05, 
    1.005623e-05, 1.009493e-05, 1.008813e-05, 1.00548e-05, 1.009286e-05, 
    1.000864e-05, 1.006613e-05, 9.957971e-06, 1.001686e-05, 9.954222e-06, 
    9.965746e-06, 9.946632e-06, 9.929355e-06, 9.907412e-06, 9.866291e-06, 
    9.875887e-06, 9.841026e-06, 9.712522e-06, 9.715632e-06, 9.715382e-06, 
    9.718082e-06, 9.71967e-06, 1.008931e-05, 1.003745e-05, 1.005712e-05, 
    1.002086e-05, 1.001349e-05, 1.006852e-05, 1.003492e-05, 9.717398e-06, 
    9.71936e-06, 9.718249e-06, 9.712788e-06, 1.00526e-05, 9.720326e-06, 
    9.999296e-06, 1.003357e-05, 9.931827e-06, 9.983076e-06, 9.88115e-06, 
    9.835971e-06, 9.792565e-06, 9.740675e-06, 9.717092e-06, 9.71525e-06, 
    9.718362e-06, 1.010151e-05, 1.007177e-05, 1.00315e-05, 1.002733e-05, 
    1.001968e-05, 9.999712e-06, 9.982766e-06, 1.001725e-05, 9.978495e-06, 
    9.719744e-06, 1.00472e-05, 9.714484e-06, 9.719056e-06, 1.010338e-05, 
    9.720326e-06, 1.005935e-05, 1.00463e-05, 9.99236e-06, 1.002043e-05, 
    9.84721e-06, 9.925681e-06, 9.700333e-06, 9.765738e-06, 9.714544e-06, 
    9.717087e-06, 1.008328e-05, 9.720476e-06, 1.002878e-05, 1.000775e-05, 
    9.990482e-06, 9.968185e-06, 9.965765e-06, 9.95242e-06, 9.974242e-06, 
    9.953287e-06, 1.003141e-05, 9.996882e-06, 1.009021e-05, 1.006791e-05, 
    1.00782e-05, 1.008943e-05, 1.005456e-05, 1.001671e-05, 1.00159e-05, 
    1.000359e-05, 9.968501e-06, 1.002844e-05, 9.83685e-06, 9.957293e-06, 
    9.71931e-06, 1.009135e-05, 1.008657e-05, 1.009952e-05, 1.000987e-05, 
    1.004283e-05, 9.952746e-06, 9.977502e-06, 9.93678e-06, 9.957119e-06, 
    9.960094e-06, 9.985879e-06, 1.000176e-05, 1.004133e-05, 1.007295e-05, 
    1.009765e-05, 1.009194e-05, 1.00647e-05, 1.001437e-05, 9.965543e-06, 
    9.976341e-06, 9.939904e-06, 1.003494e-05, 9.995639e-06, 1.001092e-05, 
    9.970827e-06, 1.005763e-05, 9.98394e-06, 1.007603e-05, 1.006813e-05, 
    1.004348e-05, 9.99294e-06, 9.98159e-06, 9.969387e-06, 9.976927e-06, 
    1.001308e-05, 1.001894e-05, 1.004409e-05, 1.005097e-05, 1.006985e-05, 
    1.008534e-05, 1.007119e-05, 1.005622e-05, 1.001306e-05, 9.973338e-06, 
    9.929107e-06, 9.918136e-06, 9.864901e-06, 9.908332e-06, 9.836158e-06, 
    9.897666e-06, 9.79003e-06, 9.979593e-06, 9.89946e-06, 1.004236e-05, 
    1.002745e-05, 1.000019e-05, 9.936224e-06, 9.971018e-06, 9.93027e-06, 
    1.001917e-05, 1.006375e-05, 1.007512e-05, 1.009616e-05, 1.007464e-05, 
    1.00764e-05, 1.00556e-05, 1.006231e-05, 1.001161e-05, 1.003901e-05, 
    9.960167e-06, 9.930596e-06, 9.844705e-06, 9.790244e-06, 9.733356e-06, 
    9.707757e-06, 9.699907e-06, 9.696616e-06,
  4.369429e-06, 4.283271e-06, 4.300009e-06, 4.230615e-06, 4.269097e-06, 
    4.223677e-06, 4.351951e-06, 4.279851e-06, 4.325866e-06, 4.361671e-06, 
    4.096314e-06, 4.227523e-06, 3.960923e-06, 4.044187e-06, 3.835547e-06, 
    3.973858e-06, 3.807759e-06, 3.839535e-06, 3.744059e-06, 3.771368e-06, 
    3.649712e-06, 3.731467e-06, 3.586968e-06, 3.669209e-06, 3.656316e-06, 
    3.734168e-06, 4.201086e-06, 4.112618e-06, 4.206333e-06, 4.193702e-06, 
    4.199371e-06, 4.268299e-06, 4.303075e-06, 4.376026e-06, 4.362775e-06, 
    4.309202e-06, 4.188024e-06, 4.229121e-06, 4.125657e-06, 4.12799e-06, 
    4.013475e-06, 4.065201e-06, 3.872888e-06, 3.927404e-06, 3.770228e-06, 
    3.809651e-06, 3.772076e-06, 3.783464e-06, 3.771928e-06, 3.829777e-06, 
    3.804972e-06, 3.855947e-06, 4.055505e-06, 3.996696e-06, 4.172084e-06, 
    4.278153e-06, 4.348785e-06, 4.398968e-06, 4.39187e-06, 4.378341e-06, 
    4.308888e-06, 4.243701e-06, 4.194095e-06, 4.160951e-06, 4.128326e-06, 
    4.030053e-06, 3.97802e-06, 3.861875e-06, 3.882803e-06, 3.847368e-06, 
    3.813577e-06, 3.756954e-06, 3.766264e-06, 3.741353e-06, 3.848308e-06, 
    3.777163e-06, 3.89473e-06, 3.862513e-06, 4.119431e-06, 4.21803e-06, 
    4.259996e-06, 4.296789e-06, 4.386413e-06, 4.3245e-06, 4.348895e-06, 
    4.290885e-06, 4.254063e-06, 4.272271e-06, 4.160045e-06, 4.203633e-06, 
    3.974939e-06, 4.073387e-06, 3.817516e-06, 3.878507e-06, 3.802923e-06, 
    3.841461e-06, 3.775467e-06, 3.834853e-06, 3.732092e-06, 3.70978e-06, 
    3.725024e-06, 3.66654e-06, 3.838149e-06, 3.772073e-06, 4.272781e-06, 
    4.26981e-06, 4.255977e-06, 4.316817e-06, 4.320544e-06, 4.376388e-06, 
    4.326697e-06, 4.305551e-06, 4.251932e-06, 4.220245e-06, 4.190151e-06, 
    4.124076e-06, 4.050743e-06, 3.948061e-06, 3.874548e-06, 3.825396e-06, 
    3.855524e-06, 3.828923e-06, 3.858661e-06, 3.872615e-06, 3.718135e-06, 
    3.804739e-06, 3.674941e-06, 3.682102e-06, 3.74076e-06, 3.681296e-06, 
    4.267725e-06, 4.28482e-06, 4.344219e-06, 4.297727e-06, 4.382474e-06, 
    4.335013e-06, 4.307744e-06, 4.202715e-06, 4.179686e-06, 4.158336e-06, 
    4.116218e-06, 4.062551e-06, 3.968075e-06, 3.886152e-06, 3.811615e-06, 
    3.817068e-06, 3.815148e-06, 3.798524e-06, 3.83972e-06, 3.791769e-06, 
    3.783729e-06, 3.804753e-06, 3.683062e-06, 3.717754e-06, 3.682255e-06, 
    3.704836e-06, 4.279263e-06, 4.250508e-06, 4.266043e-06, 4.236833e-06, 
    4.257407e-06, 4.166004e-06, 4.138646e-06, 4.011249e-06, 4.063612e-06, 
    3.98033e-06, 4.055143e-06, 4.041871e-06, 3.977606e-06, 4.051097e-06, 
    3.890656e-06, 3.999313e-06, 3.797879e-06, 3.905956e-06, 3.791123e-06, 
    3.811936e-06, 3.77749e-06, 3.746683e-06, 3.707997e-06, 3.636809e-06, 
    3.653272e-06, 3.593899e-06, 4.207682e-06, 4.170458e-06, 4.173739e-06, 
    4.134828e-06, 4.106079e-06, 4.04417e-06, 3.944633e-06, 3.982022e-06, 
    3.91343e-06, 3.899681e-06, 4.003907e-06, 3.939858e-06, 4.145573e-06, 
    4.11219e-06, 4.132066e-06, 4.204741e-06, 3.973394e-06, 4.091763e-06, 
    3.873333e-06, 3.937322e-06, 3.751072e-06, 3.843501e-06, 3.662338e-06, 
    3.585389e-06, 3.513305e-06, 3.429437e-06, 4.150166e-06, 4.175439e-06, 
    4.130206e-06, 4.068028e-06, 4.010163e-06, 3.933413e-06, 3.925576e-06, 
    3.911226e-06, 3.874102e-06, 3.842931e-06, 3.906685e-06, 3.835124e-06, 
    4.104442e-06, 3.963118e-06, 4.184993e-06, 4.117921e-06, 4.071711e-06, 
    4.091804e-06, 3.9863e-06, 3.961416e-06, 3.860543e-06, 3.91264e-06, 
    3.604345e-06, 3.740173e-06, 3.36591e-06, 3.46964e-06, 4.184272e-06, 
    4.150255e-06, 4.032438e-06, 4.088283e-06, 3.928301e-06, 3.88899e-06, 
    3.857086e-06, 3.816358e-06, 3.811969e-06, 3.787879e-06, 3.827369e-06, 
    3.78944e-06, 3.93325e-06, 3.868875e-06, 4.045927e-06, 4.002721e-06, 
    4.022591e-06, 4.044399e-06, 3.977148e-06, 3.905679e-06, 3.904163e-06, 
    3.88129e-06, 3.816937e-06, 3.927653e-06, 3.58687e-06, 3.796659e-06, 
    4.113202e-06, 4.048149e-06, 4.038834e-06, 4.064133e-06, 3.892928e-06, 
    3.954832e-06, 3.788467e-06, 3.833314e-06, 3.759885e-06, 3.796341e-06, 
    3.801709e-06, 3.848636e-06, 3.877898e-06, 3.951989e-06, 4.012433e-06, 
    4.060463e-06, 4.049289e-06, 3.996554e-06, 3.901316e-06, 3.811568e-06, 
    3.831196e-06, 3.765456e-06, 3.939891e-06, 3.866582e-06, 3.894887e-06, 
    3.821157e-06, 3.983014e-06, 3.845086e-06, 4.018386e-06, 4.003147e-06, 
    3.956063e-06, 3.861611e-06, 3.840779e-06, 3.81854e-06, 3.832262e-06, 
    3.898905e-06, 3.909845e-06, 3.957208e-06, 3.970296e-06, 4.006465e-06, 
    4.03644e-06, 4.009049e-06, 3.98031e-06, 3.89888e-06, 3.825725e-06, 
    3.746243e-06, 3.726842e-06, 3.634435e-06, 3.709612e-06, 3.585706e-06, 
    3.690978e-06, 3.509154e-06, 3.837131e-06, 3.694101e-06, 3.953925e-06, 
    3.925795e-06, 3.874986e-06, 3.758896e-06, 3.821503e-06, 3.748307e-06, 
    3.910274e-06, 3.994732e-06, 4.016639e-06, 4.057539e-06, 4.015705e-06, 
    4.019105e-06, 3.979128e-06, 3.991969e-06, 3.896181e-06, 3.94759e-06, 
    3.801842e-06, 3.748887e-06, 3.600109e-06, 3.509502e-06, 3.417803e-06, 
    3.377492e-06, 3.365245e-06, 3.360128e-06,
  4.506544e-07, 4.337498e-07, 4.370065e-07, 4.2359e-07, 4.310023e-07, 
    4.222612e-07, 4.47197e-07, 4.330859e-07, 4.420636e-07, 4.491179e-07, 
    3.982628e-07, 4.229975e-07, 3.73526e-07, 3.886024e-07, 3.514235e-07, 
    3.758472e-07, 3.466216e-07, 3.521155e-07, 3.357462e-07, 3.403862e-07, 
    3.199751e-07, 3.336182e-07, 3.097085e-07, 3.232015e-07, 3.210661e-07, 
    3.340741e-07, 4.179493e-07, 4.012929e-07, 4.189485e-07, 4.165451e-07, 
    4.176229e-07, 4.308478e-07, 4.376046e-07, 4.519634e-07, 4.493365e-07, 
    4.388008e-07, 4.15467e-07, 4.233036e-07, 4.037249e-07, 4.041609e-07, 
    3.830044e-07, 3.924579e-07, 3.579314e-07, 3.675466e-07, 3.401917e-07, 
    3.469475e-07, 3.40507e-07, 3.424522e-07, 3.404817e-07, 3.504235e-07, 
    3.46142e-07, 3.54971e-07, 3.906764e-07, 3.799644e-07, 4.124488e-07, 
    4.327566e-07, 4.465721e-07, 4.565307e-07, 4.551149e-07, 4.524229e-07, 
    4.387396e-07, 4.261028e-07, 4.166199e-07, 4.103476e-07, 4.042236e-07, 
    3.860208e-07, 3.765958e-07, 3.560055e-07, 3.5967e-07, 3.534767e-07, 
    3.476242e-07, 3.37933e-07, 3.395165e-07, 3.352883e-07, 3.536403e-07, 
    3.413751e-07, 3.617674e-07, 3.561167e-07, 4.025627e-07, 4.211811e-07, 
    4.292431e-07, 4.363791e-07, 4.540281e-07, 4.417955e-07, 4.46594e-07, 
    4.352297e-07, 4.280982e-07, 4.316168e-07, 4.101769e-07, 4.184342e-07, 
    3.760416e-07, 3.939652e-07, 3.483037e-07, 3.589161e-07, 3.457896e-07, 
    3.524501e-07, 3.410856e-07, 3.513031e-07, 3.337236e-07, 3.299697e-07, 
    3.32532e-07, 3.227589e-07, 3.518749e-07, 3.405065e-07, 4.317154e-07, 
    4.311402e-07, 4.284674e-07, 4.402903e-07, 4.410201e-07, 4.520352e-07, 
    4.422266e-07, 4.380879e-07, 4.276874e-07, 4.216045e-07, 4.158707e-07, 
    4.034295e-07, 3.89803e-07, 3.712257e-07, 3.582221e-07, 3.496653e-07, 
    3.548973e-07, 3.502756e-07, 3.554444e-07, 3.578835e-07, 3.313728e-07, 
    3.461019e-07, 3.241533e-07, 3.253444e-07, 3.35188e-07, 3.252101e-07, 
    4.307367e-07, 4.340507e-07, 4.45672e-07, 4.365618e-07, 4.532446e-07, 
    4.4386e-07, 4.385161e-07, 4.182594e-07, 4.138868e-07, 4.098551e-07, 
    4.019635e-07, 3.919706e-07, 3.748086e-07, 3.602583e-07, 3.472858e-07, 
    3.482264e-07, 3.47895e-07, 3.450337e-07, 3.521476e-07, 3.438745e-07, 
    3.424975e-07, 3.461043e-07, 3.255041e-07, 3.313087e-07, 3.253698e-07, 
    3.29141e-07, 4.329719e-07, 4.27413e-07, 4.304114e-07, 4.24783e-07, 
    4.287432e-07, 4.113005e-07, 4.061555e-07, 3.826003e-07, 3.921655e-07, 
    3.770116e-07, 3.9061e-07, 3.881787e-07, 3.765212e-07, 3.89868e-07, 
    3.610503e-07, 3.804377e-07, 3.449228e-07, 3.637475e-07, 3.437636e-07, 
    3.473413e-07, 3.414309e-07, 3.361906e-07, 3.296709e-07, 3.178495e-07, 
    3.205629e-07, 3.108338e-07, 4.192057e-07, 4.121416e-07, 4.127617e-07, 
    4.054403e-07, 4.000761e-07, 3.885993e-07, 3.706137e-07, 3.773162e-07, 
    3.650691e-07, 3.6264e-07, 3.812692e-07, 3.697623e-07, 4.074549e-07, 
    4.012132e-07, 4.049232e-07, 4.186452e-07, 3.757638e-07, 3.974193e-07, 
    3.580094e-07, 3.693106e-07, 3.369345e-07, 3.528044e-07, 3.220626e-07, 
    3.094524e-07, 2.978794e-07, 2.847059e-07, 4.083177e-07, 4.13083e-07, 
    4.045751e-07, 3.92978e-07, 3.824032e-07, 3.686148e-07, 3.672222e-07, 
    3.646792e-07, 3.58144e-07, 3.527053e-07, 3.638764e-07, 3.513501e-07, 
    3.997718e-07, 3.739194e-07, 4.148923e-07, 4.02281e-07, 3.936564e-07, 
    3.974269e-07, 3.780872e-07, 3.736143e-07, 3.557728e-07, 3.649292e-07, 
    3.125342e-07, 3.350888e-07, 2.749348e-07, 2.909818e-07, 4.147556e-07, 
    4.083346e-07, 3.864558e-07, 3.967749e-07, 3.67706e-07, 3.607573e-07, 
    3.551696e-07, 3.481038e-07, 3.47347e-07, 3.432079e-07, 3.500066e-07, 
    3.434752e-07, 3.685858e-07, 3.572289e-07, 3.889209e-07, 3.810545e-07, 
    3.846615e-07, 3.886412e-07, 3.764389e-07, 3.636986e-07, 3.63431e-07, 
    3.594044e-07, 3.482039e-07, 3.67591e-07, 3.096925e-07, 3.447133e-07, 
    4.014015e-07, 3.893278e-07, 3.876236e-07, 3.922613e-07, 3.614502e-07, 
    3.724357e-07, 3.433086e-07, 3.510362e-07, 3.38431e-07, 3.446587e-07, 
    3.455809e-07, 3.536974e-07, 3.588093e-07, 3.719272e-07, 3.828153e-07, 
    3.915868e-07, 3.895366e-07, 3.799387e-07, 3.629284e-07, 3.472778e-07, 
    3.506693e-07, 3.393789e-07, 3.697683e-07, 3.568279e-07, 3.617951e-07, 
    3.489325e-07, 3.77495e-07, 3.530799e-07, 3.838966e-07, 3.811316e-07, 
    3.726558e-07, 3.559593e-07, 3.523316e-07, 3.484806e-07, 3.508541e-07, 
    3.625031e-07, 3.644348e-07, 3.728608e-07, 3.752073e-07, 3.817327e-07, 
    3.871863e-07, 3.822012e-07, 3.770081e-07, 3.624989e-07, 3.497222e-07, 
    3.361161e-07, 3.328383e-07, 3.174591e-07, 3.299416e-07, 3.095037e-07, 
    3.268238e-07, 2.972201e-07, 3.516983e-07, 3.273454e-07, 3.722735e-07, 
    3.67261e-07, 3.58299e-07, 3.38263e-07, 3.489923e-07, 3.364659e-07, 
    3.645108e-07, 3.796093e-07, 3.835791e-07, 3.910498e-07, 3.834094e-07, 
    3.840274e-07, 3.767951e-07, 3.791101e-07, 3.620231e-07, 3.711414e-07, 
    3.456036e-07, 3.365641e-07, 3.11844e-07, 2.972754e-07, 2.829032e-07, 
    2.767029e-07, 2.748335e-07, 2.740543e-07,
  1.268738e-08, 1.195778e-08, 1.209717e-08, 1.152653e-08, 1.184061e-08, 
    1.147054e-08, 1.253694e-08, 1.192943e-08, 1.231473e-08, 1.262045e-08, 
    1.047571e-08, 1.150155e-08, 9.483516e-09, 1.008415e-08, 8.626414e-09, 
    9.575157e-09, 8.443963e-09, 8.652818e-09, 8.035792e-09, 8.209075e-09, 
    7.456517e-09, 7.956749e-09, 7.092816e-09, 7.573791e-09, 7.496101e-09, 
    7.973661e-09, 1.128949e-08, 1.059958e-08, 1.133136e-08, 1.123075e-08, 
    1.127583e-08, 1.183404e-08, 1.212283e-08, 1.27445e-08, 1.262996e-08, 
    1.217421e-08, 1.118572e-08, 1.151446e-08, 1.069937e-08, 1.07173e-08, 
    9.859638e-09, 1.02398e-08, 8.875845e-09, 9.248867e-09, 8.201788e-09, 
    8.456303e-09, 8.213603e-09, 8.286644e-09, 8.212655e-09, 8.588306e-09, 
    8.425814e-09, 8.762074e-09, 1.016778e-08, 9.73845e-09, 1.105999e-08, 
    1.191538e-08, 1.250982e-08, 1.29445e-08, 1.288239e-08, 1.276457e-08, 
    1.217158e-08, 1.163268e-08, 1.123388e-08, 1.097276e-08, 1.071988e-08, 
    9.980396e-09, 9.604773e-09, 8.801772e-09, 8.942897e-09, 8.704842e-09, 
    8.481945e-09, 8.117296e-09, 8.176499e-09, 8.018762e-09, 8.711099e-09, 
    8.246174e-09, 9.024022e-09, 8.806045e-09, 1.065164e-08, 1.14251e-08, 
    1.176581e-08, 1.207027e-08, 1.283478e-08, 1.230316e-08, 1.251077e-08, 
    1.202105e-08, 1.171721e-08, 1.186678e-08, 1.096568e-08, 1.13098e-08, 
    9.582843e-09, 1.030088e-08, 8.507721e-09, 8.913799e-09, 8.412487e-09, 
    8.665595e-09, 8.235306e-09, 8.621823e-09, 7.960659e-09, 7.821868e-09, 
    7.91651e-09, 7.557664e-09, 8.643634e-09, 8.213585e-09, 1.187098e-08, 
    1.184649e-08, 1.173287e-08, 1.223828e-08, 1.226972e-08, 1.274764e-08, 
    1.232176e-08, 1.214357e-08, 1.169979e-08, 1.14429e-08, 1.120258e-08, 
    1.068724e-08, 1.013253e-08, 9.393002e-09, 8.887043e-09, 8.559451e-09, 
    8.759249e-09, 8.582675e-09, 8.780234e-09, 8.873998e-09, 7.873645e-09, 
    8.424299e-09, 7.608508e-09, 7.652034e-09, 8.015031e-09, 7.64712e-09, 
    1.182931e-08, 1.197063e-08, 1.247079e-08, 1.20781e-08, 1.280049e-08, 
    1.239233e-08, 1.216197e-08, 1.130248e-08, 1.111983e-08, 1.095234e-08, 
    1.062706e-08, 1.022008e-08, 9.534113e-09, 8.965627e-09, 8.469119e-09, 
    8.504786e-09, 8.492215e-09, 8.383927e-09, 8.654044e-09, 8.340193e-09, 
    8.288349e-09, 8.424388e-09, 7.657877e-09, 7.871278e-09, 7.652961e-09, 
    7.791344e-09, 1.192457e-08, 1.168816e-08, 1.181547e-08, 1.157689e-08, 
    1.174458e-08, 1.101229e-08, 1.079943e-08, 9.8435e-09, 1.022797e-08, 
    9.621242e-09, 1.01651e-08, 1.00671e-08, 9.60182e-09, 1.013516e-08, 
    8.996257e-09, 9.757284e-09, 8.379739e-09, 9.10084e-09, 8.336017e-09, 
    8.47122e-09, 8.248269e-09, 8.052331e-09, 7.810856e-09, 7.379605e-09, 
    7.477835e-09, 7.127736e-09, 1.134215e-08, 1.104722e-08, 1.107301e-08, 
    1.076995e-08, 1.054978e-08, 1.008403e-08, 9.368974e-09, 9.63331e-09, 
    9.152242e-09, 9.057849e-09, 9.790404e-09, 9.335579e-09, 1.085305e-08, 
    1.059632e-08, 1.074866e-08, 1.131865e-08, 9.571856e-09, 1.044131e-08, 
    8.878849e-09, 9.317876e-09, 8.080047e-09, 8.679132e-09, 7.532321e-09, 
    7.083668e-09, 6.674738e-09, 6.219872e-09, 1.088871e-08, 1.108637e-08, 
    1.073434e-08, 1.026086e-08, 9.835631e-09, 9.290637e-09, 9.236192e-09, 
    9.137066e-09, 8.884036e-09, 8.675348e-09, 9.105851e-09, 8.623616e-09, 
    1.053733e-08, 9.499026e-09, 1.116174e-08, 1.064009e-08, 1.028836e-08, 
    1.044162e-08, 9.663881e-09, 9.486994e-09, 8.792838e-09, 9.146795e-09, 
    7.188499e-09, 8.011344e-09, 5.889936e-09, 6.435146e-09, 1.115604e-08, 
    1.088941e-08, 9.997854e-09, 1.041506e-08, 9.255094e-09, 8.984921e-09, 
    8.769692e-09, 8.500136e-09, 8.471437e-09, 8.315081e-09, 8.572438e-09, 
    8.325149e-09, 9.289502e-09, 8.848801e-09, 1.009698e-08, 9.781846e-09, 
    9.925916e-09, 1.008571e-08, 9.598565e-09, 9.098943e-09, 9.088548e-09, 
    8.932642e-09, 8.503931e-09, 9.2506e-09, 7.092244e-09, 8.371833e-09, 
    1.060403e-08, 1.011338e-08, 1.004477e-08, 1.023185e-08, 9.011737e-09, 
    9.440576e-09, 8.318874e-09, 8.611651e-09, 8.1359e-09, 8.369772e-09, 
    8.404599e-09, 8.713285e-09, 8.909682e-09, 9.420575e-09, 9.852084e-09, 
    1.020456e-08, 1.012179e-08, 9.737428e-09, 9.069038e-09, 8.468813e-09, 
    8.597669e-09, 8.171349e-09, 9.335812e-09, 8.833375e-09, 9.025095e-09, 
    8.531598e-09, 9.640394e-09, 8.689665e-09, 9.895302e-09, 9.784918e-09, 
    9.44924e-09, 8.8e-09, 8.66107e-09, 8.514434e-09, 8.604709e-09, 
    9.052539e-09, 9.127561e-09, 9.457311e-09, 9.549862e-09, 9.808877e-09, 
    1.002719e-08, 9.82757e-09, 9.621099e-09, 9.052373e-09, 8.561618e-09, 
    8.049558e-09, 7.927849e-09, 7.36551e-09, 7.820831e-09, 7.085502e-09, 
    7.706214e-09, 6.651701e-09, 8.636897e-09, 7.725347e-09, 9.434193e-09, 
    9.237707e-09, 8.890005e-09, 8.129622e-09, 8.53387e-09, 8.062583e-09, 
    9.130514e-09, 9.724329e-09, 9.882608e-09, 1.018286e-08, 9.875821e-09, 
    9.900537e-09, 9.612665e-09, 9.704491e-09, 9.033931e-09, 9.389692e-09, 
    8.405459e-09, 8.066241e-09, 7.163813e-09, 6.653632e-09, 6.158517e-09, 
    5.949162e-09, 5.886549e-09, 5.860524e-09,
  8.754802e-11, 7.986248e-11, 8.131315e-11, 7.542873e-11, 7.864973e-11, 
    7.485913e-11, 8.594478e-11, 7.956852e-11, 8.359412e-11, 8.683354e-11, 
    6.498137e-11, 7.517444e-11, 5.561127e-11, 6.122404e-11, 4.793567e-11, 
    5.645551e-11, 4.635502e-11, 4.816602e-11, 4.288975e-11, 4.434875e-11, 
    3.814694e-11, 4.223028e-11, 3.20723e-11, 3.909003e-11, 3.846427e-11, 
    4.237106e-11, 7.302717e-11, 6.618576e-11, 7.344949e-11, 7.243599e-11, 
    7.288952e-11, 7.858185e-11, 8.158111e-11, 8.81592e-11, 8.693499e-11, 
    8.211853e-11, 7.198393e-11, 7.530578e-11, 6.716138e-11, 6.733714e-11, 
    5.910426e-11, 6.270853e-11, 5.012742e-11, 5.346994e-11, 4.428703e-11, 
    4.646132e-11, 4.438711e-11, 4.500769e-11, 4.437908e-11, 4.760394e-11, 
    4.619884e-11, 4.912334e-11, 6.202012e-11, 5.797078e-11, 7.072659e-11, 
    7.942292e-11, 8.565676e-11, 9.030988e-11, 8.964021e-11, 8.837432e-11, 
    8.209098e-11, 7.651239e-11, 7.246741e-11, 6.985851e-11, 6.736244e-11, 
    6.024123e-11, 5.67293e-11, 4.947287e-11, 5.072258e-11, 4.862102e-11, 
    4.668248e-11, 4.357374e-11, 4.407309e-11, 4.274734e-11, 4.867585e-11, 
    4.466346e-11, 5.1446e-11, 4.951054e-11, 6.669415e-11, 7.439789e-11, 
    7.787856e-11, 8.103259e-11, 8.912796e-11, 8.347234e-11, 8.566681e-11, 
    8.051993e-11, 7.737894e-11, 7.89201e-11, 6.978826e-11, 7.323196e-11, 
    5.652653e-11, 6.329434e-11, 4.690519e-11, 5.0464e-11, 4.608428e-11, 
    4.827762e-11, 4.457117e-11, 4.789566e-11, 4.226281e-11, 4.111381e-11, 
    4.189603e-11, 3.895981e-11, 4.808585e-11, 4.438696e-11, 7.896352e-11, 
    7.871039e-11, 7.753988e-11, 8.279035e-11, 8.312062e-11, 8.819281e-11, 
    8.366822e-11, 8.179799e-11, 7.720011e-11, 7.457851e-11, 7.215303e-11, 
    6.704247e-11, 6.168416e-11, 5.478178e-11, 5.022665e-11, 4.735331e-11, 
    4.909851e-11, 4.755499e-11, 4.928313e-11, 5.011107e-11, 4.154106e-11, 
    4.618581e-11, 3.93709e-11, 3.972413e-11, 4.271617e-11, 3.968419e-11, 
    7.853306e-11, 7.999591e-11, 8.524279e-11, 8.111423e-11, 8.875965e-11, 
    8.441267e-11, 8.199041e-11, 7.315808e-11, 7.132409e-11, 6.965591e-11, 
    6.645397e-11, 6.251981e-11, 5.607685e-11, 5.092491e-11, 4.657181e-11, 
    4.687982e-11, 4.677117e-11, 4.583913e-11, 4.817672e-11, 4.546467e-11, 
    4.50222e-11, 4.618659e-11, 3.977164e-11, 4.15215e-11, 3.973167e-11, 
    4.086272e-11, 7.951811e-11, 7.708077e-11, 7.839027e-11, 7.594218e-11, 
    7.766022e-11, 7.025147e-11, 6.814439e-11, 5.895289e-11, 6.259526e-11, 
    5.688175e-11, 6.199454e-11, 6.106213e-11, 5.670198e-11, 6.170914e-11, 
    5.1198e-11, 5.814643e-11, 4.580323e-11, 5.213437e-11, 4.542897e-11, 
    4.658994e-11, 4.468125e-11, 4.302822e-11, 4.102316e-11, 3.753326e-11, 
    3.831772e-11, 3.555076e-11, 7.355842e-11, 7.059929e-11, 7.085636e-11, 
    6.785431e-11, 6.570065e-11, 6.122285e-11, 5.456232e-11, 5.699355e-11, 
    5.259678e-11, 5.174872e-11, 5.845578e-11, 5.425781e-11, 6.867319e-11, 
    6.615392e-11, 6.764504e-11, 7.332117e-11, 5.642503e-11, 6.464829e-11, 
    5.015403e-11, 5.409663e-11, 4.326065e-11, 4.839596e-11, 3.875553e-11, 
    3.201885e-11, 2.964211e-11, 2.702909e-11, 6.902557e-11, 7.098978e-11, 
    6.750435e-11, 6.291032e-11, 5.887912e-11, 5.384895e-11, 5.335511e-11, 
    5.246011e-11, 5.019999e-11, 4.836287e-11, 5.217939e-11, 4.791129e-11, 
    6.55796e-11, 5.575384e-11, 7.174356e-11, 6.658119e-11, 6.317408e-11, 
    6.465128e-11, 5.727709e-11, 5.564324e-11, 4.939413e-11, 5.254772e-11, 
    3.602519e-11, 4.268538e-11, 2.515545e-11, 2.826157e-11, 7.168644e-11, 
    6.903247e-11, 6.040621e-11, 6.439446e-11, 5.352638e-11, 5.109687e-11, 
    4.919035e-11, 4.683962e-11, 4.65918e-11, 4.525015e-11, 4.746605e-11, 
    4.533611e-11, 5.383864e-11, 4.988809e-11, 6.134594e-11, 5.837579e-11, 
    5.972737e-11, 6.123888e-11, 5.667187e-11, 5.211732e-11, 5.2024e-11, 
    5.06314e-11, 4.687242e-11, 5.348565e-11, 3.206896e-11, 4.573546e-11, 
    6.622917e-11, 6.150182e-11, 6.085036e-11, 6.263237e-11, 5.133622e-11, 
    5.521722e-11, 4.528253e-11, 4.780706e-11, 4.373043e-11, 4.571781e-11, 
    4.601652e-11, 4.869501e-11, 5.042745e-11, 5.503401e-11, 5.903338e-11, 
    6.23714e-11, 6.158189e-11, 5.796124e-11, 5.1849e-11, 4.656917e-11, 
    4.768537e-11, 4.402956e-11, 5.425993e-11, 4.975175e-11, 5.14556e-11, 
    4.711183e-11, 5.705921e-11, 4.848811e-11, 5.943927e-11, 5.84045e-11, 
    5.529664e-11, 4.945725e-11, 4.823808e-11, 4.696326e-11, 4.774662e-11, 
    5.170117e-11, 5.237457e-11, 5.537068e-11, 5.622204e-11, 5.862857e-11, 
    6.068383e-11, 5.880359e-11, 5.688043e-11, 5.169968e-11, 4.737212e-11, 
    4.3005e-11, 4.199013e-11, 3.74212e-11, 4.110527e-11, 3.202957e-11, 
    4.016549e-11, 2.950898e-11, 4.802708e-11, 4.032179e-11, 5.515873e-11, 
    5.336883e-11, 5.02529e-11, 4.367753e-11, 4.713152e-11, 4.311414e-11, 
    5.240115e-11, 5.783919e-11, 5.931996e-11, 6.216405e-11, 5.92562e-11, 
    5.94885e-11, 5.680233e-11, 5.765451e-11, 5.153462e-11, 5.475153e-11, 
    4.602391e-11, 4.314481e-11, 3.583215e-11, 2.952014e-11, 2.667925e-11, 
    2.549038e-11, 2.513632e-11, 2.498936e-11,
  8.438734e-14, 7.197419e-14, 7.428547e-14, 6.500878e-14, 7.005394e-14, 
    6.412516e-14, 8.176462e-14, 7.150772e-14, 7.79502e-14, 8.321646e-14, 
    4.925325e-14, 6.461399e-14, 3.606517e-14, 4.384528e-14, 2.610349e-14, 
    3.721081e-14, 2.416484e-14, 2.638947e-14, 2.006976e-14, 2.176686e-14, 
    1.485465e-14, 1.931625e-14, 1.189426e-14, 1.585229e-14, 1.518802e-14, 
    1.947638e-14, 6.130145e-14, 5.101774e-14, 6.194992e-14, 6.039626e-14, 
    6.109043e-14, 6.994678e-14, 7.471407e-14, 8.539158e-14, 8.338251e-14, 
    7.557523e-14, 5.970612e-14, 6.481783e-14, 5.245761e-14, 5.271798e-14, 
    4.086279e-14, 4.596393e-14, 2.885909e-14, 3.320133e-14, 2.169426e-14, 
    2.429388e-14, 2.181204e-14, 2.254646e-14, 2.180257e-14, 2.569314e-14, 
    2.397561e-14, 2.758727e-14, 4.497844e-14, 3.928953e-14, 5.779594e-14, 
    7.127692e-14, 8.129524e-14, 8.894423e-14, 8.783492e-14, 8.574563e-14, 
    7.553103e-14, 6.669706e-14, 6.04443e-14, 5.648536e-14, 5.275548e-14, 
    4.245609e-14, 3.758429e-14, 2.802821e-14, 2.962026e-14, 2.695693e-14, 
    2.456299e-14, 2.086031e-14, 2.144312e-14, 1.990632e-14, 2.702554e-14, 
    2.21382e-14, 3.055261e-14, 2.807586e-14, 5.176689e-14, 6.341162e-14, 
    6.883868e-14, 7.383726e-14, 8.698824e-14, 7.775361e-14, 8.131162e-14, 
    7.301977e-14, 6.805378e-14, 7.048108e-14, 5.637958e-14, 6.161571e-14, 
    3.730759e-14, 4.680655e-14, 2.483482e-14, 2.928889e-14, 2.383706e-14, 
    2.652835e-14, 2.202912e-14, 2.60539e-14, 1.935322e-14, 1.806065e-14, 
    1.893767e-14, 1.571333e-14, 2.628984e-14, 2.181186e-14, 7.054973e-14, 
    7.014972e-14, 6.83064e-14, 7.665463e-14, 7.718644e-14, 8.544689e-14, 
    7.806987e-14, 7.506134e-14, 6.77733e-14, 6.369084e-14, 5.996406e-14, 
    5.228162e-14, 4.449938e-14, 3.494854e-14, 2.898562e-14, 2.538434e-14, 
    2.755601e-14, 2.563276e-14, 2.77886e-14, 2.883825e-14, 1.853811e-14, 
    2.395983e-14, 1.615337e-14, 1.653454e-14, 1.98706e-14, 1.64913e-14, 
    6.98698e-14, 7.218613e-14, 8.062157e-14, 7.396762e-14, 8.638052e-14, 
    7.927421e-14, 7.536974e-14, 6.150232e-14, 5.870195e-14, 5.618044e-14, 
    5.141267e-14, 4.569325e-14, 3.669584e-14, 2.988024e-14, 2.442822e-14, 
    2.480381e-14, 2.467114e-14, 2.354137e-14, 2.640278e-14, 2.309175e-14, 
    2.256372e-14, 2.396077e-14, 1.658601e-14, 1.851616e-14, 1.65427e-14, 
    1.778183e-14, 7.14278e-14, 6.758628e-14, 6.964455e-14, 6.580752e-14, 
    6.849542e-14, 5.707778e-14, 5.391766e-14, 4.06518e-14, 4.580143e-14, 
    3.779265e-14, 4.494193e-14, 4.361569e-14, 3.754697e-14, 4.453496e-14, 
    3.023212e-14, 3.953232e-14, 2.349815e-14, 3.144691e-14, 2.304902e-14, 
    2.445028e-14, 2.215925e-14, 2.022907e-14, 1.795983e-14, 1.421674e-14, 
    1.503376e-14, 1.221992e-14, 6.211742e-14, 5.760332e-14, 5.799245e-14, 
    5.348585e-14, 5.030529e-14, 4.384359e-14, 3.465463e-14, 3.794565e-14, 
    3.205151e-14, 3.094505e-14, 3.996083e-14, 3.424788e-14, 5.470687e-14, 
    5.097091e-14, 5.317484e-14, 6.175273e-14, 3.716929e-14, 4.876785e-14, 
    2.8893e-14, 3.40331e-14, 2.049731e-14, 2.667583e-14, 1.549608e-14, 
    1.182557e-14, 8.950257e-15, 6.213803e-15, 5.523424e-14, 5.819463e-14, 
    5.296597e-14, 4.625377e-14, 4.054908e-14, 3.370374e-14, 3.304951e-14, 
    3.187249e-14, 2.895162e-14, 2.663457e-14, 3.150564e-14, 2.607327e-14, 
    5.012787e-14, 3.625799e-14, 5.933987e-14, 5.160021e-14, 4.663327e-14, 
    4.877221e-14, 3.833437e-14, 3.610838e-14, 2.792871e-14, 3.198721e-14, 
    1.268861e-14, 1.983532e-14, 4.543956e-15, 7.447048e-15, 5.925291e-14, 
    5.524458e-14, 4.268853e-14, 4.839871e-14, 3.327602e-14, 3.010168e-14, 
    2.767165e-14, 2.47547e-14, 2.445255e-14, 2.283531e-14, 2.552312e-14, 
    2.293798e-14, 3.369003e-14, 2.855452e-14, 4.401834e-14, 3.984992e-14, 
    4.173413e-14, 4.386634e-14, 3.750587e-14, 3.142469e-14, 3.130306e-14, 
    2.95033e-14, 2.479476e-14, 3.322211e-14, 1.188996e-14, 2.341664e-14, 
    5.108162e-14, 4.423988e-14, 4.33158e-14, 4.585465e-14, 3.041063e-14, 
    3.553358e-14, 2.287396e-14, 2.594418e-14, 2.104268e-14, 2.339543e-14, 
    2.375523e-14, 2.704952e-14, 2.924214e-14, 3.528712e-14, 4.076396e-14, 
    4.548067e-14, 4.43538e-14, 3.927636e-14, 3.107533e-14, 2.442501e-14, 
    2.57937e-14, 2.139213e-14, 3.425071e-14, 2.838141e-14, 3.056503e-14, 
    2.50878e-14, 3.803558e-14, 2.679083e-14, 4.13307e-14, 3.988971e-14, 
    3.564057e-14, 2.800847e-14, 2.647913e-14, 2.490584e-14, 2.586942e-14, 
    3.088331e-14, 3.176059e-14, 3.574037e-14, 3.689308e-14, 4.020067e-14, 
    4.308036e-14, 4.044396e-14, 3.779085e-14, 3.088138e-14, 2.540747e-14, 
    2.020233e-14, 1.904402e-14, 1.410124e-14, 1.805114e-14, 1.183932e-14, 
    1.701468e-14, 8.799815e-15, 2.621686e-14, 1.718575e-14, 3.545485e-14, 
    3.306765e-14, 2.901912e-14, 2.098106e-14, 2.511194e-14, 2.032811e-14, 
    3.179534e-14, 3.910789e-14, 4.11639e-14, 4.518406e-14, 4.107484e-14, 
    4.139957e-14, 3.768408e-14, 3.885331e-14, 3.066735e-14, 3.490799e-14, 
    2.376415e-14, 2.03635e-14, 1.249719e-14, 8.812384e-15, 5.882961e-15, 
    4.823847e-15, 4.52822e-15, 4.408219e-15,
  2.852239e-19, 2.437973e-19, 2.515188e-19, 2.20503e-19, 2.373791e-19, 
    2.175452e-19, 2.764796e-19, 2.422384e-19, 2.637542e-19, 2.813206e-19, 
    1.676607e-19, 2.191815e-19, 1.232317e-19, 1.494668e-19, 8.952005e-20, 
    1.270998e-19, 8.293947e-20, 9.04902e-20, 6.901305e-20, 7.478905e-20, 
    5.121712e-20, 6.644629e-20, 4.111686e-20, 5.462747e-20, 5.235706e-20, 
    6.699188e-20, 2.080889e-19, 1.735902e-19, 2.102611e-19, 2.050561e-19, 
    2.073819e-19, 2.370209e-19, 2.529503e-19, 2.885708e-19, 2.818742e-19, 
    2.55826e-19, 2.027433e-19, 2.198639e-19, 1.784265e-19, 1.793009e-19, 
    1.394185e-19, 1.565983e-19, 9.886149e-20, 1.135553e-19, 7.454207e-20, 
    8.337774e-20, 7.494271e-20, 7.744016e-20, 7.491052e-20, 8.812779e-20, 
    8.229674e-20, 9.455175e-20, 1.532817e-19, 1.341137e-19, 1.963399e-19, 
    2.414671e-19, 2.749142e-19, 3.004063e-19, 2.967115e-19, 2.897507e-19, 
    2.556784e-19, 2.261525e-19, 2.05217e-19, 1.919445e-19, 1.794268e-19, 
    1.447878e-19, 1.283604e-19, 9.604628e-20, 1.014395e-19, 9.24147e-20, 
    8.429159e-20, 7.170449e-20, 7.368771e-20, 6.84564e-20, 9.264733e-20, 
    7.605199e-20, 1.045959e-19, 9.620775e-20, 1.761068e-19, 2.151562e-19, 
    2.333159e-19, 2.500218e-19, 2.93891e-19, 2.630981e-19, 2.749689e-19, 
    2.472908e-19, 2.306909e-19, 2.38807e-19, 1.915897e-19, 2.091416e-19, 
    1.274264e-19, 1.594333e-19, 8.521452e-20, 1.003173e-19, 8.182613e-20, 
    9.096125e-20, 7.568104e-20, 8.935183e-20, 6.657225e-20, 6.216602e-20, 
    6.515616e-20, 5.41526e-20, 9.015224e-20, 7.49421e-20, 2.390365e-19, 
    2.376993e-19, 2.315358e-19, 2.594298e-19, 2.61205e-19, 2.887552e-19, 
    2.641536e-19, 2.5411e-19, 2.297528e-19, 2.160911e-19, 2.036078e-19, 
    1.778355e-19, 1.51669e-19, 1.194598e-19, 9.92901e-20, 8.707982e-20, 
    9.444581e-20, 8.792287e-20, 9.52342e-20, 9.87909e-20, 6.379413e-20, 
    8.224316e-20, 5.565606e-20, 5.695789e-20, 6.833474e-20, 5.681025e-20, 
    2.367635e-19, 2.445055e-19, 2.726673e-19, 2.504572e-19, 2.918662e-19, 
    2.681724e-19, 2.551398e-19, 2.087618e-19, 1.993775e-19, 1.909217e-19, 
    1.749169e-19, 1.556875e-19, 1.253613e-19, 1.023198e-19, 8.383393e-20, 
    8.510924e-20, 8.465881e-20, 8.082157e-20, 9.053534e-20, 7.929371e-20, 
    7.749884e-20, 8.224635e-20, 5.713367e-20, 6.371931e-20, 5.698577e-20, 
    6.121499e-20, 2.419713e-19, 2.291272e-19, 2.360104e-19, 2.231761e-19, 
    2.32168e-19, 1.939316e-19, 1.833286e-19, 1.387073e-19, 1.560515e-19, 
    1.290636e-19, 1.531588e-19, 1.486936e-19, 1.282344e-19, 1.517888e-19, 
    1.03511e-19, 1.349326e-19, 8.067472e-20, 1.076221e-19, 7.914847e-20, 
    8.390885e-20, 7.612357e-20, 6.955554e-20, 6.182216e-20, 4.903484e-20, 
    5.182963e-20, 4.219468e-20, 2.108222e-19, 1.95694e-19, 1.969988e-19, 
    1.81879e-19, 1.711964e-19, 1.494611e-19, 1.184667e-19, 1.295799e-19, 
    1.096673e-19, 1.05924e-19, 1.363776e-19, 1.170922e-19, 1.859774e-19, 
    1.734329e-19, 1.808348e-19, 2.096006e-19, 1.269596e-19, 1.66029e-19, 
    9.897637e-20, 1.163665e-19, 7.046883e-20, 9.146144e-20, 5.341013e-20, 
    4.0881e-20, 3.099038e-20, 2.153798e-20, 1.877471e-19, 1.976767e-19, 
    1.801336e-19, 1.575736e-19, 1.38361e-19, 1.152534e-19, 1.13042e-19, 
    1.090618e-19, 9.917492e-20, 9.13215e-20, 1.078208e-19, 8.941755e-20, 
    1.706002e-19, 1.238828e-19, 2.015158e-19, 1.755469e-19, 1.588503e-19, 
    1.660436e-19, 1.308915e-19, 1.233776e-19, 9.570906e-20, 1.094498e-19, 
    4.380148e-20, 6.821459e-20, 1.57446e-20, 2.580329e-20, 2.012243e-19, 
    1.877818e-19, 1.455709e-19, 1.647879e-19, 1.138077e-19, 1.030695e-19, 
    9.483778e-20, 8.494249e-20, 8.391657e-20, 7.842209e-20, 8.755083e-20, 
    7.877106e-20, 1.152071e-19, 9.782968e-20, 1.500495e-19, 1.360036e-19, 
    1.423552e-19, 1.495376e-19, 1.280957e-19, 1.075469e-19, 1.071355e-19, 
    1.010434e-19, 8.507851e-20, 1.136255e-19, 4.110209e-20, 8.039777e-20, 
    1.738048e-19, 1.507954e-19, 1.476837e-19, 1.562306e-19, 1.041153e-19, 
    1.214363e-19, 7.855348e-20, 8.897958e-20, 7.232514e-20, 8.032569e-20, 
    8.154814e-20, 9.272867e-20, 1.00159e-19, 1.206037e-19, 1.390854e-19, 
    1.549721e-19, 1.511789e-19, 1.340693e-19, 1.063649e-19, 8.382305e-20, 
    8.8469e-20, 7.351424e-20, 1.171018e-19, 9.724315e-20, 1.046379e-19, 
    8.607331e-20, 1.298834e-19, 9.185145e-20, 1.409957e-19, 1.361378e-19, 
    1.217976e-19, 9.597937e-20, 9.07943e-20, 8.545563e-20, 8.872591e-20, 
    1.057151e-19, 1.086833e-19, 1.221347e-19, 1.260272e-19, 1.371864e-19, 
    1.468907e-19, 1.380066e-19, 1.290575e-19, 1.057086e-19, 8.715834e-20, 
    6.946448e-20, 6.55186e-20, 4.863958e-20, 6.213359e-20, 4.092824e-20, 
    5.859719e-20, 3.047181e-20, 8.990468e-20, 5.918108e-20, 1.211703e-19, 
    1.131033e-19, 9.940358e-20, 7.211543e-20, 8.615526e-20, 6.989274e-20, 
    1.088008e-19, 1.335011e-19, 1.404335e-19, 1.539738e-19, 1.401333e-19, 
    1.412278e-19, 1.286972e-19, 1.326424e-19, 1.049842e-19, 1.193228e-19, 
    8.157843e-20, 7.001326e-20, 4.314534e-20, 3.051514e-20, 2.039194e-20, 
    1.671733e-20, 1.56899e-20, 1.52726e-20,
  2.093585e-25, 1.790998e-25, 1.847414e-25, 1.62075e-25, 1.744098e-25, 
    1.599127e-25, 2.029733e-25, 1.779607e-25, 1.936794e-25, 2.065084e-25, 
    1.234212e-25, 1.61109e-25, 9.087386e-26, 1.100992e-25, 6.613274e-26, 
    9.370968e-26, 6.129759e-26, 6.68454e-26, 5.105741e-26, 5.530588e-26, 
    3.795339e-26, 4.91688e-26, 3.051394e-26, 4.046651e-26, 3.879353e-26, 
    4.957028e-26, 1.529987e-25, 1.277613e-25, 1.545871e-25, 1.50781e-25, 
    1.524818e-25, 1.74148e-25, 1.857872e-25, 2.118023e-25, 2.069126e-25, 
    1.87888e-25, 1.490896e-25, 1.616078e-25, 1.313007e-25, 1.319405e-25, 
    1.02738e-25, 1.15322e-25, 7.299307e-26, 8.377705e-26, 5.512425e-26, 
    6.161967e-26, 5.541887e-26, 5.725521e-26, 5.53952e-26, 6.510994e-26, 
    6.082521e-26, 6.982848e-26, 1.128932e-25, 9.885074e-26, 1.444063e-25, 
    1.773971e-25, 2.018301e-25, 2.204429e-25, 2.177456e-25, 2.126637e-25, 
    1.877802e-25, 1.662048e-25, 1.508987e-25, 1.411912e-25, 1.320327e-25, 
    1.066718e-25, 9.463378e-26, 7.092599e-26, 7.48857e-26, 6.825898e-26, 
    6.229124e-26, 5.303732e-26, 5.449595e-26, 5.064787e-26, 6.842984e-26, 
    5.623456e-26, 7.72026e-26, 7.104456e-26, 1.296031e-25, 1.581662e-25, 
    1.714404e-25, 1.836477e-25, 2.156865e-25, 1.932001e-25, 2.0187e-25, 
    1.816524e-25, 1.695219e-25, 1.754533e-25, 1.409316e-25, 1.537685e-25, 
    9.394917e-26, 1.173979e-25, 6.296944e-26, 7.406187e-26, 6.047933e-26, 
    6.719141e-26, 5.59618e-26, 6.600917e-26, 4.926149e-26, 4.60184e-26, 
    4.821935e-26, 4.011664e-26, 6.659715e-26, 5.541843e-26, 1.75621e-25, 
    1.746438e-25, 1.701394e-25, 1.905206e-25, 1.918173e-25, 2.119368e-25, 
    1.939711e-25, 1.866344e-25, 1.688363e-25, 1.588497e-25, 1.497218e-25, 
    1.308682e-25, 1.117122e-25, 8.810807e-26, 7.330776e-26, 6.434e-26, 
    6.975068e-26, 6.495939e-26, 7.032966e-26, 7.294125e-26, 4.721688e-26, 
    6.078582e-26, 4.12243e-26, 4.218327e-26, 5.055835e-26, 4.207452e-26, 
    1.7396e-25, 1.796173e-25, 2.001892e-25, 1.839658e-25, 2.142083e-25, 
    1.969064e-25, 1.873868e-25, 1.534908e-25, 1.46628e-25, 1.404429e-25, 
    1.287323e-25, 1.14655e-25, 9.243518e-26, 7.553188e-26, 6.195492e-26, 
    6.289208e-26, 6.256109e-26, 5.974097e-26, 6.687856e-26, 5.861788e-26, 
    5.729836e-26, 6.078817e-26, 4.231274e-26, 4.716181e-26, 4.22038e-26, 
    4.531823e-26, 1.777656e-25, 1.68379e-25, 1.734096e-25, 1.640291e-25, 
    1.706015e-25, 1.426447e-25, 1.348877e-25, 1.022169e-25, 1.149216e-25, 
    9.514927e-26, 1.128032e-25, 1.095329e-25, 9.454147e-26, 1.117999e-25, 
    7.640634e-26, 9.945085e-26, 5.963303e-26, 7.942362e-26, 5.851111e-26, 
    6.200998e-26, 5.628719e-26, 5.145652e-26, 4.576525e-26, 3.634468e-26, 
    3.840483e-26, 3.129927e-26, 1.549973e-25, 1.439338e-25, 1.448882e-25, 
    1.338271e-25, 1.260093e-25, 1.10095e-25, 8.737979e-26, 9.552773e-26, 
    8.09244e-26, 7.817739e-26, 1.005098e-25, 8.637174e-26, 1.368258e-25, 
    1.276462e-25, 1.33063e-25, 1.541041e-25, 9.360694e-26, 1.222267e-25, 
    7.307742e-26, 8.583936e-26, 5.212839e-26, 6.755881e-26, 3.956956e-26, 
    3.03398e-26, 2.303061e-26, 1.602984e-26, 1.381205e-25, 1.45384e-25, 
    1.325499e-25, 1.160361e-25, 1.019632e-25, 8.502284e-26, 8.340051e-26, 
    8.04801e-26, 7.32232e-26, 6.745602e-26, 7.956941e-26, 6.605744e-26, 
    1.255729e-25, 9.135128e-26, 1.481919e-25, 1.291934e-25, 1.16971e-25, 
    1.222375e-25, 9.648915e-26, 9.098085e-26, 7.067836e-26, 8.076482e-26, 
    3.248492e-26, 5.046996e-26, 1.172844e-26, 1.919122e-26, 1.479787e-25, 
    1.381459e-25, 1.072454e-25, 1.213182e-25, 8.396227e-26, 7.608223e-26, 
    7.003853e-26, 6.276955e-26, 6.201565e-26, 5.797712e-26, 6.468605e-26, 
    5.823366e-26, 8.498888e-26, 7.22355e-26, 1.10526e-25, 1.002357e-25, 
    1.048897e-25, 1.101511e-25, 9.443978e-26, 7.936844e-26, 7.906645e-26, 
    7.459493e-26, 6.28695e-26, 8.382859e-26, 3.050304e-26, 5.942945e-26, 
    1.279184e-25, 1.110723e-25, 1.087931e-25, 1.150527e-25, 7.684986e-26, 
    8.955739e-26, 5.807371e-26, 6.57357e-26, 5.349382e-26, 5.937648e-26, 
    6.027501e-26, 6.848958e-26, 7.394564e-26, 8.89469e-26, 1.024939e-25, 
    1.141311e-25, 1.113532e-25, 9.88182e-26, 7.850095e-26, 6.194692e-26, 
    6.536061e-26, 5.436838e-26, 8.637875e-26, 7.180484e-26, 7.723346e-26, 
    6.360047e-26, 9.575017e-26, 6.784527e-26, 1.038936e-25, 1.003341e-25, 
    8.982237e-26, 7.087686e-26, 6.706878e-26, 6.314661e-26, 6.554935e-26, 
    7.802405e-26, 8.020232e-26, 9.006953e-26, 9.292338e-26, 1.011024e-25, 
    1.082122e-25, 1.017035e-25, 9.51448e-26, 7.801926e-26, 6.439769e-26, 
    5.138953e-26, 4.84861e-26, 3.605326e-26, 4.599452e-26, 3.037468e-26, 
    4.339063e-26, 2.264699e-26, 6.641529e-26, 4.382062e-26, 8.936238e-26, 
    8.344548e-26, 7.339108e-26, 5.333958e-26, 6.366069e-26, 5.170459e-26, 
    8.028859e-26, 9.840173e-26, 1.034817e-25, 1.134001e-25, 1.032618e-25, 
    1.040637e-25, 9.488066e-26, 9.777237e-26, 7.748764e-26, 8.80076e-26, 
    6.029727e-26, 5.179325e-26, 3.200079e-26, 2.267904e-26, 1.517969e-26, 
    1.245136e-26, 1.168777e-26, 1.137753e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.01127981, 0.01129391, 0.01129116, 0.01130253, 0.01129622, 0.01130367, 
    0.01128266, 0.01129448, 0.01128693, 0.01128106, 0.01132457, 0.01130303, 
    0.01134671, 0.01133307, 0.01136723, 0.01134461, 0.01137178, 0.01136655, 
    0.01138219, 0.01137771, 0.01139774, 0.01138426, 0.01140803, 0.0113945, 
    0.01139663, 0.01138382, 0.01130734, 0.0113219, 0.01130649, 0.01130856, 
    0.01130763, 0.01129636, 0.01129069, 0.01127871, 0.01128088, 0.01128967, 
    0.0113095, 0.01130275, 0.01131967, 0.01131929, 0.01133808, 0.01132962, 
    0.01136109, 0.01135216, 0.0113779, 0.01137144, 0.0113776, 0.01137573, 
    0.01137763, 0.01136815, 0.01137221, 0.01136386, 0.01133121, 0.01134084, 
    0.0113121, 0.01129479, 0.01128318, 0.01127496, 0.01127612, 0.01127834, 
    0.01128972, 0.01130037, 0.01130848, 0.0113139, 0.01131924, 0.01133543, 
    0.01134391, 0.01136291, 0.01135946, 0.01136528, 0.0113708, 0.01138008, 
    0.01137855, 0.01138265, 0.01136511, 0.01137678, 0.0113575, 0.01136278, 
    0.01132079, 0.01130457, 0.01129775, 0.01129169, 0.01127702, 0.01128716, 
    0.01128317, 0.01129264, 0.01129868, 0.01129569, 0.01131405, 0.01130692, 
    0.01134442, 0.0113283, 0.01137015, 0.01136016, 0.01137254, 0.01136622, 
    0.01137705, 0.01136731, 0.01138416, 0.01138784, 0.01138533, 0.01139492, 
    0.01136677, 0.01137761, 0.01129561, 0.0112961, 0.01129836, 0.01128842, 
    0.01128781, 0.01127865, 0.01128679, 0.01129026, 0.01129902, 0.01130421, 
    0.01130913, 0.01131994, 0.01133201, 0.0113488, 0.01136081, 0.01136886, 
    0.01136392, 0.01136828, 0.01136341, 0.01136112, 0.01138647, 0.01137226, 
    0.01139354, 0.01139236, 0.01138275, 0.0113925, 0.01129644, 0.01129363, 
    0.01128392, 0.01129153, 0.01127766, 0.01128544, 0.01128991, 0.0113071, 
    0.01131084, 0.01131434, 0.01132122, 0.01133005, 0.01134552, 0.01135892, 
    0.01137111, 0.01137022, 0.01137054, 0.01137327, 0.01136651, 0.01137437, 
    0.0113757, 0.01137224, 0.01139221, 0.01138651, 0.01139234, 0.01138863, 
    0.01129454, 0.01129925, 0.01129671, 0.0113015, 0.01129813, 0.01131311, 
    0.01131759, 0.01133848, 0.01132989, 0.01134352, 0.01133126, 0.01133344, 
    0.01134401, 0.01133192, 0.01135821, 0.01134044, 0.01137337, 0.01135573, 
    0.01137448, 0.01137106, 0.01137671, 0.01138177, 0.01138811, 0.01139983, 
    0.01139711, 0.01140688, 0.01130626, 0.01131237, 0.01131181, 0.01131818, 
    0.01132289, 0.01133305, 0.01134935, 0.01134322, 0.01135444, 0.0113567, 
    0.01133964, 0.01135014, 0.01131643, 0.01132192, 0.01131864, 0.01130675, 
    0.01134466, 0.01132525, 0.01136102, 0.01135054, 0.01138105, 0.01136592, 
    0.01139562, 0.01140832, 0.01142015, 0.01143405, 0.01131567, 0.01131153, 
    0.01131893, 0.01132918, 0.01133863, 0.01135118, 0.01135245, 0.01135481, 
    0.01136088, 0.01136598, 0.01135557, 0.01136726, 0.01132323, 0.01134633, 
    0.01130998, 0.01132098, 0.01132857, 0.01132522, 0.01134251, 0.01134659, 
    0.01136312, 0.01135457, 0.01140521, 0.01138287, 0.01144453, 0.01142739, 
    0.01131009, 0.01131565, 0.01133499, 0.0113258, 0.01135201, 0.01135845, 
    0.01136366, 0.01137035, 0.01137106, 0.01137502, 0.01136853, 0.01137475, 
    0.01135121, 0.01136174, 0.01133276, 0.01133984, 0.01133658, 0.01133301, 
    0.01134401, 0.01135574, 0.01135596, 0.01135972, 0.01137036, 0.01135211, 
    0.01140814, 0.01137367, 0.01132171, 0.01133244, 0.01133393, 0.01132979, 
    0.01135781, 0.01134767, 0.01137491, 0.01136756, 0.0113796, 0.01137362, 
    0.01137274, 0.01136505, 0.01136026, 0.01134815, 0.01133826, 0.01133038, 
    0.01133221, 0.01134086, 0.01135645, 0.01137114, 0.01136793, 0.01137868, 
    0.01135011, 0.01136213, 0.0113575, 0.01136956, 0.01134306, 0.01136573, 
    0.01133727, 0.01133976, 0.01134747, 0.01136296, 0.01136634, 0.01136999, 
    0.01136773, 0.01135684, 0.01135504, 0.01134728, 0.01134515, 0.01133922, 
    0.01133431, 0.0113388, 0.01134352, 0.01135683, 0.01136882, 0.01138185, 
    0.01138502, 0.01140027, 0.0113879, 0.01140834, 0.01139104, 0.01142092, 
    0.01136699, 0.01139046, 0.01134781, 0.01135242, 0.01136077, 0.0113798, 
    0.0113695, 0.01138153, 0.01135497, 0.01134117, 0.01133755, 0.01133087, 
    0.01133771, 0.01133715, 0.01134369, 0.01134159, 0.01135727, 0.01134885, 
    0.01137273, 0.01138143, 0.01140587, 0.01142081, 0.01143593, 0.0114426, 
    0.01144463, 0.01144548,
  3.677391e-05, 3.686526e-05, 3.684746e-05, 3.692118e-05, 3.688023e-05, 
    3.692854e-05, 3.679235e-05, 3.686896e-05, 3.682002e-05, 3.678202e-05, 
    3.706501e-05, 3.692445e-05, 3.721029e-05, 3.712076e-05, 3.73452e-05, 
    3.719648e-05, 3.737511e-05, 3.734072e-05, 3.74437e-05, 3.74142e-05, 
    3.754615e-05, 3.745731e-05, 3.761411e-05, 3.752483e-05, 3.753888e-05, 
    3.74544e-05, 3.695242e-05, 3.704753e-05, 3.694687e-05, 3.696034e-05, 
    3.695425e-05, 3.688114e-05, 3.684439e-05, 3.676679e-05, 3.678085e-05, 
    3.683777e-05, 3.69664e-05, 3.692263e-05, 3.703298e-05, 3.703047e-05, 
    3.715369e-05, 3.709817e-05, 3.73048e-05, 3.724609e-05, 3.741543e-05, 
    3.737291e-05, 3.741347e-05, 3.740115e-05, 3.741363e-05, 3.735125e-05, 
    3.737799e-05, 3.732301e-05, 3.710861e-05, 3.717175e-05, 3.698336e-05, 
    3.687093e-05, 3.679575e-05, 3.674249e-05, 3.675003e-05, 3.676442e-05, 
    3.683811e-05, 3.690716e-05, 3.695979e-05, 3.699519e-05, 3.703012e-05, 
    3.713624e-05, 3.719193e-05, 3.731676e-05, 3.729408e-05, 3.733236e-05, 
    3.736867e-05, 3.742982e-05, 3.741973e-05, 3.74467e-05, 3.733123e-05, 
    3.740805e-05, 3.72812e-05, 3.731594e-05, 3.704027e-05, 3.693441e-05, 
    3.689016e-05, 3.685091e-05, 3.675583e-05, 3.682154e-05, 3.679566e-05, 
    3.685708e-05, 3.689617e-05, 3.687681e-05, 3.699616e-05, 3.69497e-05, 
    3.719523e-05, 3.708949e-05, 3.736444e-05, 3.729872e-05, 3.738016e-05, 
    3.733858e-05, 3.740986e-05, 3.734571e-05, 3.745668e-05, 3.748089e-05, 
    3.746436e-05, 3.752761e-05, 3.734217e-05, 3.741353e-05, 3.68763e-05, 
    3.687946e-05, 3.689411e-05, 3.68297e-05, 3.682572e-05, 3.676644e-05, 
    3.681913e-05, 3.684161e-05, 3.689839e-05, 3.693207e-05, 3.696403e-05, 
    3.703474e-05, 3.71138e-05, 3.722402e-05, 3.730299e-05, 3.735591e-05, 
    3.732342e-05, 3.735211e-05, 3.732006e-05, 3.730501e-05, 3.747186e-05, 
    3.737828e-05, 3.751852e-05, 3.751074e-05, 3.744736e-05, 3.751162e-05, 
    3.688167e-05, 3.68635e-05, 3.680057e-05, 3.684982e-05, 3.675997e-05, 
    3.681036e-05, 3.683936e-05, 3.695081e-05, 3.697513e-05, 3.699804e-05, 
    3.704312e-05, 3.710101e-05, 3.720249e-05, 3.729056e-05, 3.737076e-05, 
    3.736488e-05, 3.736695e-05, 3.738492e-05, 3.734049e-05, 3.739221e-05, 
    3.740095e-05, 3.737819e-05, 3.75097e-05, 3.747215e-05, 3.751058e-05, 
    3.748611e-05, 3.686939e-05, 3.689994e-05, 3.688344e-05, 3.691449e-05, 
    3.689267e-05, 3.698997e-05, 3.701931e-05, 3.715624e-05, 3.709991e-05, 
    3.718936e-05, 3.710895e-05, 3.712324e-05, 3.719255e-05, 3.711326e-05, 
    3.728584e-05, 3.716912e-05, 3.738562e-05, 3.726951e-05, 3.73929e-05, 
    3.737041e-05, 3.740758e-05, 3.744092e-05, 3.748272e-05, 3.755996e-05, 
    3.754205e-05, 3.760649e-05, 3.694539e-05, 3.698512e-05, 3.698148e-05, 
    3.702318e-05, 3.705403e-05, 3.71207e-05, 3.722763e-05, 3.71874e-05, 
    3.72611e-05, 3.727594e-05, 3.716388e-05, 3.723282e-05, 3.701175e-05, 
    3.704764e-05, 3.702618e-05, 3.694859e-05, 3.719684e-05, 3.706952e-05, 
    3.730432e-05, 3.723546e-05, 3.743618e-05, 3.733657e-05, 3.753222e-05, 
    3.7616e-05, 3.769417e-05, 3.778605e-05, 3.700678e-05, 3.697966e-05, 
    3.70281e-05, 3.70953e-05, 3.715724e-05, 3.723969e-05, 3.724805e-05, 
    3.726352e-05, 3.730342e-05, 3.733701e-05, 3.726853e-05, 3.734542e-05, 
    3.705621e-05, 3.720782e-05, 3.696954e-05, 3.704153e-05, 3.709128e-05, 
    3.706934e-05, 3.718277e-05, 3.720952e-05, 3.731816e-05, 3.726195e-05, 
    3.759544e-05, 3.744814e-05, 3.785551e-05, 3.774203e-05, 3.697023e-05, 
    3.700663e-05, 3.713341e-05, 3.70731e-05, 3.724512e-05, 3.728745e-05, 
    3.732174e-05, 3.736574e-05, 3.73704e-05, 3.739644e-05, 3.735378e-05, 
    3.73947e-05, 3.723986e-05, 3.730908e-05, 3.711878e-05, 3.716522e-05, 
    3.714382e-05, 3.712042e-05, 3.719261e-05, 3.726964e-05, 3.727108e-05, 
    3.72958e-05, 3.736574e-05, 3.724581e-05, 3.76148e-05, 3.738752e-05, 
    3.704633e-05, 3.711666e-05, 3.712645e-05, 3.709927e-05, 3.728322e-05, 
    3.721665e-05, 3.739577e-05, 3.734737e-05, 3.742661e-05, 3.738726e-05, 
    3.738148e-05, 3.733086e-05, 3.729938e-05, 3.721974e-05, 3.715482e-05, 
    3.710319e-05, 3.711518e-05, 3.717187e-05, 3.72743e-05, 3.737091e-05, 
    3.734979e-05, 3.742058e-05, 3.723267e-05, 3.731164e-05, 3.728119e-05, 
    3.736051e-05, 3.718637e-05, 3.733529e-05, 3.714833e-05, 3.71647e-05, 
    3.721532e-05, 3.731712e-05, 3.733933e-05, 3.736339e-05, 3.73485e-05, 
    3.727686e-05, 3.726503e-05, 3.721405e-05, 3.720006e-05, 3.716112e-05, 
    3.712896e-05, 3.715839e-05, 3.718933e-05, 3.727681e-05, 3.735565e-05, 
    3.744143e-05, 3.746232e-05, 3.756286e-05, 3.74813e-05, 3.76161e-05, 
    3.750193e-05, 3.769922e-05, 3.734362e-05, 3.749817e-05, 3.721756e-05, 
    3.72478e-05, 3.730268e-05, 3.742793e-05, 3.736013e-05, 3.743932e-05, 
    3.726455e-05, 3.717393e-05, 3.715022e-05, 3.710636e-05, 3.715122e-05, 
    3.714756e-05, 3.719048e-05, 3.717668e-05, 3.727971e-05, 3.722437e-05, 
    3.738139e-05, 3.743864e-05, 3.759981e-05, 3.769853e-05, 3.779852e-05, 
    3.784272e-05, 3.785615e-05, 3.786177e-05,
  8.752311e-10, 8.779569e-10, 8.774257e-10, 8.796268e-10, 8.784038e-10, 
    8.798465e-10, 8.757814e-10, 8.780671e-10, 8.766067e-10, 8.754733e-10, 
    8.839304e-10, 8.797243e-10, 8.882894e-10, 8.856031e-10, 8.923423e-10, 
    8.878745e-10, 8.932601e-10, 8.922079e-10, 8.953919e-10, 8.944751e-10, 
    8.985777e-10, 8.958149e-10, 9.006945e-10, 8.97915e-10, 8.98352e-10, 
    8.957247e-10, 8.805604e-10, 8.834068e-10, 8.803943e-10, 8.807968e-10, 
    8.80615e-10, 8.78431e-10, 8.773337e-10, 8.750191e-10, 8.754384e-10, 
    8.771364e-10, 8.809777e-10, 8.796704e-10, 8.82972e-10, 8.828969e-10, 
    8.86591e-10, 8.849257e-10, 8.911282e-10, 8.893646e-10, 8.945133e-10, 
    8.931923e-10, 8.944522e-10, 8.940695e-10, 8.944572e-10, 8.925245e-10, 
    8.9335e-10, 8.916758e-10, 8.852387e-10, 8.871328e-10, 8.814854e-10, 
    8.781257e-10, 8.758826e-10, 8.742946e-10, 8.745192e-10, 8.749482e-10, 
    8.771464e-10, 8.792082e-10, 8.807807e-10, 8.818399e-10, 8.828862e-10, 
    8.860669e-10, 8.877379e-10, 8.914874e-10, 8.908063e-10, 8.919565e-10, 
    8.930606e-10, 8.949603e-10, 8.94647e-10, 8.954849e-10, 8.919228e-10, 
    8.942838e-10, 8.904193e-10, 8.914632e-10, 8.83189e-10, 8.800222e-10, 
    8.786998e-10, 8.775285e-10, 8.746921e-10, 8.76652e-10, 8.758798e-10, 
    8.777128e-10, 8.7888e-10, 8.78302e-10, 8.818689e-10, 8.804789e-10, 
    8.878371e-10, 8.846653e-10, 8.929291e-10, 8.909457e-10, 8.934174e-10, 
    8.921439e-10, 8.943398e-10, 8.923581e-10, 8.957953e-10, 8.965479e-10, 
    8.96034e-10, 8.980017e-10, 8.922517e-10, 8.94454e-10, 8.782866e-10, 
    8.78381e-10, 8.788186e-10, 8.768953e-10, 8.767767e-10, 8.750085e-10, 
    8.765802e-10, 8.772509e-10, 8.789462e-10, 8.799522e-10, 8.809072e-10, 
    8.830245e-10, 8.853942e-10, 8.887017e-10, 8.91074e-10, 8.926646e-10, 
    8.916881e-10, 8.925504e-10, 8.915871e-10, 8.911348e-10, 8.962672e-10, 
    8.933588e-10, 8.977187e-10, 8.974769e-10, 8.955056e-10, 8.975041e-10, 
    8.78447e-10, 8.779045e-10, 8.760264e-10, 8.774961e-10, 8.748157e-10, 
    8.763185e-10, 8.771837e-10, 8.805117e-10, 8.812391e-10, 8.819253e-10, 
    8.832758e-10, 8.850111e-10, 8.880554e-10, 8.907004e-10, 8.931255e-10, 
    8.929427e-10, 8.930072e-10, 8.935653e-10, 8.922011e-10, 8.937917e-10, 
    8.94063e-10, 8.933563e-10, 8.974446e-10, 8.962766e-10, 8.974718e-10, 
    8.967108e-10, 8.780803e-10, 8.789924e-10, 8.784999e-10, 8.79427e-10, 
    8.787752e-10, 8.816832e-10, 8.825618e-10, 8.866671e-10, 8.849779e-10, 
    8.876611e-10, 8.852491e-10, 8.856776e-10, 8.877563e-10, 8.853782e-10, 
    8.905581e-10, 8.870535e-10, 8.93587e-10, 8.900674e-10, 8.938133e-10, 
    8.931147e-10, 8.942694e-10, 8.953054e-10, 8.966051e-10, 8.990082e-10, 
    8.98451e-10, 9.004572e-10, 8.803502e-10, 8.815381e-10, 8.814294e-10, 
    8.826784e-10, 8.836027e-10, 8.856014e-10, 8.888102e-10, 8.876026e-10, 
    8.898156e-10, 8.90261e-10, 8.868968e-10, 8.889658e-10, 8.823358e-10, 
    8.834109e-10, 8.827682e-10, 8.804455e-10, 8.878857e-10, 8.840667e-10, 
    8.911138e-10, 8.890453e-10, 8.951582e-10, 8.920828e-10, 8.981451e-10, 
    9.007528e-10, 9.031897e-10, 9.060555e-10, 8.82187e-10, 8.813749e-10, 
    8.828259e-10, 8.848394e-10, 8.866973e-10, 8.891722e-10, 8.894235e-10, 
    8.898881e-10, 8.910869e-10, 8.920965e-10, 8.900383e-10, 8.923493e-10, 
    8.836671e-10, 8.882155e-10, 8.810719e-10, 8.832277e-10, 8.847191e-10, 
    8.840614e-10, 8.874637e-10, 8.882666e-10, 8.915296e-10, 8.89841e-10, 
    9.001124e-10, 8.955292e-10, 9.082248e-10, 9.046818e-10, 8.810926e-10, 
    8.821825e-10, 8.859823e-10, 8.841741e-10, 8.893355e-10, 8.90607e-10, 
    8.916375e-10, 8.929693e-10, 8.931142e-10, 8.939229e-10, 8.926006e-10, 
    8.938693e-10, 8.891775e-10, 8.912571e-10, 8.85544e-10, 8.86937e-10, 
    8.86295e-10, 8.855933e-10, 8.877591e-10, 8.900716e-10, 8.901154e-10, 
    8.908577e-10, 8.929677e-10, 8.893563e-10, 9.007143e-10, 8.936444e-10, 
    8.83372e-10, 8.854797e-10, 8.85774e-10, 8.849588e-10, 8.904798e-10, 
    8.884805e-10, 8.939024e-10, 8.92408e-10, 8.948606e-10, 8.93638e-10, 
    8.934584e-10, 8.919117e-10, 8.909655e-10, 8.885732e-10, 8.866247e-10, 
    8.850763e-10, 8.854359e-10, 8.871365e-10, 8.902116e-10, 8.931299e-10, 
    8.924803e-10, 8.946735e-10, 8.889616e-10, 8.913336e-10, 8.904187e-10, 
    8.928071e-10, 8.875717e-10, 8.920436e-10, 8.864303e-10, 8.869214e-10, 
    8.884407e-10, 8.914983e-10, 8.921662e-10, 8.928963e-10, 8.92442e-10, 
    8.902887e-10, 8.899333e-10, 8.884025e-10, 8.879825e-10, 8.868141e-10, 
    8.858492e-10, 8.867321e-10, 8.876604e-10, 8.902873e-10, 8.926567e-10, 
    8.95321e-10, 8.959709e-10, 8.990975e-10, 8.965602e-10, 9.007547e-10, 
    8.972004e-10, 9.03346e-10, 8.922943e-10, 8.970845e-10, 8.88508e-10, 
    8.89416e-10, 8.910641e-10, 8.949012e-10, 8.927953e-10, 8.952553e-10, 
    8.89919e-10, 8.87198e-10, 8.864869e-10, 8.851715e-10, 8.86517e-10, 
    8.864073e-10, 8.87695e-10, 8.872809e-10, 8.903744e-10, 8.887126e-10, 
    8.934554e-10, 8.952344e-10, 9.00249e-10, 9.03325e-10, 9.064454e-10, 
    9.078255e-10, 9.08245e-10, 9.084207e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  0.5836036, 0.5527475, 0.5587046, 0.53412, 0.5477114, 0.5316789, 0.5773047, 
    0.5515357, 0.5679432, 0.5808014, 0.4875063, 0.5330309, 0.4415244, 
    0.4692921, 0.4009403, 0.4458025, 0.3921618, 0.4021982, 0.3723571, 
    0.3807883, 0.3439219, 0.3684985, 0.3256117, 0.3497048, 0.3458737, 
    0.3693256, 0.5237485, 0.4930955, 0.5255864, 0.5211697, 0.5231484, 
    0.5474318, 0.5598079, 0.5859776, 0.5811993, 0.5619881, 0.5191876, 
    0.533587, 0.4975506, 0.4983542, 0.4589748, 0.4763948, 0.412854, 
    0.4305114, 0.3804343, 0.3927497, 0.3810094, 0.3845499, 0.3809634, 
    0.3991033, 0.3912807, 0.407426, 0.4731137, 0.4533758, 0.5136296, 
    0.5509421, 0.5761682, 0.5942749, 0.5917056, 0.5868175, 0.5618765, 
    0.5387259, 0.5213004, 0.5097556, 0.49847, 0.4645503, 0.4471767, 
    0.4093275, 0.4160416, 0.4046938, 0.3939853, 0.3763298, 0.3792072, 
    0.3715297, 0.4049879, 0.3825931, 0.4198897, 0.4095256, 0.4954389, 
    0.5296882, 0.5445014, 0.5575588, 0.5897326, 0.5674577, 0.5762094, 
    0.5554507, 0.5423869, 0.5488348, 0.5094411, 0.5246388, 0.4461556, 
    0.4791774, 0.3952271, 0.4146591, 0.3906353, 0.4028077, 0.3820646, 
    0.4007092, 0.3686915, 0.3619021, 0.366535, 0.3489045, 0.401756, 
    0.3810112, 0.5490169, 0.5479636, 0.5430627, 0.5647097, 0.5660411, 
    0.5861099, 0.5682405, 0.560683, 0.541631, 0.5304666, 0.5199248, 
    0.4970092, 0.4715084, 0.4372858, 0.4133863, 0.3977137, 0.4072888, 
    0.3988298, 0.4082922, 0.4127624, 0.3644394, 0.3912092, 0.3514114, 
    0.3535543, 0.3713488, 0.3533124, 0.547224, 0.553292, 0.5745265, 
    0.5578877, 0.5883073, 0.5712236, 0.56147, 0.5243242, 0.516272, 0.5088512, 
    0.4943042, 0.475497, 0.4438801, 0.4171253, 0.3933657, 0.3950836, 
    0.3944786, 0.3892571, 0.4022555, 0.3871429, 0.3846362, 0.3912102, 
    0.3538419, 0.3643184, 0.3535999, 0.3603998, 0.5513167, 0.5411296, 
    0.5466271, 0.5363056, 0.5435722, 0.5115204, 0.5020435, 0.458238, 
    0.475858, 0.4479384, 0.4729892, 0.4685113, 0.4470479, 0.4716201, 
    0.4185848, 0.4542569, 0.3890548, 0.4235451, 0.3869408, 0.3934671, 
    0.3826893, 0.373166, 0.361358, 0.3401091, 0.3449659, 0.3276046, 
    0.5260569, 0.513065, 0.5142003, 0.5007142, 0.4908258, 0.4692824, 
    0.4361562, 0.4484926, 0.4259561, 0.4214951, 0.4557735, 0.4345924, 
    0.5044313, 0.492931, 0.4997635, 0.5250304, 0.4456419, 0.4859323, 
    0.4129971, 0.4337573, 0.3745168, 0.4034647, 0.3476566, 0.3251646, 
    0.3047841, 0.2820172, 0.5060185, 0.5147917, 0.499118, 0.4773613, 
    0.4578665, 0.4324787, 0.4299144, 0.4252416, 0.4132407, 0.4032754, 
    0.4237725, 0.400795, 0.4902859, 0.4422432, 0.5181263, 0.4949015, 
    0.4786083, 0.4859391, 0.4499109, 0.441675, 0.4088996, 0.4256988, 
    0.3306386, 0.371175, 0.265451, 0.2928063, 0.5178706, 0.5060468, 
    0.4653383, 0.4847353, 0.4308042, 0.4180388, 0.4077876, 0.3948643, 
    0.3934784, 0.3859292, 0.3983378, 0.3864143, 0.4324253, 0.4115642, 
    0.4698736, 0.4553812, 0.462024, 0.4693583, 0.4468758, 0.423447, 
    0.4229467, 0.4155583, 0.3950754, 0.4305926, 0.3256068, 0.3886994, 
    0.4932668, 0.4706363, 0.4674858, 0.4760303, 0.4193109, 0.4395082, 
    0.3861115, 0.400221, 0.3772328, 0.3885725, 0.3902552, 0.4050917, 
    0.4144633, 0.4385741, 0.4586265, 0.4747865, 0.4710084, 0.4533272, 
    0.4220307, 0.3933555, 0.3995559, 0.378956, 0.4345979, 0.4108327, 
    0.4199482, 0.3963759, 0.4488238, 0.4039889, 0.4606142, 0.4555201, 
    0.4399133, 0.4092468, 0.4025913, 0.3955526, 0.3998876, 0.421248, 
    0.4247937, 0.4402884, 0.444612, 0.4566267, 0.4666768, 0.4574924, 
    0.4479297, 0.4212365, 0.3978226, 0.3730322, 0.3670866, 0.3394244, 
    0.3618614, 0.3252737, 0.3562539, 0.3036537, 0.4014488, 0.3571778, 
    0.4392066, 0.4299852, 0.4135347, 0.3769389, 0.3964851, 0.3736725, 
    0.4249324, 0.4527252, 0.46003, 0.4737988, 0.4597172, 0.4608558, 
    0.4475311, 0.4517949, 0.4203626, 0.4371235, 0.390299, 0.3738486, 
    0.3294018, 0.3037378, 0.278929, 0.2684214, 0.2652779, 0.2639718,
  0.9312378, 0.9125337, 0.9161377, 0.9012924, 0.9094925, 0.8998227, 
    0.9274133, 0.9117996, 0.9217339, 0.9295377, 0.8733478, 0.900637, 
    0.8114799, 0.8239906, 0.7934842, 0.8133957, 0.7896399, 0.794039, 
    0.7810352, 0.7846878, 0.7688482, 0.7793695, 0.761126, 0.7713102, 
    0.7696786, 0.779726, 0.8950546, 0.8766815, 0.8961593, 0.8935034, 
    0.8946939, 0.9093221, 0.9168011, 0.9326841, 0.9297795, 0.918124, 
    0.8923125, 0.9009746, 0.8793552, 0.8798355, 0.8193254, 0.8272153, 
    0.7987326, 0.8065652, 0.7845341, 0.789899, 0.7847834, 0.786323, 
    0.7847634, 0.7926804, 0.7892567, 0.7963389, 0.8257242, 0.8168017, 
    0.8889784, 0.9114366, 0.9267224, 0.9377323, 0.936168, 0.9331928, 
    0.9180562, 0.9040711, 0.893585, 0.8866581, 0.8799046, 0.8218389, 
    0.8140136, 0.797175, 0.800142, 0.7951349, 0.7904393, 0.7827534, 
    0.7840012, 0.7806767, 0.7952659, 0.7854705, 0.8018464, 0.7972642, 
    0.8780798, 0.8986273, 0.907548, 0.9154437, 0.9349669, 0.9214379, 
    0.9267468, 0.9141707, 0.9062788, 0.9101722, 0.8864697, 0.8955904, 
    0.8135555, 0.8284793, 0.7909825, 0.7995304, 0.7889755, 0.7943076, 
    0.7852412, 0.7933859, 0.7794521, 0.7765291, 0.7785223, 0.7709706, 
    0.7938454, 0.7847834, 0.9102815, 0.9096451, 0.9066871, 0.9197723, 
    0.9205797, 0.9327638, 0.9219142, 0.9173346, 0.9058239, 0.8990956, 
    0.8927576, 0.8790303, 0.8249944, 0.8095855, 0.798968, 0.7920721, 
    0.7962791, 0.7925614, 0.7967209, 0.7986932, 0.7776196, 0.789225, 
    0.7720393, 0.7729544, 0.7805983, 0.772851, 0.9091985, 0.9128658, 
    0.9257265, 0.915645, 0.9341006, 0.923722, 0.9178092, 0.8953983, 
    0.8905656, 0.886115, 0.8774155, 0.8268072, 0.8125368, 0.8006204, 
    0.7901688, 0.7909204, 0.7906556, 0.7883737, 0.7940646, 0.7874519, 
    0.7863594, 0.7892264, 0.7730773, 0.7775691, 0.7729739, 0.7758857, 
    0.9116719, 0.9055206, 0.9088384, 0.9026114, 0.9069929, 0.8877115, 
    0.8820357, 0.8189907, 0.8269707, 0.8143569, 0.8256683, 0.8236368, 
    0.8139532, 0.8250476, 0.8012648, 0.8171955, 0.7882854, 0.8034623, 
    0.7873638, 0.7902131, 0.7855139, 0.7813841, 0.7762967, 0.7672337, 
    0.7692943, 0.7619628, 0.8964432, 0.8886393, 0.8893231, 0.8812457, 
    0.8753385, 0.8239874, 0.809082, 0.8146078, 0.8045386, 0.8025573, 
    0.8178834, 0.808383, 0.8834675, 0.8765911, 0.8806762, 0.8958243, 
    0.8133258, 0.8724176, 0.7987958, 0.8080117, 0.7819683, 0.7945939, 
    0.7704386, 0.7609368, 0.7524727, 0.7431926, 0.8844188, 0.8896779, 
    0.880292, 0.8276522, 0.8188257, 0.8074411, 0.8062994, 0.8042204, 
    0.7989044, 0.794513, 0.8035661, 0.7934237, 0.8750069, 0.8118033, 
    0.8916769, 0.8777669, 0.8282204, 0.8724248, 0.8152455, 0.8115509, 
    0.7969869, 0.8044243, 0.763234, 0.7805214, 0.7365851, 0.7475638, 
    0.8915253, 0.884437, 0.8221996, 0.8717081, 0.8066958, 0.8010255, 
    0.7964989, 0.790823, 0.7902178, 0.7869227, 0.7923457, 0.7871346, 
    0.8074173, 0.7981636, 0.8242559, 0.8177056, 0.8207035, 0.8240222, 
    0.8138822, 0.8034213, 0.8032018, 0.7999271, 0.790907, 0.8066015, 
    0.7611173, 0.7881225, 0.8767966, 0.8245977, 0.8231731, 0.8270503, 
    0.8015889, 0.8105804, 0.7870025, 0.7931716, 0.7831452, 0.7880753, 
    0.7888094, 0.7953117, 0.7994439, 0.8101622, 0.8191683, 0.8264854, 
    0.8247704, 0.8167801, 0.8027931, 0.790163, 0.792878, 0.7838925, 
    0.8083872, 0.7978396, 0.8018701, 0.7914855, 0.8147559, 0.7948184, 
    0.8200669, 0.8177691, 0.8107616, 0.7971383, 0.7942125, 0.7911243, 
    0.7930254, 0.8024465, 0.8040211, 0.8109302, 0.8128656, 0.8182681, 
    0.8228077, 0.8186576, 0.8143536, 0.8024424, 0.7921184, 0.7813258, 
    0.7787607, 0.76694, 0.7765087, 0.7609774, 0.7740989, 0.7520016, 
    0.7937057, 0.7744992, 0.8104464, 0.8063312, 0.7990313, 0.7830145, 
    0.7915334, 0.7816011, 0.804083, 0.8165078, 0.8198029, 0.8260362, 
    0.8196617, 0.8201758, 0.8141766, 0.8160926, 0.8020551, 0.8095152, 
    0.7888278, 0.781678, 0.7627168, 0.7520397, 0.7419535, 0.7377611, 
    0.7365175, 0.7360022,
  1.172322, 1.173099, 1.172974, 1.173412, 1.173196, 1.173443, 1.172505, 
    1.173123, 1.172755, 1.172405, 1.173604, 1.173426, 1.212348, 1.218197, 
    1.203276, 1.213266, 1.20122, 1.20357, 1.196442, 1.198501, 1.189195, 
    1.195487, 1.184258, 1.19071, 1.189709, 1.195692, 1.17353, 1.173629, 
    1.173512, 1.173553, 1.173536, 1.173201, 1.172949, 1.172249, 1.172393, 
    1.172899, 1.173569, 1.173419, 1.17364, 1.173641, 1.216056, 1.219652, 
    1.206012, 1.209955, 1.198416, 1.20136, 1.198555, 1.199408, 1.198543, 
    1.20285, 1.201012, 1.204775, 1.218982, 1.214878, 1.173606, 1.173135, 
    1.172537, 1.171983, 1.172067, 1.172223, 1.172902, 1.173346, 1.173552, 
    1.173624, 1.173641, 1.217214, 1.213561, 1.205208, 1.206734, 1.204145, 
    1.201652, 1.197416, 1.198118, 1.196237, 1.204214, 1.198936, 1.2076, 
    1.205255, 1.173635, 1.173468, 1.173253, 1.172999, 1.172131, 1.172767, 
    1.172536, 1.173044, 1.173289, 1.173175, 1.173625, 1.173522, 1.213343, 
    1.220216, 1.201944, 1.206422, 1.20086, 1.203711, 1.198809, 1.203225, 
    1.195534, 1.193833, 1.194996, 1.190503, 1.203467, 1.198554, 1.173172, 
    1.173191, 1.173277, 1.172835, 1.172802, 1.172245, 1.172748, 1.172929, 
    1.173301, 1.173458, 1.173564, 1.173639, 1.218652, 1.211433, 1.206133, 
    1.202527, 1.204744, 1.202787, 1.204973, 1.205993, 1.194471, 1.200995, 
    1.191153, 1.191706, 1.196192, 1.191644, 1.173205, 1.173088, 1.172582, 
    1.172992, 1.172176, 1.172671, 1.172911, 1.173525, 1.17359, 1.173627, 
    1.173634, 1.219469, 1.212856, 1.206977, 1.201506, 1.20191, 1.201768, 
    1.200533, 1.203583, 1.200029, 1.199428, 1.200996, 1.19178, 1.194442, 
    1.191718, 1.193454, 1.173128, 1.173309, 1.173216, 1.173382, 1.173269, 
    1.173616, 1.173641, 1.2159, 1.219542, 1.213724, 1.218956, 1.218036, 
    1.213531, 1.218676, 1.207304, 1.215062, 1.200485, 1.208411, 1.199981, 
    1.20153, 1.198961, 1.19664, 1.193696, 1.188188, 1.189472, 1.184808, 
    1.173508, 1.173609, 1.173603, 1.173642, 1.173622, 1.218196, 1.211188, 
    1.213844, 1.20895, 1.207958, 1.215385, 1.210847, 1.173639, 1.173629, 
    1.173642, 1.173518, 1.213233, 1.173595, 1.206045, 1.210666, 1.196972, 
    1.203861, 1.190177, 1.184133, 1.178337, 1.171424, 1.173635, 1.173599, 
    1.173642, 1.219846, 1.215824, 1.210386, 1.209824, 1.208791, 1.206101, 
    1.203819, 1.208464, 1.203245, 1.173619, 1.212505, 1.173577, 1.173635, 
    1.2201, 1.173596, 1.214146, 1.212384, 1.205111, 1.208893, 1.185635, 
    1.196147, 1.166061, 1.174761, 1.173579, 1.173636, 1.21738, 1.173588, 
    1.210019, 1.207183, 1.204858, 1.201858, 1.201532, 1.199738, 1.202672, 
    1.199855, 1.210374, 1.20572, 1.218318, 1.215302, 1.216693, 1.218212, 
    1.213499, 1.208391, 1.208282, 1.206624, 1.2019, 1.209973, 1.18425, 
    1.200393, 1.173631, 1.218472, 1.217825, 1.219578, 1.207469, 1.211915, 
    1.199782, 1.203111, 1.197637, 1.20037, 1.20077, 1.204238, 1.206377, 
    1.211713, 1.215983, 1.219324, 1.218551, 1.214868, 1.208076, 1.201502, 
    1.202955, 1.198057, 1.210849, 1.205552, 1.207611, 1.202213, 1.213914, 
    1.203977, 1.216399, 1.215332, 1.212003, 1.205189, 1.203661, 1.202019, 
    1.203034, 1.207902, 1.208692, 1.212084, 1.213014, 1.215564, 1.217659, 
    1.215746, 1.213723, 1.2079, 1.202551, 1.196607, 1.195135, 1.188002, 
    1.19382, 1.184157, 1.19239, 1.177999, 1.203392, 1.19263, 1.211851, 
    1.20984, 1.206165, 1.197563, 1.202239, 1.196763, 1.208723, 1.21474, 
    1.216277, 1.219122, 1.216212, 1.21645, 1.213639, 1.214545, 1.207705, 
    1.211399, 1.20078, 1.196807, 1.1853, 1.178028, 1.17045, 1.167047, 
    1.166004, 1.165567,
  0.506425, 0.4962071, 0.4981915, 0.4899662, 0.4945269, 0.4891443, 0.5043516, 
    0.4958016, 0.5012577, 0.5055046, 0.4740624, 0.4895999, 0.4580597, 
    0.467906, 0.4432479, 0.4595888, 0.4399673, 0.4437187, 0.4324504, 
    0.4356725, 0.4213253, 0.430965, 0.4139324, 0.4236236, 0.4221037, 
    0.4312837, 0.4864678, 0.4759921, 0.4870893, 0.4855931, 0.4862646, 
    0.4944323, 0.4985551, 0.5072078, 0.5056357, 0.4992816, 0.4849205, 
    0.4897892, 0.4775355, 0.4778117, 0.4642733, 0.4703923, 0.4476575, 
    0.4540981, 0.4355379, 0.4401907, 0.435756, 0.4370999, 0.4357385, 
    0.4425665, 0.4396383, 0.4456567, 0.469245, 0.4622892, 0.4830327, 
    0.4956004, 0.503976, 0.5099301, 0.5090877, 0.5074824, 0.4992444, 
    0.491517, 0.4856397, 0.4817142, 0.4778514, 0.4662341, 0.4600809, 
    0.4463569, 0.4488286, 0.4446436, 0.4406542, 0.4339717, 0.4350703, 
    0.4321312, 0.4447546, 0.4363563, 0.4502375, 0.4464321, 0.4767985, 
    0.4884752, 0.4934482, 0.4978098, 0.5084402, 0.5010957, 0.5039892, 
    0.4971098, 0.492745, 0.4949032, 0.4816069, 0.4867695, 0.4597166, 
    0.4713609, 0.4411191, 0.4483211, 0.4393965, 0.4439462, 0.4361562, 
    0.4431659, 0.4310387, 0.4284072, 0.430205, 0.423309, 0.443555, 0.4357557, 
    0.4949635, 0.4946114, 0.4929719, 0.5001846, 0.5006265, 0.5072508, 
    0.5013562, 0.4988487, 0.4924924, 0.4887376, 0.4851725, 0.4773483, 
    0.4686816, 0.4565395, 0.4478535, 0.4420493, 0.4456068, 0.4424657, 
    0.4459773, 0.4476252, 0.4293925, 0.4396109, 0.4242993, 0.4251436, 
    0.4320612, 0.4250485, 0.4943643, 0.4963908, 0.5034345, 0.497921, 
    0.5079729, 0.5023425, 0.4991087, 0.4866607, 0.483933, 0.4814046, 
    0.4764181, 0.4700787, 0.4589052, 0.4492242, 0.4404224, 0.4410662, 
    0.4408395, 0.4388773, 0.4437405, 0.43808, 0.4371311, 0.4396125, 
    0.4252567, 0.4293476, 0.4251616, 0.4278242, 0.495732, 0.4923236, 
    0.4941649, 0.4907031, 0.4931413, 0.4823126, 0.4790732, 0.4640101, 
    0.4702042, 0.4603541, 0.4692023, 0.467632, 0.4600319, 0.4687236, 
    0.4497563, 0.4625986, 0.4388011, 0.4515637, 0.4380037, 0.4404604, 
    0.4363948, 0.43276, 0.428197, 0.4198047, 0.4217449, 0.4147488, 0.4872492, 
    0.4828401, 0.4832287, 0.4786212, 0.4752181, 0.467904, 0.4561343, 
    0.4605541, 0.4524469, 0.4508224, 0.4631418, 0.4555699, 0.4798933, 
    0.4759414, 0.4782942, 0.4869007, 0.4595339, 0.4735239, 0.4477101, 
    0.4552702, 0.4332777, 0.444187, 0.4228136, 0.4137463, 0.4052582, 
    0.3953901, 0.4804372, 0.48343, 0.478074, 0.4707267, 0.4638816, 0.4548083, 
    0.4538822, 0.4521865, 0.4478009, 0.4441197, 0.45165, 0.4431979, 
    0.4750243, 0.4583192, 0.4845616, 0.4766198, 0.4711626, 0.4735287, 
    0.4610599, 0.4581179, 0.4461995, 0.4523535, 0.4159794, 0.4319921, 
    0.3879206, 0.4001195, 0.4844761, 0.4804478, 0.4665163, 0.473112, 
    0.4542041, 0.4495595, 0.4457912, 0.4409824, 0.4404643, 0.4376209, 
    0.4422823, 0.4378051, 0.454789, 0.4471835, 0.4681119, 0.4630016, 
    0.4653515, 0.4679311, 0.4599778, 0.4515311, 0.451352, 0.4486499, 
    0.4410508, 0.4541276, 0.4139207, 0.4386571, 0.4760611, 0.4683748, 
    0.4672728, 0.4702658, 0.4500247, 0.4573398, 0.4376903, 0.4429842, 
    0.4343175, 0.4386196, 0.4392532, 0.4447933, 0.4482493, 0.4570037, 
    0.4641501, 0.4698317, 0.4685096, 0.4622723, 0.4510156, 0.4404169, 
    0.4427342, 0.4349749, 0.4555739, 0.4469127, 0.4502561, 0.4415489, 
    0.4606714, 0.4443741, 0.4648541, 0.4630519, 0.4574852, 0.4463257, 
    0.4438657, 0.44124, 0.4428601, 0.4507307, 0.4520233, 0.4576206, 
    0.4591678, 0.4634443, 0.4669897, 0.4637499, 0.4603517, 0.4507279, 
    0.4420882, 0.4327081, 0.4304195, 0.4195248, 0.4283874, 0.4137837, 
    0.42619, 0.4047697, 0.4434349, 0.4265583, 0.4572326, 0.453908, 0.4479053, 
    0.4342009, 0.4415898, 0.4329516, 0.452074, 0.4620568, 0.4646476, 
    0.4694857, 0.4645371, 0.4649393, 0.4602118, 0.4617301, 0.450409, 
    0.4564837, 0.4392689, 0.43302, 0.4154803, 0.4048107, 0.3940219, 0.389282, 
    0.3878424, 0.387241,
  0.04991171, 0.04802241, 0.04838632, 0.04688735, 0.04771542, 0.04673892, 
    0.04952523, 0.04794823, 0.04895147, 0.04973995, 0.04405922, 0.04682116, 
    0.04129905, 0.04298105, 0.03883456, 0.04155796, 0.03829936, 0.03891169, 
    0.03708753, 0.0376045, 0.03533095, 0.03685046, 0.03418794, 0.03569023, 
    0.03545243, 0.03690125, 0.04625731, 0.04439746, 0.04636891, 0.04610048, 
    0.04622085, 0.04769816, 0.04845315, 0.05005804, 0.04976439, 0.04858683, 
    0.04598008, 0.04685536, 0.04466896, 0.04471764, 0.04235642, 0.04341131, 
    0.03956003, 0.04063216, 0.03758284, 0.03833568, 0.03761796, 0.03783472, 
    0.03761515, 0.03872309, 0.03824591, 0.03923, 0.0432125, 0.04201725, 
    0.04564302, 0.04791144, 0.04945539, 0.05056867, 0.05041038, 0.05010942, 
    0.04857999, 0.04716805, 0.04610883, 0.04540839, 0.04472464, 0.04269298, 
    0.04164146, 0.03934532, 0.03975386, 0.03906343, 0.0384111, 0.03733116, 
    0.0375076, 0.03703652, 0.03908166, 0.0377147, 0.03998772, 0.03935772, 
    0.04453921, 0.04661828, 0.04751887, 0.04831621, 0.05028887, 0.04892151, 
    0.04945783, 0.04818777, 0.04739096, 0.04778408, 0.04538933, 0.04631147, 
    0.04157964, 0.04357954, 0.03848683, 0.03966981, 0.03820663, 0.03894898, 
    0.03768244, 0.03882113, 0.03686221, 0.03644404, 0.03672946, 0.03564094, 
    0.03888487, 0.03761791, 0.04779509, 0.04773083, 0.04743221, 0.04875328, 
    0.04883484, 0.05006608, 0.04896969, 0.04850715, 0.04734507, 0.04666556, 
    0.04602517, 0.04463599, 0.04311503, 0.04104247, 0.03959244, 0.03863858, 
    0.03922179, 0.03870661, 0.03928278, 0.03955469, 0.03660033, 0.03824144, 
    0.03579622, 0.03592888, 0.03702534, 0.03591391, 0.04768575, 0.04805603, 
    0.04935478, 0.04833663, 0.05020127, 0.04915224, 0.04855501, 0.04629194, 
    0.04580361, 0.0453534, 0.04447232, 0.04335693, 0.0414421, 0.03981946, 
    0.03837338, 0.03847821, 0.03844128, 0.03812239, 0.03891527, 0.03799321, 
    0.03783976, 0.03824171, 0.03594667, 0.0365932, 0.0359317, 0.03635174, 
    0.04793549, 0.04731442, 0.04764941, 0.04702062, 0.04746303, 0.0455148, 
    0.04494032, 0.04231134, 0.04337869, 0.04168785, 0.04320509, 0.04293377, 
    0.04163314, 0.04312228, 0.03990776, 0.04207005, 0.03811003, 0.0402085, 
    0.03798086, 0.03837956, 0.03772091, 0.03713704, 0.03641075, 0.03509426, 
    0.0353964, 0.03431321, 0.04639764, 0.04560872, 0.04567796, 0.04486047, 
    0.04426163, 0.0429807, 0.04097422, 0.04172183, 0.04035588, 0.04008502, 
    0.04216283, 0.04087926, 0.0450854, 0.04438856, 0.04480275, 0.04633504, 
    0.04154865, 0.04396506, 0.03956872, 0.04082888, 0.03721993, 0.03898847, 
    0.0355634, 0.03415943, 0.03287147, 0.03140602, 0.04518174, 0.04571385, 
    0.04476389, 0.04346936, 0.04228934, 0.04075129, 0.04059597, 0.0403124, 
    0.03958374, 0.03897744, 0.04022288, 0.03882638, 0.04422766, 0.04134292, 
    0.0459159, 0.04450776, 0.04354508, 0.04396591, 0.04180784, 0.04130889, 
    0.03931938, 0.04034027, 0.03450249, 0.03701429, 0.03031947, 0.03210407, 
    0.04590063, 0.04518363, 0.04274152, 0.04389313, 0.04064993, 0.03987509, 
    0.03925214, 0.03846455, 0.0383802, 0.03791893, 0.03867663, 0.03794872, 
    0.04074805, 0.03948171, 0.0430166, 0.04213887, 0.04254131, 0.04298538, 
    0.04162396, 0.04020305, 0.04017321, 0.03972425, 0.0384757, 0.04063711, 
    0.03418616, 0.03808669, 0.04440958, 0.043062, 0.04287183, 0.04338938, 
    0.03995235, 0.04117743, 0.03793015, 0.03879139, 0.03738666, 0.03808061, 
    0.03818337, 0.03908802, 0.03965791, 0.04112072, 0.04233532, 0.0433141, 
    0.0430853, 0.04201438, 0.04011717, 0.03837248, 0.03875049, 0.03749227, 
    0.04087992, 0.039437, 0.03999081, 0.03855691, 0.04174177, 0.03901919, 
    0.04245596, 0.04214747, 0.04120198, 0.03934018, 0.03893578, 0.03850654, 
    0.03877109, 0.04006976, 0.04028515, 0.04122485, 0.04148658, 0.04221453, 
    0.04282303, 0.04226681, 0.04168745, 0.04006927, 0.03864493, 0.03712875, 
    0.03676358, 0.0350508, 0.03644091, 0.03416515, 0.03609364, 0.03279811, 
    0.03886519, 0.03615174, 0.04115934, 0.0406003, 0.03960101, 0.03736794, 
    0.03856358, 0.03716771, 0.04029362, 0.04197764, 0.04242054, 0.04325417, 
    0.0424016, 0.04247056, 0.0416637, 0.04192195, 0.04001623, 0.04103307, 
    0.03818591, 0.03717865, 0.03442566, 0.03280426, 0.03120552, 0.03051606, 
    0.03030821, 0.03022159,
  0.001340993, 0.001263546, 0.00127834, 0.00121778, 0.001251111, 0.001211838, 
    0.001325022, 0.001260537, 0.001301433, 0.001333887, 0.001106295, 
    0.001215129, 0.001001077, 0.001064767, 0.000910224, 0.001010793, 
    0.000890889, 0.0009130223, 0.0008476401, 0.0008659997, 0.0007862776, 
    0.000839266, 0.0007477448, 0.0007986988, 0.00079047, 0.0008410577, 
    0.001192627, 0.001119435, 0.00119707, 0.001186395, 0.001191178, 
    0.001250413, 0.001281064, 0.001347057, 0.001334897, 0.001286517, 
    0.001181617, 0.001216499, 0.00113002, 0.001131922, 0.001040958, 
    0.001081274, 0.0009366599, 0.0009762007, 0.0008652276, 0.0008921967, 
    0.0008664795, 0.0008742188, 0.0008663791, 0.0009061854, 0.0008889658, 
    0.0009246015, 0.001073636, 0.001028107, 0.001168278, 0.001259046, 
    0.001322143, 0.00136829, 0.001361696, 0.001349188, 0.001286238, 
    0.001229044, 0.001186726, 0.001159022, 0.001132195, 0.001053764, 
    0.001013934, 0.000928809, 0.000943767, 0.0009185359, 0.000894914, 
    0.0008562755, 0.0008625481, 0.0008458358, 0.000919199, 0.0008699307, 
    0.000952366, 0.0009292618, 0.001124957, 0.001207016, 0.001243172, 
    0.001275486, 0.001356641, 0.001300205, 0.001322243, 0.001270261, 
    0.001238015, 0.001253888, 0.001158272, 0.001194783, 0.001011608, 
    0.001087752, 0.0008976455, 0.0009406828, 0.0008875536, 0.0009143764, 
    0.0008687791, 0.0009097375, 0.0008396802, 0.0008249769, 0.0008350031, 
    0.0007969906, 0.000912049, 0.0008664777, 0.001254334, 0.001251734, 
    0.001239677, 0.001293319, 0.001296656, 0.00134739, 0.00130218, 
    0.001283266, 0.001236166, 0.001208906, 0.001183405, 0.001128733, 
    0.001069898, 0.0009914809, 0.0009378469, 0.0009031275, 0.0009243022, 
    0.0009055887, 0.0009265263, 0.0009364642, 0.000830462, 0.0008888052, 
    0.000802376, 0.0008069865, 0.0008454406, 0.000806466, 0.001249911, 
    0.00126491, 0.001317999, 0.001276317, 0.001353001, 0.001309671, 
    0.001285218, 0.001194005, 0.001174626, 0.001156857, 0.00112235, 
    0.001079183, 0.001006442, 0.0009461763, 0.0008935548, 0.0008973345, 
    0.0008960023, 0.0008845272, 0.0009131522, 0.000879893, 0.0008743994, 
    0.0008888147, 0.0008076054, 0.0008302113, 0.0008070847, 0.0008217435, 
    0.001260021, 0.001234932, 0.001248443, 0.001223124, 0.001240919, 
    0.001163217, 0.001140634, 0.001039247, 0.001080019, 0.00101568, 
    0.001073351, 0.001062958, 0.00101362, 0.001070176, 0.000949423, 
    0.001030105, 0.0008840834, 0.0009605088, 0.0008794505, 0.0008937775, 
    0.0008701526, 0.0008493924, 0.0008238104, 0.0007781317, 0.0007885354, 
    0.0007514584, 0.001198214, 0.001166923, 0.001169658, 0.001137507, 
    0.001114152, 0.001064753, 0.0009889336, 0.001016959, 0.0009659576, 
    0.0009559516, 0.001033616, 0.0009853932, 0.001146323, 0.001119088, 
    0.001135249, 0.001195721, 0.001010443, 0.001102647, 0.0009369783, 
    0.0009835165, 0.0008523289, 0.000915811, 0.0007943063, 0.0007467762, 
    0.0007034834, 0.0006553394, 0.001150106, 0.001171076, 0.001133729, 
    0.001083508, 0.001038412, 0.0009806288, 0.000974857, 0.000964349, 
    0.0009375282, 0.00091541, 0.00096104, 0.0009099276, 0.001112832, 
    0.001002722, 0.001179073, 0.001123731, 0.001086424, 0.001102679, 
    0.001020201, 0.001001446, 0.000927862, 0.0009653803, 0.000757893, 
    0.0008450501, 0.0006204264, 0.0006781227, 0.001178468, 0.00115018, 
    0.001055615, 0.001099862, 0.0009768608, 0.0009482214, 0.0009254089, 
    0.0008968417, 0.0008938004, 0.0008772321, 0.0009045038, 0.0008782989, 
    0.0009805084, 0.0009337935, 0.001066127, 0.001032709, 0.001047986, 
    0.001064932, 0.001013275, 0.0009603077, 0.0009592058, 0.0009426801, 
    0.0008972438, 0.0009763844, 0.0007476842, 0.0008832457, 0.001119907, 
    0.001067866, 0.00106059, 0.00108043, 0.0009510638, 0.0009965247, 
    0.000877634, 0.0009086594, 0.0008582466, 0.0008830273, 0.0008867177, 
    0.0009194307, 0.0009402464, 0.0009944042, 0.001040157, 0.001077537, 
    0.001068758, 0.001027999, 0.0009571377, 0.0008935224, 0.0009071777, 
    0.0008620024, 0.0009854179, 0.0009321585, 0.0009524798, 0.0009001758, 
    0.00101771, 0.0009169274, 0.00104474, 0.001033035, 0.0009974432, 
    0.0009286212, 0.0009138969, 0.000898357, 0.0009079237, 0.0009553888, 
    0.0009633413, 0.000998299, 0.001008112, 0.001035575, 0.001058726, 
    0.001037557, 0.001015665, 0.0009553712, 0.0009033572, 0.0008490987, 
    0.0008362044, 0.0007766389, 0.0008248671, 0.0007469704, 0.0008127256, 
    0.0007010447, 0.000911335, 0.0008147523, 0.000995848, 0.0009750177, 
    0.0009381608, 0.0008575814, 0.0009004166, 0.0008504786, 0.0009636544, 
    0.00102661, 0.001043394, 0.001075235, 0.001042674, 0.001045295, 
    0.00101477, 0.001024507, 0.0009534164, 0.00099113, 0.0008868088, 
    0.0008508662, 0.0007552789, 0.0007012492, 0.0006488464, 0.0006266931, 
    0.0006200682, 0.0006173145,
  8.818053e-06, 8.041774e-06, 8.188288e-06, 7.594008e-06, 7.919293e-06, 
    7.536487e-06, 8.656107e-06, 8.012084e-06, 8.418671e-06, 8.745881e-06, 
    6.53915e-06, 7.568329e-06, 5.593382e-06, 6.159864e-06, 4.818942e-06, 
    5.678581e-06, 4.659501e-06, 4.842178e-06, 4.310014e-06, 4.45715e-06, 
    3.831832e-06, 4.243514e-06, 3.213126e-06, 3.926901e-06, 3.863819e-06, 
    4.25771e-06, 7.351496e-06, 6.660738e-06, 7.394141e-06, 7.291801e-06, 
    7.337596e-06, 7.912437e-06, 8.215352e-06, 8.879791e-06, 8.756128e-06, 
    8.269632e-06, 7.246154e-06, 7.581592e-06, 6.759235e-06, 6.776979e-06, 
    5.945905e-06, 6.309711e-06, 5.04005e-06, 5.3773e-06, 4.450925e-06, 
    4.670223e-06, 4.461019e-06, 4.523607e-06, 4.460209e-06, 4.785479e-06, 
    4.643748e-06, 4.938754e-06, 6.240221e-06, 5.831505e-06, 7.119197e-06, 
    7.997381e-06, 8.627014e-06, 9.097049e-06, 9.0294e-06, 8.901522e-06, 
    8.266848e-06, 7.703443e-06, 7.294973e-06, 7.031548e-06, 6.779533e-06, 
    6.060662e-06, 5.706211e-06, 4.974015e-06, 5.100096e-06, 4.888078e-06, 
    4.692531e-06, 4.378991e-06, 4.429349e-06, 4.295654e-06, 4.893609e-06, 
    4.488889e-06, 5.173084e-06, 4.977815e-06, 6.712064e-06, 7.489911e-06, 
    7.841411e-06, 8.159952e-06, 8.977651e-06, 8.40637e-06, 8.628029e-06, 
    8.108174e-06, 7.790954e-06, 7.946598e-06, 7.024454e-06, 7.372175e-06, 
    5.685748e-06, 6.368845e-06, 4.714995e-06, 5.074007e-06, 4.632193e-06, 
    4.853437e-06, 4.479582e-06, 4.814906e-06, 4.246794e-06, 4.130937e-06, 
    4.20981e-06, 3.913774e-06, 4.834092e-06, 4.461004e-06, 7.950983e-06, 
    7.925418e-06, 7.807207e-06, 8.337487e-06, 8.370846e-06, 8.883188e-06, 
    8.426156e-06, 8.237256e-06, 7.772894e-06, 7.50815e-06, 7.263228e-06, 
    6.74723e-06, 6.206309e-06, 5.509675e-06, 5.050061e-06, 4.760197e-06, 
    4.936248e-06, 4.780542e-06, 4.954873e-06, 5.038401e-06, 4.174016e-06, 
    4.642433e-06, 3.955216e-06, 3.990827e-06, 4.29251e-06, 3.9868e-06, 
    7.90751e-06, 8.05525e-06, 8.585198e-06, 8.168196e-06, 8.940447e-06, 
    8.50135e-06, 8.256691e-06, 7.364716e-06, 7.179528e-06, 7.011091e-06, 
    6.687816e-06, 6.29066e-06, 5.640367e-06, 5.120509e-06, 4.681367e-06, 
    4.712436e-06, 4.701477e-06, 4.607467e-06, 4.843258e-06, 4.569697e-06, 
    4.525071e-06, 4.642512e-06, 3.995616e-06, 4.172044e-06, 3.991587e-06, 
    4.10562e-06, 8.006994e-06, 7.760842e-06, 7.893089e-06, 7.645858e-06, 
    7.81936e-06, 7.071224e-06, 6.85848e-06, 5.930627e-06, 6.298277e-06, 
    5.721596e-06, 6.237638e-06, 6.143522e-06, 5.703454e-06, 6.20883e-06, 
    5.148062e-06, 5.849233e-06, 4.603845e-06, 5.242538e-06, 4.566097e-06, 
    4.683196e-06, 4.490684e-06, 4.323978e-06, 4.121797e-06, 3.769973e-06, 
    3.849046e-06, 3.570166e-06, 7.40514e-06, 7.106343e-06, 7.1323e-06, 
    6.829193e-06, 6.611763e-06, 6.159743e-06, 5.487529e-06, 5.732879e-06, 
    5.289196e-06, 5.203627e-06, 5.880455e-06, 5.456801e-06, 6.91187e-06, 
    6.657523e-06, 6.808065e-06, 7.381183e-06, 5.675504e-06, 6.505524e-06, 
    5.042734e-06, 5.440537e-06, 4.347417e-06, 4.865375e-06, 3.89318e-06, 
    3.207772e-06, 2.969701e-06, 2.707985e-06, 6.947448e-06, 7.145772e-06, 
    6.793861e-06, 6.33008e-06, 5.923182e-06, 5.415545e-06, 5.365713e-06, 
    5.275405e-06, 5.047372e-06, 4.862036e-06, 5.24708e-06, 4.816483e-06, 
    6.599543e-06, 5.60777e-06, 7.221883e-06, 6.700659e-06, 6.356705e-06, 
    6.505826e-06, 5.761495e-06, 5.596608e-06, 4.966071e-06, 5.284245e-06, 
    3.617978e-06, 4.289405e-06, 2.520336e-06, 2.831425e-06, 7.216115e-06, 
    6.948145e-06, 6.077315e-06, 6.4799e-06, 5.382995e-06, 5.137859e-06, 
    4.945513e-06, 4.70838e-06, 4.683384e-06, 4.548061e-06, 4.77157e-06, 
    4.556732e-06, 5.414504e-06, 5.015905e-06, 6.172168e-06, 5.872381e-06, 
    6.008796e-06, 6.161361e-06, 5.700415e-06, 5.240818e-06, 5.231402e-06, 
    5.090896e-06, 4.711689e-06, 5.378884e-06, 3.212792e-06, 4.59701e-06, 
    6.665121e-06, 6.187903e-06, 6.122145e-06, 6.302022e-06, 5.162008e-06, 
    5.553617e-06, 4.551327e-06, 4.805968e-06, 4.394792e-06, 4.59523e-06, 
    4.625359e-06, 4.895542e-06, 5.07032e-06, 5.535128e-06, 5.938751e-06, 
    6.275679e-06, 6.195985e-06, 5.830543e-06, 5.213744e-06, 4.681102e-06, 
    4.793693e-06, 4.42496e-06, 5.457015e-06, 5.00215e-06, 5.174052e-06, 
    4.735839e-06, 5.739506e-06, 4.874671e-06, 5.979718e-06, 5.875279e-06, 
    5.561632e-06, 4.972439e-06, 4.849448e-06, 4.720853e-06, 4.799872e-06, 
    5.198829e-06, 5.266774e-06, 5.569103e-06, 5.655019e-06, 5.897894e-06, 
    6.105337e-06, 5.915558e-06, 5.721463e-06, 5.198679e-06, 4.762094e-06, 
    4.321636e-06, 4.219298e-06, 3.758678e-06, 4.130076e-06, 3.208846e-06, 
    4.035324e-06, 2.956366e-06, 4.828163e-06, 4.051083e-06, 5.547714e-06, 
    5.367098e-06, 5.05271e-06, 4.389457e-06, 4.737825e-06, 4.332642e-06, 
    5.269455e-06, 5.818225e-06, 5.967675e-06, 6.254749e-06, 5.96124e-06, 
    5.984687e-06, 5.713582e-06, 5.799586e-06, 5.182025e-06, 5.506623e-06, 
    4.626104e-06, 4.335735e-06, 3.598523e-06, 2.957484e-06, 2.672946e-06, 
    2.553879e-06, 2.51842e-06, 2.503702e-06,
  8.089843e-09, 6.90219e-09, 7.123345e-09, 6.235644e-09, 6.718444e-09, 
    6.151081e-09, 7.838929e-09, 6.857555e-09, 7.473987e-09, 7.977826e-09, 
    4.727548e-09, 6.197863e-09, 3.464641e-09, 4.209748e-09, 2.510203e-09, 
    3.574375e-09, 2.324393e-09, 2.537612e-09, 1.931808e-09, 2.094521e-09, 
    1.431628e-09, 1.859556e-09, 1.147179e-09, 1.527334e-09, 1.46361e-09, 
    1.874911e-09, 5.880837e-09, 4.896473e-09, 5.942901e-09, 5.794202e-09, 
    5.86064e-09, 6.70819e-09, 7.164355e-09, 8.185915e-09, 7.993712e-09, 
    7.246752e-09, 5.728148e-09, 6.217371e-09, 5.034315e-09, 5.05924e-09, 
    3.92414e-09, 4.412615e-09, 2.774273e-09, 3.190306e-09, 2.08756e-09, 
    2.336762e-09, 2.098852e-09, 2.169258e-09, 2.097944e-09, 2.470876e-09, 
    2.306254e-09, 2.6524e-09, 4.318253e-09, 3.773469e-09, 5.545317e-09, 
    6.83547e-09, 7.794022e-09, 8.525775e-09, 8.419656e-09, 8.219785e-09, 
    7.242523e-09, 6.397211e-09, 5.7988e-09, 5.41987e-09, 5.06283e-09, 
    4.076721e-09, 3.610147e-09, 2.694655e-09, 2.847209e-09, 2.591994e-09, 
    2.362556e-09, 2.007607e-09, 2.063483e-09, 1.916136e-09, 2.598569e-09, 
    2.13012e-09, 2.936543e-09, 2.699221e-09, 4.968191e-09, 6.082792e-09, 
    6.602153e-09, 7.08046e-09, 8.33866e-09, 7.455179e-09, 7.795589e-09, 
    7.002237e-09, 6.527043e-09, 6.759317e-09, 5.409745e-09, 5.910914e-09, 
    3.583645e-09, 4.493294e-09, 2.38861e-09, 2.815457e-09, 2.292974e-09, 
    2.550921e-09, 2.119663e-09, 2.505451e-09, 1.8631e-09, 1.739147e-09, 
    1.823252e-09, 1.514003e-09, 2.528063e-09, 2.098835e-09, 6.765885e-09, 
    6.727608e-09, 6.551217e-09, 7.350029e-09, 7.400912e-09, 8.191207e-09, 
    7.485436e-09, 7.197583e-09, 6.500203e-09, 6.109515e-09, 5.752836e-09, 
    5.017468e-09, 4.272381e-09, 3.35768e-09, 2.786398e-09, 2.441279e-09, 
    2.649405e-09, 2.465088e-09, 2.671694e-09, 2.772277e-09, 1.784935e-09, 
    2.304742e-09, 1.556215e-09, 1.592776e-09, 1.912711e-09, 1.58863e-09, 
    6.700823e-09, 6.92247e-09, 7.729571e-09, 7.092932e-09, 8.280523e-09, 
    7.600662e-09, 7.22709e-09, 5.900061e-09, 5.632035e-09, 5.390683e-09, 
    4.934281e-09, 4.386697e-09, 3.525049e-09, 2.872119e-09, 2.349638e-09, 
    2.385638e-09, 2.372922e-09, 2.264631e-09, 2.538887e-09, 2.221531e-09, 
    2.170913e-09, 2.304832e-09, 1.597714e-09, 1.782831e-09, 1.59356e-09, 
    1.712407e-09, 6.849908e-09, 6.482305e-09, 6.679269e-09, 6.312084e-09, 
    6.569306e-09, 5.476577e-09, 5.174083e-09, 3.903934e-09, 4.397055e-09, 
    3.630104e-09, 4.314757e-09, 4.187763e-09, 3.606573e-09, 4.275788e-09, 
    2.905835e-09, 3.796722e-09, 2.260488e-09, 3.022226e-09, 2.217434e-09, 
    2.351753e-09, 2.132138e-09, 1.947083e-09, 1.729478e-09, 1.370425e-09, 
    1.448811e-09, 1.17881e-09, 5.958931e-09, 5.52688e-09, 5.564126e-09, 
    5.132748e-09, 4.828267e-09, 4.209586e-09, 3.329526e-09, 3.644758e-09, 
    3.08015e-09, 2.974143e-09, 3.83776e-09, 3.290562e-09, 5.24963e-09, 
    4.89199e-09, 5.102974e-09, 5.924027e-09, 3.570398e-09, 4.681076e-09, 
    2.777523e-09, 3.269987e-09, 1.972803e-09, 2.565055e-09, 1.493163e-09, 
    1.140588e-09, 8.646351e-10, 6.018308e-10, 5.300111e-09, 5.583478e-09, 
    5.08298e-09, 4.440366e-09, 3.894097e-09, 3.238435e-09, 3.175762e-09, 
    3.063e-09, 2.78314e-09, 2.561101e-09, 3.027853e-09, 2.507307e-09, 
    4.811282e-09, 3.483111e-09, 5.693093e-09, 4.952236e-09, 4.476703e-09, 
    4.681492e-09, 3.681988e-09, 3.46878e-09, 2.68512e-09, 3.07399e-09, 
    1.223791e-09, 1.909328e-09, 4.413376e-10, 7.202954e-10, 5.68477e-09, 
    5.301101e-09, 4.09898e-09, 4.645734e-09, 3.197461e-09, 2.893338e-09, 
    2.660486e-09, 2.38093e-09, 2.35197e-09, 2.196948e-09, 2.45458e-09, 
    2.20679e-09, 3.237123e-09, 2.745089e-09, 4.226319e-09, 3.827138e-09, 
    4.007584e-09, 4.211764e-09, 3.602636e-09, 3.020097e-09, 3.008444e-09, 
    2.836002e-09, 2.384771e-09, 3.192297e-09, 1.146766e-09, 2.252675e-09, 
    4.902589e-09, 4.247533e-09, 4.159046e-09, 4.402151e-09, 2.922939e-09, 
    3.413722e-09, 2.200654e-09, 2.494935e-09, 2.025091e-09, 2.250641e-09, 
    2.28513e-09, 2.600868e-09, 2.810978e-09, 3.390113e-09, 3.914675e-09, 
    4.366342e-09, 4.258441e-09, 3.772208e-09, 2.986626e-09, 2.349331e-09, 
    2.480513e-09, 2.058595e-09, 3.290833e-09, 2.728501e-09, 2.937733e-09, 
    2.412857e-09, 3.653371e-09, 2.576076e-09, 3.96895e-09, 3.830949e-09, 
    3.42397e-09, 2.692763e-09, 2.546204e-09, 2.395417e-09, 2.48777e-09, 
    2.968228e-09, 3.052279e-09, 3.433529e-09, 3.543942e-09, 3.86073e-09, 
    4.136501e-09, 3.88403e-09, 3.629931e-09, 2.968043e-09, 2.443496e-09, 
    1.944519e-09, 1.83345e-09, 1.359344e-09, 1.738235e-09, 1.141908e-09, 
    1.638831e-09, 8.50192e-10, 2.521069e-09, 1.655238e-09, 3.40618e-09, 
    3.177499e-09, 2.789608e-09, 2.019183e-09, 2.415171e-09, 1.956579e-09, 
    3.055608e-09, 3.756072e-09, 3.952976e-09, 4.337941e-09, 3.944447e-09, 
    3.975545e-09, 3.619705e-09, 3.731691e-09, 2.947536e-09, 3.353796e-09, 
    2.285985e-09, 1.959972e-09, 1.20542e-09, 8.513987e-10, 5.700416e-10, 
    4.682471e-10, 4.398246e-10, 4.28286e-10,
  4.32761e-13, 4.280987e-13, 4.289675e-13, 4.254785e-13, 4.273767e-13, 
    4.251458e-13, 4.317767e-13, 4.279234e-13, 4.303444e-13, 4.323216e-13, 
    4.195388e-13, 4.253299e-13, 4.14551e-13, 4.174954e-13, 4.107719e-13, 
    4.149849e-13, 4.100349e-13, 4.108805e-13, 4.084764e-13, 4.091226e-13, 
    4.064874e-13, 4.081893e-13, 4.053598e-13, 4.068683e-13, 4.066147e-13, 
    4.082503e-13, 4.240825e-13, 4.20205e-13, 4.243268e-13, 4.237415e-13, 
    4.24003e-13, 4.273364e-13, 4.291286e-13, 4.331378e-13, 4.323839e-13, 
    4.294522e-13, 4.234815e-13, 4.254066e-13, 4.207484e-13, 4.208466e-13, 
    4.163674e-13, 4.182963e-13, 4.118184e-13, 4.134656e-13, 4.09095e-13, 
    4.10084e-13, 4.091398e-13, 4.094193e-13, 4.091362e-13, 4.106159e-13, 
    4.099629e-13, 4.113355e-13, 4.179238e-13, 4.15772e-13, 4.227616e-13, 
    4.278366e-13, 4.316004e-13, 4.344703e-13, 4.340543e-13, 4.332706e-13, 
    4.294356e-13, 4.261139e-13, 4.237596e-13, 4.222676e-13, 4.208608e-13, 
    4.169701e-13, 4.151264e-13, 4.11503e-13, 4.121074e-13, 4.110961e-13, 
    4.101863e-13, 4.087775e-13, 4.089994e-13, 4.084141e-13, 4.111222e-13, 
    4.092639e-13, 4.124612e-13, 4.115211e-13, 4.204877e-13, 4.248772e-13, 
    4.269196e-13, 4.287991e-13, 4.337367e-13, 4.302706e-13, 4.316066e-13, 
    4.284918e-13, 4.266243e-13, 4.275373e-13, 4.222277e-13, 4.242009e-13, 
    4.150216e-13, 4.186147e-13, 4.102897e-13, 4.119816e-13, 4.099103e-13, 
    4.109333e-13, 4.092224e-13, 4.10753e-13, 4.082034e-13, 4.077107e-13, 
    4.08045e-13, 4.068152e-13, 4.108427e-13, 4.091397e-13, 4.275631e-13, 
    4.274127e-13, 4.267194e-13, 4.298577e-13, 4.300575e-13, 4.331585e-13, 
    4.303893e-13, 4.292591e-13, 4.265188e-13, 4.249823e-13, 4.235787e-13, 
    4.20682e-13, 4.177427e-13, 4.141279e-13, 4.118665e-13, 4.104985e-13, 
    4.113236e-13, 4.10593e-13, 4.11412e-13, 4.118105e-13, 4.078927e-13, 
    4.09957e-13, 4.069832e-13, 4.071286e-13, 4.084005e-13, 4.071121e-13, 
    4.273074e-13, 4.281784e-13, 4.313476e-13, 4.288481e-13, 4.335088e-13, 
    4.308416e-13, 4.29375e-13, 4.241582e-13, 4.231031e-13, 4.221526e-13, 
    4.20354e-13, 4.18194e-13, 4.147899e-13, 4.12206e-13, 4.101351e-13, 
    4.102779e-13, 4.102274e-13, 4.097978e-13, 4.108856e-13, 4.096268e-13, 
    4.094259e-13, 4.099573e-13, 4.071483e-13, 4.078844e-13, 4.071318e-13, 
    4.076044e-13, 4.278933e-13, 4.264485e-13, 4.272227e-13, 4.257791e-13, 
    4.267905e-13, 4.224909e-13, 4.212992e-13, 4.162876e-13, 4.182349e-13, 
    4.152053e-13, 4.1791e-13, 4.174086e-13, 4.151123e-13, 4.177562e-13, 
    4.123395e-13, 4.158639e-13, 4.097814e-13, 4.128004e-13, 4.096105e-13, 
    4.101435e-13, 4.09272e-13, 4.085371e-13, 4.076723e-13, 4.062438e-13, 
    4.065558e-13, 4.054805e-13, 4.243898e-13, 4.22689e-13, 4.228357e-13, 
    4.211363e-13, 4.19936e-13, 4.174948e-13, 4.140165e-13, 4.152632e-13, 
    4.130297e-13, 4.1261e-13, 4.160261e-13, 4.138623e-13, 4.215969e-13, 
    4.201873e-13, 4.21019e-13, 4.242525e-13, 4.149692e-13, 4.193555e-13, 
    4.118313e-13, 4.137809e-13, 4.086392e-13, 4.109893e-13, 4.067323e-13, 
    4.053335e-13, 4.042316e-13, 4.031807e-13, 4.217958e-13, 4.229119e-13, 
    4.209402e-13, 4.184058e-13, 4.162487e-13, 4.136561e-13, 4.134081e-13, 
    4.129618e-13, 4.118536e-13, 4.109736e-13, 4.128227e-13, 4.107604e-13, 
    4.19869e-13, 4.14624e-13, 4.233435e-13, 4.204248e-13, 4.185492e-13, 
    4.193571e-13, 4.154104e-13, 4.145674e-13, 4.114652e-13, 4.130053e-13, 
    4.056597e-13, 4.083871e-13, 4.025382e-13, 4.036546e-13, 4.233107e-13, 
    4.217997e-13, 4.17058e-13, 4.192161e-13, 4.13494e-13, 4.1229e-13, 
    4.113676e-13, 4.102592e-13, 4.101443e-13, 4.095292e-13, 4.105513e-13, 
    4.095683e-13, 4.136509e-13, 4.117028e-13, 4.175609e-13, 4.159841e-13, 
    4.166971e-13, 4.175034e-13, 4.150967e-13, 4.12792e-13, 4.127458e-13, 
    4.12063e-13, 4.102744e-13, 4.134735e-13, 4.053582e-13, 4.097504e-13, 
    4.202291e-13, 4.176446e-13, 4.172952e-13, 4.18255e-13, 4.124073e-13, 
    4.143496e-13, 4.095439e-13, 4.107113e-13, 4.088469e-13, 4.097423e-13, 
    4.098791e-13, 4.111313e-13, 4.119638e-13, 4.142562e-13, 4.1633e-13, 
    4.181137e-13, 4.176877e-13, 4.15767e-13, 4.126595e-13, 4.101338e-13, 
    4.106541e-13, 4.0898e-13, 4.138634e-13, 4.116371e-13, 4.124659e-13, 
    4.103858e-13, 4.152973e-13, 4.11033e-13, 4.165444e-13, 4.159992e-13, 
    4.143901e-13, 4.114955e-13, 4.109146e-13, 4.103167e-13, 4.106829e-13, 
    4.125866e-13, 4.129194e-13, 4.144279e-13, 4.148646e-13, 4.161168e-13, 
    4.172062e-13, 4.162089e-13, 4.152046e-13, 4.125859e-13, 4.105073e-13, 
    4.085269e-13, 4.080856e-13, 4.061996e-13, 4.077071e-13, 4.053388e-13, 
    4.073118e-13, 4.041739e-13, 4.108149e-13, 4.073771e-13, 4.143197e-13, 
    4.13415e-13, 4.118792e-13, 4.088234e-13, 4.10395e-13, 4.085748e-13, 
    4.129325e-13, 4.157033e-13, 4.164813e-13, 4.180015e-13, 4.164476e-13, 
    4.165705e-13, 4.151642e-13, 4.156069e-13, 4.125047e-13, 4.141125e-13, 
    4.098825e-13, 4.085883e-13, 4.055865e-13, 4.041787e-13, 4.030535e-13, 
    4.02646e-13, 4.025321e-13, 4.024859e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.94965e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949653e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.94965e-07, 8.949651e-07, 8.949648e-07, 8.949649e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.94965e-07, 8.949651e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.01737e-16, 6.033623e-16, 6.030466e-16, 6.043563e-16, 6.036301e-16, 
    6.044873e-16, 6.020669e-16, 6.034266e-16, 6.025589e-16, 6.018837e-16, 
    6.068941e-16, 6.044148e-16, 6.094675e-16, 6.07889e-16, 6.118515e-16, 
    6.092216e-16, 6.123814e-16, 6.117762e-16, 6.135982e-16, 6.130765e-16, 
    6.154034e-16, 6.13839e-16, 6.166091e-16, 6.150302e-16, 6.152771e-16, 
    6.137872e-16, 6.049145e-16, 6.065855e-16, 6.048154e-16, 6.050538e-16, 
    6.049469e-16, 6.036449e-16, 6.029881e-16, 6.016131e-16, 6.018629e-16, 
    6.028729e-16, 6.05161e-16, 6.04385e-16, 6.06341e-16, 6.062969e-16, 
    6.084711e-16, 6.074912e-16, 6.111412e-16, 6.10105e-16, 6.130983e-16, 
    6.123459e-16, 6.130629e-16, 6.128456e-16, 6.130657e-16, 6.119621e-16, 
    6.12435e-16, 6.114637e-16, 6.076746e-16, 6.087892e-16, 6.054625e-16, 
    6.03458e-16, 6.021265e-16, 6.011806e-16, 6.013143e-16, 6.015692e-16, 
    6.028788e-16, 6.041097e-16, 6.050469e-16, 6.056733e-16, 6.062905e-16, 
    6.081556e-16, 6.09143e-16, 6.113504e-16, 6.109526e-16, 6.116267e-16, 
    6.122711e-16, 6.133516e-16, 6.131739e-16, 6.136496e-16, 6.116093e-16, 
    6.129655e-16, 6.107263e-16, 6.113387e-16, 6.064564e-16, 6.045945e-16, 
    6.038009e-16, 6.031073e-16, 6.014171e-16, 6.025844e-16, 6.021243e-16, 
    6.03219e-16, 6.03914e-16, 6.035704e-16, 6.056905e-16, 6.048665e-16, 
    6.092015e-16, 6.073358e-16, 6.121959e-16, 6.110343e-16, 6.124743e-16, 
    6.117398e-16, 6.12998e-16, 6.118656e-16, 6.138268e-16, 6.142533e-16, 
    6.139619e-16, 6.150819e-16, 6.118028e-16, 6.130627e-16, 6.035607e-16, 
    6.036167e-16, 6.03878e-16, 6.027293e-16, 6.026591e-16, 6.016062e-16, 
    6.025432e-16, 6.029419e-16, 6.039544e-16, 6.045526e-16, 6.051212e-16, 
    6.063707e-16, 6.077645e-16, 6.097121e-16, 6.111097e-16, 6.120459e-16, 
    6.11472e-16, 6.119787e-16, 6.114122e-16, 6.111467e-16, 6.140934e-16, 
    6.124393e-16, 6.149208e-16, 6.147837e-16, 6.136609e-16, 6.147991e-16, 
    6.036561e-16, 6.033335e-16, 6.022126e-16, 6.030899e-16, 6.014915e-16, 
    6.023862e-16, 6.029003e-16, 6.048833e-16, 6.053191e-16, 6.057226e-16, 
    6.065195e-16, 6.075413e-16, 6.093322e-16, 6.108886e-16, 6.123086e-16, 
    6.122047e-16, 6.122412e-16, 6.125581e-16, 6.117728e-16, 6.12687e-16, 
    6.128402e-16, 6.124393e-16, 6.147653e-16, 6.141012e-16, 6.147807e-16, 
    6.143484e-16, 6.034384e-16, 6.039811e-16, 6.036879e-16, 6.042392e-16, 
    6.038507e-16, 6.055771e-16, 6.060943e-16, 6.085128e-16, 6.075211e-16, 
    6.090995e-16, 6.076817e-16, 6.079329e-16, 6.091501e-16, 6.077584e-16, 
    6.108024e-16, 6.087388e-16, 6.125704e-16, 6.105113e-16, 6.126994e-16, 
    6.123025e-16, 6.129597e-16, 6.135478e-16, 6.142878e-16, 6.156517e-16, 
    6.15336e-16, 6.164761e-16, 6.0479e-16, 6.054931e-16, 6.054316e-16, 
    6.061674e-16, 6.067112e-16, 6.078896e-16, 6.097774e-16, 6.090679e-16, 
    6.103706e-16, 6.106319e-16, 6.086529e-16, 6.09868e-16, 6.059638e-16, 
    6.065949e-16, 6.062194e-16, 6.048453e-16, 6.09231e-16, 6.069816e-16, 
    6.111327e-16, 6.099164e-16, 6.13464e-16, 6.117002e-16, 6.151621e-16, 
    6.166387e-16, 6.180287e-16, 6.196494e-16, 6.058772e-16, 6.053995e-16, 
    6.062549e-16, 6.07437e-16, 6.08534e-16, 6.099906e-16, 6.101397e-16, 
    6.104123e-16, 6.111183e-16, 6.117117e-16, 6.104982e-16, 6.118605e-16, 
    6.067406e-16, 6.094262e-16, 6.052185e-16, 6.064863e-16, 6.073675e-16, 
    6.069814e-16, 6.089869e-16, 6.094591e-16, 6.113759e-16, 6.103857e-16, 
    6.162741e-16, 6.136716e-16, 6.208835e-16, 6.188714e-16, 6.052325e-16, 
    6.058756e-16, 6.081114e-16, 6.070481e-16, 6.10088e-16, 6.108348e-16, 
    6.114423e-16, 6.122178e-16, 6.123018e-16, 6.127611e-16, 6.120083e-16, 
    6.127315e-16, 6.099937e-16, 6.112177e-16, 6.078565e-16, 6.086751e-16, 
    6.082987e-16, 6.078854e-16, 6.091605e-16, 6.105172e-16, 6.105467e-16, 
    6.109811e-16, 6.122043e-16, 6.101003e-16, 6.166086e-16, 6.125914e-16, 
    6.065767e-16, 6.078134e-16, 6.079906e-16, 6.075116e-16, 6.107603e-16, 
    6.095838e-16, 6.1275e-16, 6.11895e-16, 6.132958e-16, 6.125999e-16, 
    6.124974e-16, 6.116031e-16, 6.110459e-16, 6.096377e-16, 6.084909e-16, 
    6.075811e-16, 6.077927e-16, 6.087919e-16, 6.106003e-16, 6.123092e-16, 
    6.119348e-16, 6.131894e-16, 6.098677e-16, 6.11261e-16, 6.107227e-16, 
    6.121266e-16, 6.090489e-16, 6.116684e-16, 6.083784e-16, 6.086673e-16, 
    6.095605e-16, 6.113551e-16, 6.117527e-16, 6.121762e-16, 6.11915e-16, 
    6.106463e-16, 6.104385e-16, 6.095389e-16, 6.092902e-16, 6.086044e-16, 
    6.080362e-16, 6.085553e-16, 6.091e-16, 6.106471e-16, 6.120392e-16, 
    6.135562e-16, 6.139274e-16, 6.15696e-16, 6.142556e-16, 6.166309e-16, 
    6.146105e-16, 6.181067e-16, 6.118208e-16, 6.145522e-16, 6.096013e-16, 
    6.101356e-16, 6.111007e-16, 6.133137e-16, 6.1212e-16, 6.135162e-16, 
    6.104304e-16, 6.088261e-16, 6.084114e-16, 6.076363e-16, 6.084292e-16, 
    6.083647e-16, 6.09123e-16, 6.088794e-16, 6.106984e-16, 6.097216e-16, 
    6.124947e-16, 6.135053e-16, 6.163565e-16, 6.181012e-16, 6.19876e-16, 
    6.206586e-16, 6.208967e-16, 6.209962e-16 ;

 CWDC_TO_LITR2C =
  4.573201e-16, 4.585554e-16, 4.583154e-16, 4.593108e-16, 4.587589e-16, 
    4.594104e-16, 4.575709e-16, 4.586042e-16, 4.579448e-16, 4.574316e-16, 
    4.612395e-16, 4.593552e-16, 4.631953e-16, 4.619956e-16, 4.650072e-16, 
    4.630084e-16, 4.654099e-16, 4.649499e-16, 4.663347e-16, 4.659382e-16, 
    4.677066e-16, 4.665176e-16, 4.686229e-16, 4.67423e-16, 4.676106e-16, 
    4.664783e-16, 4.59735e-16, 4.61005e-16, 4.596597e-16, 4.598409e-16, 
    4.597597e-16, 4.587701e-16, 4.582709e-16, 4.572259e-16, 4.574158e-16, 
    4.581834e-16, 4.599224e-16, 4.593326e-16, 4.608192e-16, 4.607856e-16, 
    4.624381e-16, 4.616933e-16, 4.644673e-16, 4.636798e-16, 4.659547e-16, 
    4.653829e-16, 4.659278e-16, 4.657627e-16, 4.6593e-16, 4.650912e-16, 
    4.654506e-16, 4.647125e-16, 4.618328e-16, 4.626797e-16, 4.601515e-16, 
    4.586281e-16, 4.576161e-16, 4.568972e-16, 4.569989e-16, 4.571925e-16, 
    4.581879e-16, 4.591234e-16, 4.598356e-16, 4.603117e-16, 4.607808e-16, 
    4.621982e-16, 4.629487e-16, 4.646263e-16, 4.64324e-16, 4.648363e-16, 
    4.65326e-16, 4.661472e-16, 4.660122e-16, 4.663737e-16, 4.64823e-16, 
    4.658538e-16, 4.64152e-16, 4.646174e-16, 4.609069e-16, 4.594918e-16, 
    4.588887e-16, 4.583615e-16, 4.57077e-16, 4.579641e-16, 4.576145e-16, 
    4.584465e-16, 4.589746e-16, 4.587135e-16, 4.603248e-16, 4.596985e-16, 
    4.629931e-16, 4.615752e-16, 4.652689e-16, 4.643861e-16, 4.654804e-16, 
    4.649222e-16, 4.658784e-16, 4.650179e-16, 4.665084e-16, 4.668325e-16, 
    4.66611e-16, 4.674622e-16, 4.649701e-16, 4.659277e-16, 4.587061e-16, 
    4.587487e-16, 4.589472e-16, 4.580743e-16, 4.580209e-16, 4.572207e-16, 
    4.579329e-16, 4.582359e-16, 4.590054e-16, 4.5946e-16, 4.598921e-16, 
    4.608417e-16, 4.61901e-16, 4.633812e-16, 4.644433e-16, 4.651549e-16, 
    4.647187e-16, 4.651038e-16, 4.646732e-16, 4.644715e-16, 4.66711e-16, 
    4.654539e-16, 4.673398e-16, 4.672356e-16, 4.663823e-16, 4.672474e-16, 
    4.587786e-16, 4.585335e-16, 4.576816e-16, 4.583483e-16, 4.571335e-16, 
    4.578135e-16, 4.582042e-16, 4.597114e-16, 4.600425e-16, 4.603492e-16, 
    4.609548e-16, 4.617314e-16, 4.630924e-16, 4.642753e-16, 4.653546e-16, 
    4.652756e-16, 4.653034e-16, 4.655442e-16, 4.649473e-16, 4.656421e-16, 
    4.657585e-16, 4.654539e-16, 4.672216e-16, 4.667169e-16, 4.672334e-16, 
    4.669048e-16, 4.586132e-16, 4.590257e-16, 4.588028e-16, 4.592218e-16, 
    4.589265e-16, 4.602386e-16, 4.606317e-16, 4.624697e-16, 4.61716e-16, 
    4.629156e-16, 4.61838e-16, 4.62029e-16, 4.629541e-16, 4.618964e-16, 
    4.642099e-16, 4.626415e-16, 4.655536e-16, 4.639886e-16, 4.656515e-16, 
    4.653499e-16, 4.658494e-16, 4.662963e-16, 4.668587e-16, 4.678952e-16, 
    4.676554e-16, 4.685219e-16, 4.596404e-16, 4.601748e-16, 4.60128e-16, 
    4.606872e-16, 4.611005e-16, 4.619961e-16, 4.634308e-16, 4.628916e-16, 
    4.638817e-16, 4.640802e-16, 4.625762e-16, 4.634996e-16, 4.605325e-16, 
    4.610121e-16, 4.607268e-16, 4.596825e-16, 4.630155e-16, 4.61306e-16, 
    4.644608e-16, 4.635365e-16, 4.662326e-16, 4.648922e-16, 4.675232e-16, 
    4.686454e-16, 4.697018e-16, 4.709336e-16, 4.604666e-16, 4.601036e-16, 
    4.607537e-16, 4.616521e-16, 4.624858e-16, 4.635929e-16, 4.637062e-16, 
    4.639134e-16, 4.644499e-16, 4.649009e-16, 4.639786e-16, 4.65014e-16, 
    4.611228e-16, 4.63164e-16, 4.599661e-16, 4.609297e-16, 4.615993e-16, 
    4.613058e-16, 4.6283e-16, 4.631889e-16, 4.646456e-16, 4.638931e-16, 
    4.683684e-16, 4.663904e-16, 4.718714e-16, 4.703423e-16, 4.599767e-16, 
    4.604655e-16, 4.621647e-16, 4.613566e-16, 4.636668e-16, 4.642345e-16, 
    4.646961e-16, 4.652855e-16, 4.653494e-16, 4.656984e-16, 4.651263e-16, 
    4.65676e-16, 4.635952e-16, 4.645254e-16, 4.619709e-16, 4.625931e-16, 
    4.62307e-16, 4.619929e-16, 4.62962e-16, 4.639931e-16, 4.640156e-16, 
    4.643456e-16, 4.652753e-16, 4.636762e-16, 4.686226e-16, 4.655694e-16, 
    4.609983e-16, 4.619382e-16, 4.620728e-16, 4.617088e-16, 4.641778e-16, 
    4.632837e-16, 4.6569e-16, 4.650402e-16, 4.661048e-16, 4.655759e-16, 
    4.65498e-16, 4.648183e-16, 4.643949e-16, 4.633246e-16, 4.62453e-16, 
    4.617617e-16, 4.619225e-16, 4.626818e-16, 4.640562e-16, 4.653549e-16, 
    4.650705e-16, 4.66024e-16, 4.634995e-16, 4.645583e-16, 4.641492e-16, 
    4.652162e-16, 4.628772e-16, 4.648679e-16, 4.623676e-16, 4.625871e-16, 
    4.63266e-16, 4.646299e-16, 4.649321e-16, 4.652539e-16, 4.650554e-16, 
    4.640912e-16, 4.639333e-16, 4.632496e-16, 4.630605e-16, 4.625394e-16, 
    4.621075e-16, 4.62502e-16, 4.62916e-16, 4.640918e-16, 4.651498e-16, 
    4.663026e-16, 4.665848e-16, 4.679289e-16, 4.668343e-16, 4.686395e-16, 
    4.67104e-16, 4.697611e-16, 4.649838e-16, 4.670597e-16, 4.63297e-16, 
    4.637031e-16, 4.644365e-16, 4.661184e-16, 4.652111e-16, 4.662723e-16, 
    4.639271e-16, 4.627078e-16, 4.623927e-16, 4.618036e-16, 4.624061e-16, 
    4.623572e-16, 4.629335e-16, 4.627483e-16, 4.641308e-16, 4.633884e-16, 
    4.65496e-16, 4.662641e-16, 4.684309e-16, 4.69757e-16, 4.711058e-16, 
    4.717005e-16, 4.718815e-16, 4.719571e-16 ;

 CWDC_TO_LITR3C =
  1.444169e-16, 1.44807e-16, 1.447312e-16, 1.450455e-16, 1.448712e-16, 
    1.45077e-16, 1.444961e-16, 1.448224e-16, 1.446141e-16, 1.444521e-16, 
    1.456546e-16, 1.450595e-16, 1.462722e-16, 1.458934e-16, 1.468444e-16, 
    1.462132e-16, 1.469715e-16, 1.468263e-16, 1.472636e-16, 1.471384e-16, 
    1.476968e-16, 1.473214e-16, 1.479862e-16, 1.476073e-16, 1.476665e-16, 
    1.473089e-16, 1.451795e-16, 1.455805e-16, 1.451557e-16, 1.452129e-16, 
    1.451873e-16, 1.448748e-16, 1.447171e-16, 1.443871e-16, 1.444471e-16, 
    1.446895e-16, 1.452386e-16, 1.450524e-16, 1.455218e-16, 1.455112e-16, 
    1.460331e-16, 1.457979e-16, 1.466739e-16, 1.464252e-16, 1.471436e-16, 
    1.46963e-16, 1.471351e-16, 1.470829e-16, 1.471358e-16, 1.468709e-16, 
    1.469844e-16, 1.467513e-16, 1.458419e-16, 1.461094e-16, 1.45311e-16, 
    1.448299e-16, 1.445104e-16, 1.442833e-16, 1.443154e-16, 1.443766e-16, 
    1.446909e-16, 1.449863e-16, 1.452112e-16, 1.453616e-16, 1.455097e-16, 
    1.459573e-16, 1.461943e-16, 1.467241e-16, 1.466286e-16, 1.467904e-16, 
    1.469451e-16, 1.472044e-16, 1.471617e-16, 1.472759e-16, 1.467862e-16, 
    1.471117e-16, 1.465743e-16, 1.467213e-16, 1.455495e-16, 1.451027e-16, 
    1.449122e-16, 1.447457e-16, 1.443401e-16, 1.446202e-16, 1.445098e-16, 
    1.447726e-16, 1.449394e-16, 1.448569e-16, 1.453657e-16, 1.45168e-16, 
    1.462084e-16, 1.457606e-16, 1.46927e-16, 1.466482e-16, 1.469938e-16, 
    1.468175e-16, 1.471195e-16, 1.468478e-16, 1.473184e-16, 1.474208e-16, 
    1.473508e-16, 1.476196e-16, 1.468327e-16, 1.47135e-16, 1.448546e-16, 
    1.44868e-16, 1.449307e-16, 1.44655e-16, 1.446382e-16, 1.443855e-16, 
    1.446104e-16, 1.447061e-16, 1.449491e-16, 1.450926e-16, 1.452291e-16, 
    1.45529e-16, 1.458635e-16, 1.463309e-16, 1.466663e-16, 1.46891e-16, 
    1.467533e-16, 1.468749e-16, 1.467389e-16, 1.466752e-16, 1.473824e-16, 
    1.469854e-16, 1.47581e-16, 1.475481e-16, 1.472786e-16, 1.475518e-16, 
    1.448775e-16, 1.448e-16, 1.44531e-16, 1.447416e-16, 1.44358e-16, 
    1.445727e-16, 1.446961e-16, 1.45172e-16, 1.452766e-16, 1.453734e-16, 
    1.455647e-16, 1.458099e-16, 1.462397e-16, 1.466133e-16, 1.469541e-16, 
    1.469291e-16, 1.469379e-16, 1.47014e-16, 1.468255e-16, 1.470449e-16, 
    1.470816e-16, 1.469854e-16, 1.475437e-16, 1.473843e-16, 1.475474e-16, 
    1.474436e-16, 1.448252e-16, 1.449555e-16, 1.448851e-16, 1.450174e-16, 
    1.449242e-16, 1.453385e-16, 1.454626e-16, 1.460431e-16, 1.458051e-16, 
    1.461839e-16, 1.458436e-16, 1.459039e-16, 1.46196e-16, 1.45862e-16, 
    1.465926e-16, 1.460973e-16, 1.470169e-16, 1.465227e-16, 1.470478e-16, 
    1.469526e-16, 1.471103e-16, 1.472515e-16, 1.474291e-16, 1.477564e-16, 
    1.476806e-16, 1.479543e-16, 1.451496e-16, 1.453184e-16, 1.453036e-16, 
    1.454802e-16, 1.456107e-16, 1.458935e-16, 1.463466e-16, 1.461763e-16, 
    1.464889e-16, 1.465517e-16, 1.460767e-16, 1.463683e-16, 1.454313e-16, 
    1.455828e-16, 1.454927e-16, 1.451629e-16, 1.462154e-16, 1.456756e-16, 
    1.466718e-16, 1.463799e-16, 1.472313e-16, 1.468081e-16, 1.476389e-16, 
    1.479933e-16, 1.483269e-16, 1.487159e-16, 1.454105e-16, 1.452959e-16, 
    1.455012e-16, 1.457849e-16, 1.460482e-16, 1.463977e-16, 1.464335e-16, 
    1.46499e-16, 1.466684e-16, 1.468108e-16, 1.465196e-16, 1.468465e-16, 
    1.456177e-16, 1.462623e-16, 1.452525e-16, 1.455567e-16, 1.457682e-16, 
    1.456755e-16, 1.461569e-16, 1.462702e-16, 1.467302e-16, 1.464926e-16, 
    1.479058e-16, 1.472812e-16, 1.49012e-16, 1.485291e-16, 1.452558e-16, 
    1.454102e-16, 1.459467e-16, 1.456915e-16, 1.464211e-16, 1.466004e-16, 
    1.467461e-16, 1.469323e-16, 1.469524e-16, 1.470627e-16, 1.46882e-16, 
    1.470556e-16, 1.463985e-16, 1.466922e-16, 1.458855e-16, 1.46082e-16, 
    1.459917e-16, 1.458925e-16, 1.461985e-16, 1.465241e-16, 1.465312e-16, 
    1.466355e-16, 1.46929e-16, 1.464241e-16, 1.479861e-16, 1.470219e-16, 
    1.455784e-16, 1.458752e-16, 1.459177e-16, 1.458028e-16, 1.465825e-16, 
    1.463001e-16, 1.4706e-16, 1.468548e-16, 1.47191e-16, 1.47024e-16, 
    1.469994e-16, 1.467847e-16, 1.46651e-16, 1.46313e-16, 1.460378e-16, 
    1.458195e-16, 1.458703e-16, 1.461101e-16, 1.465441e-16, 1.469542e-16, 
    1.468644e-16, 1.471655e-16, 1.463683e-16, 1.467026e-16, 1.465734e-16, 
    1.469104e-16, 1.461717e-16, 1.468004e-16, 1.460108e-16, 1.460801e-16, 
    1.462945e-16, 1.467252e-16, 1.468207e-16, 1.469223e-16, 1.468596e-16, 
    1.465551e-16, 1.465052e-16, 1.462893e-16, 1.462297e-16, 1.460651e-16, 
    1.459287e-16, 1.460533e-16, 1.46184e-16, 1.465553e-16, 1.468894e-16, 
    1.472535e-16, 1.473426e-16, 1.47767e-16, 1.474213e-16, 1.479914e-16, 
    1.475065e-16, 1.483456e-16, 1.46837e-16, 1.474925e-16, 1.463043e-16, 
    1.464326e-16, 1.466642e-16, 1.471953e-16, 1.469088e-16, 1.472439e-16, 
    1.465033e-16, 1.461183e-16, 1.460188e-16, 1.458327e-16, 1.46023e-16, 
    1.460075e-16, 1.461895e-16, 1.461311e-16, 1.465676e-16, 1.463332e-16, 
    1.469987e-16, 1.472413e-16, 1.479256e-16, 1.483443e-16, 1.487702e-16, 
    1.489581e-16, 1.490152e-16, 1.490391e-16 ;

 CWDC_vr =
  5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  9.146403e-19, 9.171108e-19, 9.166309e-19, 9.186216e-19, 9.175177e-19, 
    9.188207e-19, 9.151417e-19, 9.172085e-19, 9.158895e-19, 9.148633e-19, 
    9.224791e-19, 9.187104e-19, 9.263906e-19, 9.239912e-19, 9.300143e-19, 
    9.260169e-19, 9.308197e-19, 9.298999e-19, 9.326693e-19, 9.318763e-19, 
    9.354132e-19, 9.330352e-19, 9.372458e-19, 9.348459e-19, 9.352213e-19, 
    9.329566e-19, 9.194701e-19, 9.220099e-19, 9.193193e-19, 9.196817e-19, 
    9.195193e-19, 9.175403e-19, 9.165419e-19, 9.144519e-19, 9.148316e-19, 
    9.163669e-19, 9.198447e-19, 9.186652e-19, 9.216383e-19, 9.215712e-19, 
    9.248761e-19, 9.233866e-19, 9.289346e-19, 9.273596e-19, 9.319094e-19, 
    9.307658e-19, 9.318556e-19, 9.315253e-19, 9.318599e-19, 9.301824e-19, 
    9.309012e-19, 9.294249e-19, 9.236654e-19, 9.253595e-19, 9.203031e-19, 
    9.172561e-19, 9.152322e-19, 9.137945e-19, 9.139978e-19, 9.143851e-19, 
    9.163758e-19, 9.182467e-19, 9.196712e-19, 9.206235e-19, 9.215615e-19, 
    9.243965e-19, 9.258973e-19, 9.292526e-19, 9.286481e-19, 9.296726e-19, 
    9.30652e-19, 9.322945e-19, 9.320243e-19, 9.327475e-19, 9.296461e-19, 
    9.317075e-19, 9.28304e-19, 9.292348e-19, 9.218138e-19, 9.189836e-19, 
    9.177774e-19, 9.16723e-19, 9.14154e-19, 9.159283e-19, 9.152289e-19, 
    9.168929e-19, 9.179492e-19, 9.174269e-19, 9.206495e-19, 9.193971e-19, 
    9.259863e-19, 9.231504e-19, 9.305379e-19, 9.287721e-19, 9.30961e-19, 
    9.298445e-19, 9.317569e-19, 9.300358e-19, 9.330168e-19, 9.33665e-19, 
    9.332221e-19, 9.349244e-19, 9.299402e-19, 9.318554e-19, 9.174122e-19, 
    9.174974e-19, 9.178945e-19, 9.161484e-19, 9.160417e-19, 9.144413e-19, 
    9.158657e-19, 9.164718e-19, 9.180107e-19, 9.1892e-19, 9.197842e-19, 
    9.216834e-19, 9.23802e-19, 9.267623e-19, 9.288866e-19, 9.303098e-19, 
    9.294374e-19, 9.302076e-19, 9.293465e-19, 9.28943e-19, 9.33422e-19, 
    9.309077e-19, 9.346797e-19, 9.344712e-19, 9.327645e-19, 9.344947e-19, 
    9.175572e-19, 9.17067e-19, 9.153632e-19, 9.166967e-19, 9.14267e-19, 
    9.15627e-19, 9.164084e-19, 9.194227e-19, 9.200851e-19, 9.206983e-19, 
    9.219096e-19, 9.234628e-19, 9.261848e-19, 9.285507e-19, 9.307091e-19, 
    9.305511e-19, 9.306067e-19, 9.310884e-19, 9.298947e-19, 9.312843e-19, 
    9.315171e-19, 9.309078e-19, 9.344432e-19, 9.334338e-19, 9.344668e-19, 
    9.338096e-19, 9.172265e-19, 9.180514e-19, 9.176056e-19, 9.184436e-19, 
    9.17853e-19, 9.204772e-19, 9.212633e-19, 9.249394e-19, 9.234321e-19, 
    9.258312e-19, 9.236761e-19, 9.240579e-19, 9.259082e-19, 9.237928e-19, 
    9.284198e-19, 9.252829e-19, 9.311071e-19, 9.279771e-19, 9.31303e-19, 
    9.306998e-19, 9.316987e-19, 9.325928e-19, 9.337174e-19, 9.357905e-19, 
    9.353107e-19, 9.370437e-19, 9.192809e-19, 9.203496e-19, 9.20256e-19, 
    9.213744e-19, 9.22201e-19, 9.239923e-19, 9.268618e-19, 9.257832e-19, 
    9.277634e-19, 9.281604e-19, 9.251524e-19, 9.269993e-19, 9.21065e-19, 
    9.220242e-19, 9.214536e-19, 9.193648e-19, 9.260311e-19, 9.22612e-19, 
    9.289217e-19, 9.27073e-19, 9.324652e-19, 9.297843e-19, 9.350464e-19, 
    9.372909e-19, 9.394036e-19, 9.418671e-19, 9.209333e-19, 9.202072e-19, 
    9.215075e-19, 9.233043e-19, 9.249717e-19, 9.271857e-19, 9.274124e-19, 
    9.278268e-19, 9.288998e-19, 9.298019e-19, 9.279573e-19, 9.30028e-19, 
    9.222456e-19, 9.263279e-19, 9.199322e-19, 9.218593e-19, 9.231986e-19, 
    9.226117e-19, 9.256601e-19, 9.263778e-19, 9.292913e-19, 9.277862e-19, 
    9.367367e-19, 9.327808e-19, 9.437429e-19, 9.406846e-19, 9.199534e-19, 
    9.20931e-19, 9.243294e-19, 9.227131e-19, 9.273337e-19, 9.284689e-19, 
    9.293922e-19, 9.305711e-19, 9.306986e-19, 9.313969e-19, 9.302526e-19, 
    9.313519e-19, 9.271904e-19, 9.290508e-19, 9.239418e-19, 9.251861e-19, 
    9.24614e-19, 9.239858e-19, 9.25924e-19, 9.279862e-19, 9.280311e-19, 
    9.286913e-19, 9.305506e-19, 9.273524e-19, 9.372452e-19, 9.311389e-19, 
    9.219965e-19, 9.238763e-19, 9.241457e-19, 9.234176e-19, 9.283556e-19, 
    9.265675e-19, 9.3138e-19, 9.300804e-19, 9.322097e-19, 9.311517e-19, 
    9.30996e-19, 9.296367e-19, 9.287898e-19, 9.266493e-19, 9.249061e-19, 
    9.235233e-19, 9.238449e-19, 9.253637e-19, 9.281125e-19, 9.307099e-19, 
    9.301409e-19, 9.320479e-19, 9.26999e-19, 9.291167e-19, 9.282985e-19, 
    9.304324e-19, 9.257544e-19, 9.297359e-19, 9.247352e-19, 9.251742e-19, 
    9.265319e-19, 9.292598e-19, 9.298641e-19, 9.305079e-19, 9.301108e-19, 
    9.281824e-19, 9.278666e-19, 9.264992e-19, 9.261211e-19, 9.250788e-19, 
    9.24215e-19, 9.250039e-19, 9.25832e-19, 9.281835e-19, 9.302996e-19, 
    9.326053e-19, 9.331695e-19, 9.358579e-19, 9.336685e-19, 9.37279e-19, 
    9.34208e-19, 9.395222e-19, 9.299676e-19, 9.341193e-19, 9.26594e-19, 
    9.274062e-19, 9.288731e-19, 9.322368e-19, 9.304224e-19, 9.325446e-19, 
    9.278543e-19, 9.254157e-19, 9.247854e-19, 9.236072e-19, 9.248123e-19, 
    9.247144e-19, 9.258669e-19, 9.254967e-19, 9.282616e-19, 9.267768e-19, 
    9.309919e-19, 9.325281e-19, 9.368619e-19, 9.395139e-19, 9.422116e-19, 
    9.43401e-19, 9.43763e-19, 9.439143e-19 ;

 CWDN_TO_LITR3N =
  2.888338e-19, 2.896139e-19, 2.894624e-19, 2.90091e-19, 2.897424e-19, 
    2.901539e-19, 2.889921e-19, 2.896448e-19, 2.892283e-19, 2.889042e-19, 
    2.913092e-19, 2.901191e-19, 2.925444e-19, 2.917867e-19, 2.936887e-19, 
    2.924264e-19, 2.939431e-19, 2.936526e-19, 2.945271e-19, 2.942767e-19, 
    2.953936e-19, 2.946427e-19, 2.959723e-19, 2.952145e-19, 2.95333e-19, 
    2.946179e-19, 2.90359e-19, 2.91161e-19, 2.903114e-19, 2.904258e-19, 
    2.903745e-19, 2.897496e-19, 2.894343e-19, 2.887743e-19, 2.888942e-19, 
    2.89379e-19, 2.904773e-19, 2.901048e-19, 2.910437e-19, 2.910225e-19, 
    2.920662e-19, 2.915957e-19, 2.933477e-19, 2.928504e-19, 2.942872e-19, 
    2.93926e-19, 2.942702e-19, 2.941659e-19, 2.942715e-19, 2.937418e-19, 
    2.939688e-19, 2.935026e-19, 2.916838e-19, 2.922188e-19, 2.90622e-19, 
    2.896598e-19, 2.890207e-19, 2.885667e-19, 2.886309e-19, 2.887532e-19, 
    2.893818e-19, 2.899726e-19, 2.904225e-19, 2.907232e-19, 2.910194e-19, 
    2.919147e-19, 2.923886e-19, 2.934482e-19, 2.932573e-19, 2.935808e-19, 
    2.938901e-19, 2.944088e-19, 2.943235e-19, 2.945518e-19, 2.935724e-19, 
    2.942234e-19, 2.931486e-19, 2.934426e-19, 2.910991e-19, 2.902054e-19, 
    2.898244e-19, 2.894915e-19, 2.886802e-19, 2.892405e-19, 2.890197e-19, 
    2.895451e-19, 2.898787e-19, 2.897138e-19, 2.907314e-19, 2.903359e-19, 
    2.924167e-19, 2.915212e-19, 2.938541e-19, 2.932965e-19, 2.939877e-19, 
    2.936351e-19, 2.94239e-19, 2.936955e-19, 2.946369e-19, 2.948416e-19, 
    2.947017e-19, 2.952393e-19, 2.936654e-19, 2.942701e-19, 2.897091e-19, 
    2.89736e-19, 2.898614e-19, 2.8931e-19, 2.892764e-19, 2.887709e-19, 
    2.892208e-19, 2.894121e-19, 2.898981e-19, 2.901852e-19, 2.904582e-19, 
    2.910579e-19, 2.91727e-19, 2.926618e-19, 2.933326e-19, 2.93782e-19, 
    2.935066e-19, 2.937497e-19, 2.934778e-19, 2.933504e-19, 2.947649e-19, 
    2.939709e-19, 2.95162e-19, 2.950962e-19, 2.945572e-19, 2.951036e-19, 
    2.897549e-19, 2.896001e-19, 2.890621e-19, 2.894832e-19, 2.887159e-19, 
    2.891454e-19, 2.893921e-19, 2.90344e-19, 2.905532e-19, 2.907468e-19, 
    2.911293e-19, 2.916198e-19, 2.924794e-19, 2.932265e-19, 2.939082e-19, 
    2.938582e-19, 2.938758e-19, 2.940279e-19, 2.93651e-19, 2.940898e-19, 
    2.941633e-19, 2.939709e-19, 2.950873e-19, 2.947686e-19, 2.950948e-19, 
    2.948873e-19, 2.896504e-19, 2.89911e-19, 2.897702e-19, 2.900348e-19, 
    2.898483e-19, 2.90677e-19, 2.909253e-19, 2.920861e-19, 2.916101e-19, 
    2.923678e-19, 2.916872e-19, 2.918078e-19, 2.923921e-19, 2.91724e-19, 
    2.931852e-19, 2.921946e-19, 2.940338e-19, 2.930454e-19, 2.940957e-19, 
    2.939052e-19, 2.942206e-19, 2.94503e-19, 2.948581e-19, 2.955128e-19, 
    2.953613e-19, 2.959085e-19, 2.902992e-19, 2.906367e-19, 2.906072e-19, 
    2.909603e-19, 2.912214e-19, 2.91787e-19, 2.926932e-19, 2.923526e-19, 
    2.929779e-19, 2.931033e-19, 2.921534e-19, 2.927366e-19, 2.908626e-19, 
    2.911656e-19, 2.909853e-19, 2.903257e-19, 2.924309e-19, 2.913512e-19, 
    2.933437e-19, 2.927599e-19, 2.944627e-19, 2.936161e-19, 2.952778e-19, 
    2.959866e-19, 2.966538e-19, 2.974317e-19, 2.90821e-19, 2.905918e-19, 
    2.910024e-19, 2.915698e-19, 2.920963e-19, 2.927955e-19, 2.928671e-19, 
    2.929979e-19, 2.933368e-19, 2.936216e-19, 2.930391e-19, 2.93693e-19, 
    2.912355e-19, 2.925246e-19, 2.905049e-19, 2.911134e-19, 2.915364e-19, 
    2.913511e-19, 2.923137e-19, 2.925404e-19, 2.934604e-19, 2.929851e-19, 
    2.958116e-19, 2.945624e-19, 2.98024e-19, 2.970583e-19, 2.905116e-19, 
    2.908203e-19, 2.918935e-19, 2.913831e-19, 2.928422e-19, 2.932007e-19, 
    2.934923e-19, 2.938645e-19, 2.939048e-19, 2.941253e-19, 2.93764e-19, 
    2.941111e-19, 2.92797e-19, 2.933845e-19, 2.917711e-19, 2.92164e-19, 
    2.919834e-19, 2.91785e-19, 2.92397e-19, 2.930483e-19, 2.930624e-19, 
    2.932709e-19, 2.938581e-19, 2.928481e-19, 2.959722e-19, 2.940439e-19, 
    2.911568e-19, 2.917504e-19, 2.918355e-19, 2.916056e-19, 2.931649e-19, 
    2.926003e-19, 2.9412e-19, 2.937096e-19, 2.94382e-19, 2.940479e-19, 
    2.939988e-19, 2.935695e-19, 2.93302e-19, 2.926261e-19, 2.920756e-19, 
    2.916389e-19, 2.917405e-19, 2.922201e-19, 2.930881e-19, 2.939084e-19, 
    2.937287e-19, 2.943309e-19, 2.927365e-19, 2.934053e-19, 2.931469e-19, 
    2.938207e-19, 2.923435e-19, 2.936008e-19, 2.920216e-19, 2.921603e-19, 
    2.92589e-19, 2.934504e-19, 2.936413e-19, 2.938446e-19, 2.937192e-19, 
    2.931102e-19, 2.930105e-19, 2.925787e-19, 2.924593e-19, 2.921301e-19, 
    2.918574e-19, 2.921065e-19, 2.92368e-19, 2.931106e-19, 2.937788e-19, 
    2.94507e-19, 2.946851e-19, 2.955341e-19, 2.948427e-19, 2.959828e-19, 
    2.950131e-19, 2.966912e-19, 2.93674e-19, 2.949851e-19, 2.926086e-19, 
    2.928651e-19, 2.933283e-19, 2.943906e-19, 2.938176e-19, 2.944878e-19, 
    2.930066e-19, 2.922365e-19, 2.920375e-19, 2.916654e-19, 2.92046e-19, 
    2.920151e-19, 2.92379e-19, 2.922621e-19, 2.931352e-19, 2.926664e-19, 
    2.939974e-19, 2.944826e-19, 2.958511e-19, 2.966886e-19, 2.975405e-19, 
    2.979161e-19, 2.980304e-19, 2.980782e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  2.809604e-14, 2.822128e-14, 2.819686e-14, 2.829796e-14, 2.824182e-14, 
    2.830801e-14, 2.812127e-14, 2.822611e-14, 2.815912e-14, 2.810706e-14, 
    2.849423e-14, 2.830228e-14, 2.869358e-14, 2.857098e-14, 2.88789e-14, 
    2.867447e-14, 2.892011e-14, 2.887287e-14, 2.901481e-14, 2.897409e-14, 
    2.915586e-14, 2.903352e-14, 2.925002e-14, 2.912656e-14, 2.914586e-14, 
    2.902938e-14, 2.8341e-14, 2.847052e-14, 2.83333e-14, 2.835176e-14, 
    2.834343e-14, 2.82429e-14, 2.81923e-14, 2.80862e-14, 2.810541e-14, 
    2.81833e-14, 2.835988e-14, 2.829983e-14, 2.845097e-14, 2.844756e-14, 
    2.861602e-14, 2.854003e-14, 2.882342e-14, 2.874277e-14, 2.897576e-14, 
    2.891711e-14, 2.897297e-14, 2.895598e-14, 2.897312e-14, 2.888716e-14, 
    2.892394e-14, 2.88483e-14, 2.855456e-14, 2.864098e-14, 2.838328e-14, 
    2.822859e-14, 2.812577e-14, 2.805293e-14, 2.806317e-14, 2.808282e-14, 
    2.81837e-14, 2.827855e-14, 2.835091e-14, 2.83993e-14, 2.8447e-14, 
    2.859172e-14, 2.86682e-14, 2.88397e-14, 2.880867e-14, 2.886115e-14, 
    2.891125e-14, 2.899544e-14, 2.898155e-14, 2.901864e-14, 2.885959e-14, 
    2.896528e-14, 2.87908e-14, 2.88385e-14, 2.846044e-14, 2.831612e-14, 
    2.8255e-14, 2.820134e-14, 2.807108e-14, 2.816101e-14, 2.812553e-14, 
    2.820981e-14, 2.826342e-14, 2.823685e-14, 2.84006e-14, 2.833688e-14, 
    2.86727e-14, 2.852796e-14, 2.890543e-14, 2.881498e-14, 2.892703e-14, 
    2.886982e-14, 2.896783e-14, 2.887958e-14, 2.90324e-14, 2.906573e-14, 
    2.90429e-14, 2.913032e-14, 2.887454e-14, 2.897274e-14, 2.823626e-14, 
    2.82406e-14, 2.826071e-14, 2.817215e-14, 2.816671e-14, 2.808554e-14, 
    2.815768e-14, 2.818845e-14, 2.826645e-14, 2.831263e-14, 2.835653e-14, 
    2.845316e-14, 2.856115e-14, 2.871222e-14, 2.882081e-14, 2.889362e-14, 
    2.884892e-14, 2.888834e-14, 2.884423e-14, 2.882352e-14, 2.905318e-14, 
    2.89242e-14, 2.911768e-14, 2.910696e-14, 2.901934e-14, 2.91081e-14, 
    2.824358e-14, 2.821864e-14, 2.813227e-14, 2.819981e-14, 2.807665e-14, 
    2.814559e-14, 2.818523e-14, 2.833823e-14, 2.837179e-14, 2.840301e-14, 
    2.846461e-14, 2.854373e-14, 2.868267e-14, 2.88036e-14, 2.891405e-14, 
    2.890591e-14, 2.890875e-14, 2.893342e-14, 2.887225e-14, 2.894341e-14, 
    2.895535e-14, 2.892409e-14, 2.910545e-14, 2.905361e-14, 2.910663e-14, 
    2.907283e-14, 2.82267e-14, 2.826856e-14, 2.824589e-14, 2.828848e-14, 
    2.825844e-14, 2.839187e-14, 2.843186e-14, 2.861918e-14, 2.854218e-14, 
    2.866464e-14, 2.855455e-14, 2.857406e-14, 2.866864e-14, 2.856042e-14, 
    2.879689e-14, 2.863656e-14, 2.893435e-14, 2.877422e-14, 2.894435e-14, 
    2.891337e-14, 2.896455e-14, 2.901045e-14, 2.906811e-14, 2.917472e-14, 
    2.914996e-14, 2.923912e-14, 2.833099e-14, 2.838535e-14, 2.838051e-14, 
    2.843739e-14, 2.847947e-14, 2.857074e-14, 2.871724e-14, 2.866207e-14, 
    2.876322e-14, 2.878356e-14, 2.862977e-14, 2.872418e-14, 2.842148e-14, 
    2.847035e-14, 2.844119e-14, 2.833492e-14, 2.867462e-14, 2.850018e-14, 
    2.882232e-14, 2.872769e-14, 2.900383e-14, 2.886648e-14, 2.913636e-14, 
    2.925198e-14, 2.936063e-14, 2.948788e-14, 2.841497e-14, 2.837797e-14, 
    2.844409e-14, 2.853575e-14, 2.862067e-14, 2.873376e-14, 2.874528e-14, 
    2.876645e-14, 2.882132e-14, 2.886751e-14, 2.877314e-14, 2.887902e-14, 
    2.848174e-14, 2.868974e-14, 2.836371e-14, 2.846187e-14, 2.852998e-14, 
    2.850004e-14, 2.865544e-14, 2.869207e-14, 2.884114e-14, 2.876403e-14, 
    2.92234e-14, 2.902002e-14, 2.958466e-14, 2.942673e-14, 2.836504e-14, 
    2.841472e-14, 2.858792e-14, 2.850547e-14, 2.874122e-14, 2.879934e-14, 
    2.88465e-14, 2.890694e-14, 2.891339e-14, 2.894921e-14, 2.889047e-14, 
    2.894683e-14, 2.873374e-14, 2.882891e-14, 2.856779e-14, 2.863129e-14, 
    2.860203e-14, 2.856995e-14, 2.866884e-14, 2.877435e-14, 2.877651e-14, 
    2.881033e-14, 2.890587e-14, 2.874172e-14, 2.924969e-14, 2.893589e-14, 
    2.846894e-14, 2.856483e-14, 2.857843e-14, 2.854128e-14, 2.879344e-14, 
    2.870203e-14, 2.894833e-14, 2.888167e-14, 2.899079e-14, 2.893655e-14, 
    2.892852e-14, 2.885887e-14, 2.881548e-14, 2.870603e-14, 2.861695e-14, 
    2.854637e-14, 2.856272e-14, 2.864028e-14, 2.878072e-14, 2.89137e-14, 
    2.888454e-14, 2.898217e-14, 2.872361e-14, 2.883201e-14, 2.879007e-14, 
    2.889929e-14, 2.866052e-14, 2.886447e-14, 2.860843e-14, 2.86308e-14, 
    2.870014e-14, 2.883978e-14, 2.887054e-14, 2.890357e-14, 2.888313e-14, 
    2.878446e-14, 2.876824e-14, 2.869827e-14, 2.867897e-14, 2.86257e-14, 
    2.858157e-14, 2.862186e-14, 2.866412e-14, 2.878428e-14, 2.889263e-14, 
    2.90108e-14, 2.903971e-14, 2.917806e-14, 2.906547e-14, 2.925133e-14, 
    2.90934e-14, 2.936673e-14, 2.887613e-14, 2.908913e-14, 2.870328e-14, 
    2.874475e-14, 2.881992e-14, 2.899227e-14, 2.889908e-14, 2.900801e-14, 
    2.876758e-14, 2.864303e-14, 2.861071e-14, 2.855063e-14, 2.861204e-14, 
    2.860704e-14, 2.866584e-14, 2.864689e-14, 2.87882e-14, 2.871227e-14, 
    2.8928e-14, 2.900684e-14, 2.922951e-14, 2.936615e-14, 2.950526e-14, 
    2.95667e-14, 2.95854e-14, 2.95932e-14 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  6.531128, 6.547447, 6.544277, 6.557425, 6.550149, 6.558741, 6.534445, 
    6.548085, 6.539382, 6.532613, 6.582907, 6.558012, 6.608951, 6.592999, 
    6.634775, 6.606448, 6.64019, 6.63403, 6.652662, 6.64732, 6.671146, 
    6.655128, 6.683582, 6.667334, 6.669861, 6.654596, 6.563043, 6.579797, 
    6.562045, 6.564433, 6.563368, 6.55029, 6.543667, 6.529902, 6.532404, 
    6.542525, 6.565508, 6.557729, 6.577405, 6.576961, 6.598885, 6.58899, 
    6.627558, 6.615445, 6.647544, 6.639848, 6.647177, 6.644958, 6.647206, 
    6.635925, 6.640754, 6.630847, 6.590837, 6.602097, 6.568547, 6.548378, 
    6.535038, 6.525569, 6.526907, 6.529452, 6.542583, 6.554966, 6.564379, 
    6.570679, 6.576897, 6.595653, 6.605663, 6.629677, 6.625644, 6.632495, 
    6.639084, 6.65013, 6.648314, 6.653179, 6.632332, 6.64617, 6.621759, 
    6.629574, 6.578494, 6.559831, 6.551834, 6.544883, 6.527934, 6.539629, 
    6.535013, 6.546019, 6.553003, 6.549554, 6.570852, 6.562563, 6.606257, 
    6.58741, 6.638316, 6.626473, 6.641162, 6.633666, 6.646506, 6.634949, 
    6.654998, 6.65936, 6.656377, 6.667881, 6.634306, 6.647167, 6.549453, 
    6.550015, 6.552646, 6.541081, 6.54038, 6.529829, 6.539225, 6.543223, 
    6.553414, 6.55941, 6.565121, 6.577697, 6.591733, 6.611441, 6.627239, 
    6.636789, 6.630938, 6.636103, 6.630326, 6.627625, 6.657719, 6.640793, 
    6.666224, 6.664818, 6.65329, 6.664977, 6.550412, 6.547172, 6.535905, 
    6.544721, 6.528682, 6.537643, 6.542794, 6.562717, 6.567115, 6.571168, 
    6.579199, 6.589495, 6.607593, 6.624981, 6.639472, 6.638411, 6.638783, 
    6.642015, 6.633999, 6.643333, 6.644891, 6.640803, 6.664629, 6.657815, 
    6.664788, 6.660352, 6.548227, 6.553678, 6.550734, 6.556261, 6.552363, 
    6.569687, 6.57489, 6.599286, 6.589287, 6.605234, 6.590912, 6.593442, 
    6.605714, 6.591691, 6.624088, 6.601563, 6.642142, 6.619524, 6.64346, 
    6.639409, 6.646127, 6.652138, 6.659727, 6.673724, 6.670484, 6.682224, 
    6.561796, 6.568852, 6.568248, 6.575653, 6.581124, 6.593015, 6.612114, 
    6.604932, 6.618143, 6.620792, 6.600734, 6.613024, 6.573592, 6.579934, 
    6.576172, 6.562342, 6.606562, 6.583831, 6.627471, 6.613527, 6.651278, 
    6.633239, 6.668697, 6.683864, 6.698265, 6.715024, 6.572726, 6.567925, 
    6.576539, 6.588424, 6.599522, 6.614276, 6.615798, 6.618561, 6.627335, 
    6.633379, 6.619417, 6.634898, 6.581368, 6.608547, 6.566095, 6.578838, 
    6.587731, 6.583847, 6.604116, 6.608896, 6.629941, 6.618296, 6.6801, 
    6.653381, 6.727882, 6.706962, 6.566245, 6.572717, 6.595241, 6.584521, 
    6.615273, 6.624441, 6.630635, 6.638532, 6.6394, 6.644087, 6.636405, 
    6.643791, 6.614307, 6.628342, 6.592684, 6.60095, 6.597152, 6.592976, 
    6.605871, 6.619607, 6.619931, 6.625923, 6.638312, 6.615397, 6.683498, 
    6.642277, 6.579777, 6.592217, 6.594031, 6.589201, 6.622095, 6.610153, 
    6.643977, 6.635249, 6.649565, 6.642444, 6.641396, 6.632272, 6.626592, 
    6.610694, 6.599084, 6.589905, 6.59204, 6.602128, 6.620455, 6.639465, 
    6.635638, 6.648476, 6.613036, 6.628772, 6.621701, 6.637608, 6.604734, 
    6.632859, 6.597959, 6.600879, 6.609917, 6.629714, 6.633797, 6.638107, 
    6.635454, 6.620926, 6.618824, 6.609704, 6.607174, 6.600245, 6.5945, 
    6.599741, 6.605244, 6.620944, 6.636707, 6.652219, 6.656033, 6.674136, 
    6.659352, 6.683722, 6.662931, 6.698997, 6.634445, 6.662386, 6.610338, 
    6.615758, 6.627128, 6.649713, 6.63754, 6.651793, 6.618744, 6.602461, 
    6.598291, 6.590457, 6.59847, 6.597819, 6.605494, 6.603028, 6.621467, 
    6.611557, 6.641361, 6.651688, 6.680981, 6.698986, 6.717416, 6.725552, 
    6.728033, 6.729068 ;

 EFLX_LH_TOT_R =
  6.531128, 6.547447, 6.544277, 6.557425, 6.550149, 6.558741, 6.534445, 
    6.548085, 6.539382, 6.532613, 6.582907, 6.558012, 6.608951, 6.592999, 
    6.634775, 6.606448, 6.64019, 6.63403, 6.652662, 6.64732, 6.671146, 
    6.655128, 6.683582, 6.667334, 6.669861, 6.654596, 6.563043, 6.579797, 
    6.562045, 6.564433, 6.563368, 6.55029, 6.543667, 6.529902, 6.532404, 
    6.542525, 6.565508, 6.557729, 6.577405, 6.576961, 6.598885, 6.58899, 
    6.627558, 6.615445, 6.647544, 6.639848, 6.647177, 6.644958, 6.647206, 
    6.635925, 6.640754, 6.630847, 6.590837, 6.602097, 6.568547, 6.548378, 
    6.535038, 6.525569, 6.526907, 6.529452, 6.542583, 6.554966, 6.564379, 
    6.570679, 6.576897, 6.595653, 6.605663, 6.629677, 6.625644, 6.632495, 
    6.639084, 6.65013, 6.648314, 6.653179, 6.632332, 6.64617, 6.621759, 
    6.629574, 6.578494, 6.559831, 6.551834, 6.544883, 6.527934, 6.539629, 
    6.535013, 6.546019, 6.553003, 6.549554, 6.570852, 6.562563, 6.606257, 
    6.58741, 6.638316, 6.626473, 6.641162, 6.633666, 6.646506, 6.634949, 
    6.654998, 6.65936, 6.656377, 6.667881, 6.634306, 6.647167, 6.549453, 
    6.550015, 6.552646, 6.541081, 6.54038, 6.529829, 6.539225, 6.543223, 
    6.553414, 6.55941, 6.565121, 6.577697, 6.591733, 6.611441, 6.627239, 
    6.636789, 6.630938, 6.636103, 6.630326, 6.627625, 6.657719, 6.640793, 
    6.666224, 6.664818, 6.65329, 6.664977, 6.550412, 6.547172, 6.535905, 
    6.544721, 6.528682, 6.537643, 6.542794, 6.562717, 6.567115, 6.571168, 
    6.579199, 6.589495, 6.607593, 6.624981, 6.639472, 6.638411, 6.638783, 
    6.642015, 6.633999, 6.643333, 6.644891, 6.640803, 6.664629, 6.657815, 
    6.664788, 6.660352, 6.548227, 6.553678, 6.550734, 6.556261, 6.552363, 
    6.569687, 6.57489, 6.599286, 6.589287, 6.605234, 6.590912, 6.593442, 
    6.605714, 6.591691, 6.624088, 6.601563, 6.642142, 6.619524, 6.64346, 
    6.639409, 6.646127, 6.652138, 6.659727, 6.673724, 6.670484, 6.682224, 
    6.561796, 6.568852, 6.568248, 6.575653, 6.581124, 6.593015, 6.612114, 
    6.604932, 6.618143, 6.620792, 6.600734, 6.613024, 6.573592, 6.579934, 
    6.576172, 6.562342, 6.606562, 6.583831, 6.627471, 6.613527, 6.651278, 
    6.633239, 6.668697, 6.683864, 6.698265, 6.715024, 6.572726, 6.567925, 
    6.576539, 6.588424, 6.599522, 6.614276, 6.615798, 6.618561, 6.627335, 
    6.633379, 6.619417, 6.634898, 6.581368, 6.608547, 6.566095, 6.578838, 
    6.587731, 6.583847, 6.604116, 6.608896, 6.629941, 6.618296, 6.6801, 
    6.653381, 6.727882, 6.706962, 6.566245, 6.572717, 6.595241, 6.584521, 
    6.615273, 6.624441, 6.630635, 6.638532, 6.6394, 6.644087, 6.636405, 
    6.643791, 6.614307, 6.628342, 6.592684, 6.60095, 6.597152, 6.592976, 
    6.605871, 6.619607, 6.619931, 6.625923, 6.638312, 6.615397, 6.683498, 
    6.642277, 6.579777, 6.592217, 6.594031, 6.589201, 6.622095, 6.610153, 
    6.643977, 6.635249, 6.649565, 6.642444, 6.641396, 6.632272, 6.626592, 
    6.610694, 6.599084, 6.589905, 6.59204, 6.602128, 6.620455, 6.639465, 
    6.635638, 6.648476, 6.613036, 6.628772, 6.621701, 6.637608, 6.604734, 
    6.632859, 6.597959, 6.600879, 6.609917, 6.629714, 6.633797, 6.638107, 
    6.635454, 6.620926, 6.618824, 6.609704, 6.607174, 6.600245, 6.5945, 
    6.599741, 6.605244, 6.620944, 6.636707, 6.652219, 6.656033, 6.674136, 
    6.659352, 6.683722, 6.662931, 6.698997, 6.634445, 6.662386, 6.610338, 
    6.615758, 6.627128, 6.649713, 6.63754, 6.651793, 6.618744, 6.602461, 
    6.598291, 6.590457, 6.59847, 6.597819, 6.605494, 6.603028, 6.621467, 
    6.611557, 6.641361, 6.651688, 6.680981, 6.698986, 6.717416, 6.725552, 
    6.728033, 6.729068 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371698e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441075e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379093e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377207e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523353e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.56315e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529406e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.532169e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547246e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.46224e-08, 6.465288e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532766e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472856e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRSEB =
  -6.253161e-15, -1.553191e-14, -1.131726e-14, 2.712503e-15, -1.487663e-15, 
    -1.81218e-14, -7.820266e-15, -4.416874e-15, 9.396942e-16, -9.224797e-15, 
    -1.651936e-14, -3.697176e-15, -7.343926e-15, -8.668344e-15, 
    -1.381564e-14, -4.52826e-15, -1.121069e-15, -7.544976e-15, -4.216774e-15, 
    -1.136348e-14, -3.639895e-15, -1.250076e-14, -3.072584e-15, 
    -1.148642e-15, -3.553257e-15, -8.177055e-18, -1.654158e-14, 
    -1.158891e-14, -6.638382e-15, -1.304099e-14, -4.495705e-15, 
    -4.051431e-15, -1.154651e-14, -1.297752e-14, -1.674446e-14, 
    -4.036189e-15, -1.326929e-14, -1.460674e-14, -2.268408e-15, 
    -3.739606e-15, -1.834292e-14, -8.073438e-15, -4.391388e-15, 2.207524e-15, 
    -2.469389e-15, -1.607202e-14, -3.29813e-15, -9.449302e-15, -1.185917e-14, 
    -7.891191e-15, -1.095381e-14, -8.831358e-15, -7.592978e-15, 
    -1.545608e-14, -1.596736e-14, -1.102812e-14, -1.06755e-14, -1.414296e-14, 
    -8.053845e-15, 4.916204e-15, -1.819847e-14, -1.027414e-14, -1.579538e-15, 
    -9.120188e-15, -6.195468e-15, -2.778516e-15, -6.521608e-16, 
    -1.095961e-14, -8.126923e-15, -1.832852e-14, -9.730378e-16, 
    -9.107361e-15, -6.675286e-15, -6.110429e-15, -3.61843e-15, -1.683952e-14, 
    -6.768975e-15, -2.10034e-15, -2.271991e-14, -1.021729e-14, -1.048557e-14, 
    -1.116528e-14, -2.648113e-15, -1.197956e-14, -6.189682e-15, 
    -5.468605e-15, -4.622675e-15, -5.644731e-15, -8.126547e-15, 
    -8.202248e-15, -4.67631e-15, -1.216326e-14, -2.968904e-15, -3.803049e-15, 
    -8.886355e-15, -6.989818e-15, -8.88481e-15, -1.627541e-14, -6.515737e-15, 
    -1.172322e-15, -1.411588e-14, -1.025841e-14, -9.549709e-15, 
    -1.310095e-14, 2.304777e-15, -4.312879e-15, -1.255311e-14, -1.057639e-14, 
    -1.865242e-14, -4.966483e-15, -8.726252e-15, -1.356977e-14, 
    -1.041762e-14, -8.528809e-15, -1.393112e-14, -4.27783e-15, 1.044454e-16, 
    -8.699055e-15, -3.983469e-15, -9.796853e-15, -2.680628e-15, 
    -9.146635e-15, -1.212463e-14, -6.609626e-15, -7.280891e-15, -1.14109e-14, 
    -8.296778e-15, -9.154156e-15, -5.49142e-15, 2.796892e-15, -1.05701e-14, 
    -4.614876e-15, -5.730083e-15, -2.3988e-15, -8.326622e-15, -3.598409e-15, 
    -9.486214e-15, -2.240083e-15, -1.724124e-14, 4.414643e-15, -7.805861e-15, 
    -1.53877e-14, -9.936718e-15, -1.807631e-14, -1.441534e-14, -1.246955e-14, 
    -3.550641e-15, -1.326267e-14, -5.277666e-15, -5.114171e-15, 
    -4.907365e-15, -9.372885e-15, -3.302205e-16, -1.899493e-15, 
    -8.029791e-16, -1.354811e-14, -9.738074e-15, -6.565266e-15, -1.23684e-14, 
    -1.383411e-14, -1.357697e-14, -1.517481e-14, -8.957373e-15, 
    -4.715903e-15, -4.547141e-15, -1.811438e-14, -1.265612e-14, 
    -1.640331e-14, -2.90959e-15, -5.169011e-15, -1.596064e-14, -1.141599e-14, 
    -7.218749e-15, -2.424933e-15, -6.699321e-15, -1.079221e-14, 
    -6.057789e-15, -3.722356e-16, -1.486633e-14, -2.103712e-14, 
    -8.106033e-15, -8.057749e-15, -7.57973e-15, -1.251528e-14, -4.294976e-15, 
    -2.833555e-15, -9.215005e-15, -1.243491e-14, -1.368951e-15, 
    -1.808665e-15, -6.926151e-15, -8.727122e-15, -1.075766e-14, 
    -8.085985e-15, -5.213762e-15, -1.124694e-14, -8.450777e-15, 
    -4.870672e-15, -1.163313e-14, -7.48031e-15, -8.996749e-15, -7.954369e-15, 
    -3.909571e-15, -9.978624e-15, -7.748619e-15, -4.176187e-15, 
    -1.104897e-14, -1.450791e-14, -9.895406e-15, -9.25823e-15, -1.54121e-14, 
    -8.594477e-15, -1.281552e-14, -5.665371e-15, -7.612801e-15, 
    -1.053351e-14, -1.084867e-14, -1.447422e-15, -1.498358e-14, 
    -1.521876e-14, -1.275265e-14, -6.84949e-15, -1.206105e-14, -3.789708e-15, 
    -1.336663e-14, -1.226966e-14, -9.755463e-15, -1.596606e-14, 
    -9.217696e-15, -9.923532e-15, -8.091169e-16, -2.062669e-14, 
    -1.907824e-14, -1.520397e-14, -1.088743e-14, -9.99849e-15, -1.470407e-14, 
    -1.040991e-14, -1.175404e-14, -6.031384e-15, -2.0699e-15, -1.009195e-15, 
    4.483923e-15, -8.775565e-15, -1.320182e-14, -1.085643e-14, -5.323367e-15, 
    -8.279515e-15, -1.61334e-14, -1.673462e-14, 1.490803e-15, -1.00047e-14, 
    -9.486221e-15, -1.397551e-14, -3.547385e-15, -6.518539e-15, 
    -7.442845e-15, -9.1902e-15, -1.118584e-14, -1.483589e-14, -1.622965e-14, 
    -9.254132e-15, -8.646704e-15, -1.381016e-14, -1.147194e-14, -3.94859e-15, 
    -3.630855e-15, -1.861975e-14, -9.746882e-15, -4.013426e-15, 
    -5.368026e-15, -1.386825e-14, -1.244192e-14, -4.175092e-15, 
    -7.166103e-15, -1.164187e-14, -2.068687e-15, -1.025228e-14, 
    -9.182051e-15, -1.02617e-14, -7.671859e-16, -1.042099e-14, -1.761199e-14, 
    -8.813181e-15, 1.409223e-15, -1.860168e-14, 4.855328e-15, -6.174119e-15, 
    -1.067627e-14, -1.463606e-14, -1.103473e-14, -1.157287e-14, 
    -4.504936e-15, -2.286842e-15, -6.444776e-15, -1.094942e-14, 
    -1.070439e-14, -6.110848e-15, -4.900457e-15, -7.940894e-15, 
    -6.917319e-15, -6.806471e-15, 6.751981e-15, 3.629188e-15, -2.92161e-15, 
    -8.984932e-15, -2.281e-14, -1.206147e-14, -9.343113e-15, -1.150389e-14, 
    -7.380786e-15, -1.840556e-14, -7.039468e-15, -3.321711e-15, -1.73534e-14, 
    -9.434207e-15, -1.034618e-14, -1.368323e-14, -4.54852e-15, -9.620026e-15, 
    -1.626562e-14, -1.636982e-14, -1.222475e-14, -4.112137e-15, 
    -3.541481e-15, -3.608429e-15, -4.327759e-15, -8.500582e-15, 
    -1.950778e-14, -1.757483e-14, -1.726668e-15, -1.284552e-15, 
    -3.085501e-15, -1.942044e-14, -9.303465e-15, -2.421472e-15, 
    -4.605947e-15, -6.884782e-15 ;

 ERRSOI =
  -71.27113, -71.36424, -71.34656, -71.42079, -71.38028, -71.4284, -71.2908, 
    -71.36723, -71.31889, -71.28061, -71.56287, -71.4243, -71.71505, 
    -71.62503, -71.85405, -71.69992, -71.88551, -71.85145, -71.95857, 
    -71.92797, -72.06138, -71.97272, -72.13376, -72.04118, -72.05495, 
    -71.96949, -71.45391, -71.54501, -71.4481, -71.46118, -71.45573, 
    -71.38047, -71.34142, -71.26527, -71.27942, -71.33604, -71.46711, 
    -71.42377, -71.53664, -71.53413, -71.65892, -71.60257, -71.81436, 
    -71.7544, -71.92928, -71.88497, -71.92688, -71.91441, -71.92704, 
    -71.86218, -71.88986, -71.83343, -71.61278, -71.6769, -71.48499, 
    -71.36727, -71.29382, -71.24039, -71.24794, -71.26196, -71.33633, 
    -71.40796, -71.46207, -71.49802, -71.53374, -71.63728, -71.69622, 
    -71.82558, -71.80378, -71.84192, -71.88065, -71.9436, -71.93346, 
    -71.96085, -71.84206, -71.9204, -71.7909, -71.82615, -71.53722, 
    -71.43575, -71.38734, -71.34972, -71.25361, -71.31963, -71.29344, 
    -71.35708, -71.39665, -71.37733, -71.49902, -71.45142, -71.69971, 
    -71.59263, -71.87614, -71.80838, -71.89262, -71.84992, -71.92259, 
    -71.8572, -71.97156, -71.99578, -71.97909, -72.04538, -71.85341, 
    -71.92628, -71.3765, -71.3796, -71.39484, -71.32779, -71.32405, 
    -71.26457, -71.31805, -71.34034, -71.39944, -71.43327, -71.46587, 
    -71.53774, -71.61711, -71.73019, -71.8127, -71.86777, -71.8344, 
    -71.86381, -71.8307, -71.81547, -71.9863, -71.88973, -72.03583, 
    -72.02795, -71.96126, -72.02885, -71.3819, -71.36378, -71.29896, 
    -71.3497, -71.25819, -71.3086, -71.33715, -71.45107, -71.47762, 
    -71.50032, -71.54665, -71.60542, -71.70834, -71.79922, -71.88316, 
    -71.87713, -71.8792, -71.89732, -71.85156, -71.9049, -71.91325, 
    -71.89046, -72.02686, -71.98792, -72.02777, -72.00257, -71.36983, 
    -71.4006, -71.38387, -71.41499, -71.39256, -71.49059, -71.52, -71.65977, 
    -71.60391, -71.69457, -71.61361, -71.62759, -71.69489, -71.61839, 
    -71.79301, -71.67213, -71.89804, -71.7745, -71.90564, -71.88279, 
    -71.92125, -71.95504, -71.99876, -72.07774, -72.05968, -72.12685, 
    -71.4471, -71.48653, -71.48421, -71.52635, -71.55727, -71.62586, 
    -71.73473, -71.69412, -71.76999, -71.78481, -71.67029, -71.73944, 
    -71.51383, -71.54897, -71.52892, -71.44952, -71.70186, -71.57143, 
    -71.81384, -71.74308, -71.95007, -71.84581, -72.04948, -72.1338, 
    -72.21884, -72.31203, -71.50935, -71.4824, -71.5317, -71.59785, 
    -71.66268, -71.74718, -71.75648, -71.77197, -71.81373, -71.84819, 
    -71.77573, -71.85696, -71.55476, -71.71375, -71.47113, -71.54245, 
    -71.59447, -71.57283, -71.68979, -71.71698, -71.82738, -71.7709, 
    -72.11193, -71.96052, -72.38713, -72.26662, -71.4727, -71.5098, 
    -71.63747, -71.57686, -71.75345, -71.79661, -71.83268, -71.87691, 
    -71.88255, -71.90894, -71.86557, -71.90769, -71.74734, -71.81915, 
    -71.62426, -71.67089, -71.64984, -71.62589, -71.6997, -71.77658, 
    -71.78012, -71.80458, -71.86993, -71.75419, -72.12801, -71.89344, 
    -71.55017, -71.61921, -71.63139, -71.60421, -71.79212, -71.72368, 
    -71.90857, -71.85894, -71.94079, -71.89993, -71.89383, -71.84187, 
    -71.80904, -71.72646, -71.66003, -71.60838, -71.62053, -71.67732, 
    -71.78172, -71.88222, -71.85993, -71.93459, -71.74053, -71.82085, 
    -71.7891, -71.87213, -71.69262, -71.83971, -71.65449, -71.67107, 
    -71.72234, -71.82504, -71.85059, -71.87447, -71.86013, -71.78473, 
    -71.77326, -71.72156, -71.70636, -71.6676, -71.63465, -71.66428, 
    -71.69502, -71.78555, -71.86636, -71.95525, -71.97775, -72.07717, 
    -71.9936, -72.12894, -72.00988, -72.21819, -71.85103, -72.01026, 
    -71.72531, -71.75636, -71.81062, -71.93929, -71.87177, -71.95166, 
    -71.77296, -71.67833, -71.65625, -71.61117, -71.65728, -71.6536, 
    -71.69765, -71.6836, -71.78859, -71.73223, -71.89316, -71.9515, 
    -72.11911, -72.22104, -72.32815, -72.37451, -72.38882, -72.39468 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  -1.621223, -1.620124, -1.620332, -1.619455, -1.619934, -1.619365, -1.62099, 
    -1.620089, -1.620659, -1.621111, -1.617776, -1.619413, -1.615986, 
    -1.617043, -1.614353, -1.616164, -1.613981, -1.614383, -1.613114, 
    -1.613477, -1.611894, -1.612946, -1.61103, -1.612133, -1.61197, 
    -1.612984, -1.619062, -1.617986, -1.619131, -1.618977, -1.619041, 
    -1.619932, -1.620394, -1.621291, -1.621125, -1.620457, -1.618907, 
    -1.619419, -1.61808, -1.61811, -1.616645, -1.617306, -1.614821, 
    -1.615521, -1.613461, -1.613986, -1.61349, -1.613637, -1.613488, 
    -1.614256, -1.613928, -1.614595, -1.617187, -1.616433, -1.618694, 
    -1.62009, -1.620955, -1.621584, -1.621496, -1.621331, -1.620454, 
    -1.619606, -1.618965, -1.618539, -1.618115, -1.616901, -1.616207, 
    -1.614689, -1.614945, -1.614496, -1.614037, -1.613292, -1.613412, 
    -1.613087, -1.614493, -1.613567, -1.615091, -1.614681, -1.618078, 
    -1.619277, -1.619852, -1.620295, -1.621429, -1.620651, -1.62096, 
    -1.620208, -1.61974, -1.619968, -1.618527, -1.619092, -1.616166, 
    -1.617424, -1.614091, -1.614891, -1.613895, -1.6144, -1.613541, 
    -1.614314, -1.61296, -1.612673, -1.612871, -1.612082, -1.614359, 
    -1.613497, -1.619978, -1.619942, -1.619761, -1.620555, -1.620599, 
    -1.6213, -1.620669, -1.620406, -1.619707, -1.619307, -1.61892, -1.618068, 
    -1.617136, -1.615807, -1.61484, -1.614189, -1.614584, -1.614236, 
    -1.614627, -1.614807, -1.612785, -1.61393, -1.612196, -1.61229, 
    -1.613082, -1.612279, -1.619915, -1.620128, -1.620894, -1.620295, 
    -1.621375, -1.620781, -1.620444, -1.619097, -1.618781, -1.618512, 
    -1.617963, -1.617273, -1.616064, -1.615, -1.614007, -1.614079, -1.614054, 
    -1.61384, -1.614381, -1.61375, -1.613652, -1.613921, -1.612303, 
    -1.612765, -1.612292, -1.612591, -1.620057, -1.619693, -1.619891, 
    -1.619523, -1.619789, -1.618628, -1.61828, -1.616636, -1.617291, 
    -1.616226, -1.617177, -1.617013, -1.616224, -1.61712, -1.615074, 
    -1.61649, -1.613831, -1.615287, -1.613741, -1.614012, -1.613556, 
    -1.613156, -1.612637, -1.611698, -1.611912, -1.611112, -1.619143, 
    -1.618676, -1.618703, -1.618203, -1.617838, -1.617033, -1.615753, 
    -1.61623, -1.615337, -1.615163, -1.61651, -1.615698, -1.618352, 
    -1.617937, -1.618173, -1.619115, -1.61614, -1.617673, -1.614827, 
    -1.615654, -1.613215, -1.61445, -1.612034, -1.61103, -1.610011, 
    -1.608896, -1.618405, -1.618724, -1.618139, -1.617363, -1.6166, 
    -1.615607, -1.615497, -1.615314, -1.614828, -1.614421, -1.615271, 
    -1.614317, -1.617871, -1.616, -1.618858, -1.618014, -1.617402, -1.617655, 
    -1.616281, -1.615961, -1.614667, -1.615327, -1.611292, -1.613092, 
    -1.607992, -1.60944, -1.618839, -1.618399, -1.616897, -1.617608, 
    -1.615532, -1.61503, -1.614604, -1.614082, -1.614015, -1.613702, 
    -1.614215, -1.613717, -1.615605, -1.614764, -1.617051, -1.616504, 
    -1.616751, -1.617032, -1.616164, -1.615261, -1.615218, -1.614937, 
    -1.614168, -1.615523, -1.611102, -1.613889, -1.617921, -1.617112, 
    -1.616968, -1.617287, -1.615077, -1.615883, -1.613707, -1.614294, 
    -1.613325, -1.613809, -1.613881, -1.614496, -1.614883, -1.61585, 
    -1.616632, -1.617238, -1.617095, -1.616428, -1.6152, -1.614019, 
    -1.614283, -1.613398, -1.615684, -1.614744, -1.615113, -1.614138, 
    -1.616248, -1.614525, -1.616696, -1.616501, -1.615898, -1.614696, 
    -1.614393, -1.614111, -1.61428, -1.615164, -1.615299, -1.615907, 
    -1.616087, -1.616542, -1.616929, -1.616581, -1.61622, -1.615154, 
    -1.614207, -1.613154, -1.612886, -1.611706, -1.6127, -1.611091, 
    -1.612509, -1.610023, -1.61439, -1.612503, -1.615863, -1.615498, 
    -1.614866, -1.613344, -1.614142, -1.613197, -1.615303, -1.616417, 
    -1.616675, -1.617205, -1.616663, -1.616706, -1.616188, -1.616353, 
    -1.615118, -1.615782, -1.613889, -1.613199, -1.611204, -1.609986, 
    -1.608701, -1.608143, -1.607971, -1.6079 ;

 FCH4 =
  1.822083e-13, 1.821208e-13, 1.821389e-13, 1.820604e-13, 1.821052e-13, 
    1.82052e-13, 1.821917e-13, 1.821169e-13, 1.821658e-13, 1.822011e-13, 
    1.818792e-13, 1.820567e-13, 1.806653e-13, 1.806556e-13, 1.806189e-13, 
    1.806657e-13, 1.80598e-13, 1.806218e-13, 1.805344e-13, 1.805645e-13, 
    1.803976e-13, 1.805192e-13, 1.802775e-13, 1.804303e-13, 1.80409e-13, 
    1.805225e-13, 1.820242e-13, 1.819033e-13, 1.820308e-13, 1.820148e-13, 
    1.820221e-13, 1.821042e-13, 1.821419e-13, 1.822146e-13, 1.822021e-13, 
    1.821485e-13, 1.820075e-13, 1.820588e-13, 1.819229e-13, 1.819263e-13, 
    1.806629e-13, 1.806484e-13, 1.806411e-13, 1.806607e-13, 1.805633e-13, 
    1.805997e-13, 1.805652e-13, 1.805764e-13, 1.80565e-13, 1.806151e-13, 
    1.805958e-13, 1.80632e-13, 1.80652e-13, 1.80665e-13, 1.819867e-13, 
    1.821148e-13, 1.821886e-13, 1.822355e-13, 1.822291e-13, 1.822166e-13, 
    1.821482e-13, 1.820761e-13, 1.820155e-13, 1.81972e-13, 1.819267e-13, 
    1.806591e-13, 1.806659e-13, 1.806352e-13, 1.806458e-13, 1.806267e-13, 
    1.806029e-13, 1.805491e-13, 1.805591e-13, 1.805311e-13, 1.806275e-13, 
    1.805702e-13, 1.806507e-13, 1.806357e-13, 1.819132e-13, 1.820453e-13, 
    1.820945e-13, 1.821354e-13, 1.822241e-13, 1.821643e-13, 1.821886e-13, 
    1.821292e-13, 1.820881e-13, 1.821088e-13, 1.819707e-13, 1.820275e-13, 
    1.806659e-13, 1.80645e-13, 1.80606e-13, 1.806438e-13, 1.805941e-13, 
    1.806231e-13, 1.805685e-13, 1.806187e-13, 1.805199e-13, 1.804907e-13, 
    1.805109e-13, 1.804261e-13, 1.806209e-13, 1.805651e-13, 1.821093e-13, 
    1.82106e-13, 1.820903e-13, 1.821564e-13, 1.821603e-13, 1.822149e-13, 
    1.821666e-13, 1.821447e-13, 1.820857e-13, 1.82048e-13, 1.820103e-13, 
    1.819206e-13, 1.806535e-13, 1.806642e-13, 1.806419e-13, 1.80612e-13, 
    1.806318e-13, 1.806145e-13, 1.806336e-13, 1.80641e-13, 1.805019e-13, 
    1.805955e-13, 1.804395e-13, 1.804506e-13, 1.805304e-13, 1.804494e-13, 
    1.821037e-13, 1.821226e-13, 1.821841e-13, 1.821366e-13, 1.822205e-13, 
    1.82175e-13, 1.821469e-13, 1.820261e-13, 1.819968e-13, 1.819683e-13, 
    1.819093e-13, 1.806494e-13, 1.806659e-13, 1.806471e-13, 1.806013e-13, 
    1.806057e-13, 1.806042e-13, 1.805903e-13, 1.80622e-13, 1.805842e-13, 
    1.805766e-13, 1.805956e-13, 1.804521e-13, 1.805015e-13, 1.804509e-13, 
    1.80484e-13, 1.821166e-13, 1.82084e-13, 1.821018e-13, 1.820679e-13, 
    1.820919e-13, 1.819785e-13, 1.81941e-13, 1.806631e-13, 1.80649e-13, 
    1.806659e-13, 1.806522e-13, 1.806563e-13, 1.806656e-13, 1.806536e-13, 
    1.806488e-13, 1.806645e-13, 1.805897e-13, 1.806543e-13, 1.805836e-13, 
    1.806016e-13, 1.805706e-13, 1.805374e-13, 1.804883e-13, 1.80375e-13, 
    1.80404e-13, 1.802921e-13, 1.820326e-13, 1.819845e-13, 1.81989e-13, 
    1.819359e-13, 1.818944e-13, 1.806557e-13, 1.806638e-13, 1.806661e-13, 
    1.806571e-13, 1.806525e-13, 1.806644e-13, 1.80663e-13, 1.819508e-13, 
    1.819031e-13, 1.81932e-13, 1.820288e-13, 1.806659e-13, 1.818728e-13, 
    1.806413e-13, 1.806627e-13, 1.805425e-13, 1.806242e-13, 1.804191e-13, 
    1.802739e-13, 1.801044e-13, 1.798625e-13, 1.819572e-13, 1.819913e-13, 
    1.819294e-13, 1.806471e-13, 1.806634e-13, 1.806619e-13, 1.806603e-13, 
    1.806564e-13, 1.806417e-13, 1.806241e-13, 1.806548e-13, 1.806189e-13, 
    1.818914e-13, 1.806656e-13, 1.820036e-13, 1.819115e-13, 1.806457e-13, 
    1.81873e-13, 1.806659e-13, 1.806657e-13, 1.806345e-13, 1.806568e-13, 
    1.80313e-13, 1.805295e-13, 1.796464e-13, 1.799845e-13, 1.820028e-13, 
    1.819574e-13, 1.806588e-13, 1.818677e-13, 1.806609e-13, 1.806484e-13, 
    1.806327e-13, 1.80605e-13, 1.806016e-13, 1.805806e-13, 1.806134e-13, 
    1.805821e-13, 1.806619e-13, 1.806391e-13, 1.806553e-13, 1.806645e-13, 
    1.806613e-13, 1.806557e-13, 1.806662e-13, 1.806544e-13, 1.806541e-13, 
    1.80645e-13, 1.806047e-13, 1.806607e-13, 1.802767e-13, 1.805879e-13, 
    1.819049e-13, 1.806542e-13, 1.806573e-13, 1.806489e-13, 1.8065e-13, 
    1.806651e-13, 1.805811e-13, 1.806176e-13, 1.805523e-13, 1.805883e-13, 
    1.80593e-13, 1.806277e-13, 1.806435e-13, 1.806647e-13, 1.806631e-13, 
    1.806503e-13, 1.806542e-13, 1.806651e-13, 1.80653e-13, 1.806012e-13, 
    1.80616e-13, 1.805583e-13, 1.806631e-13, 1.806378e-13, 1.806506e-13, 
    1.806088e-13, 1.80666e-13, 1.806247e-13, 1.806621e-13, 1.806645e-13, 
    1.806652e-13, 1.80635e-13, 1.806227e-13, 1.806067e-13, 1.806169e-13, 
    1.806521e-13, 1.806559e-13, 1.806654e-13, 1.80666e-13, 1.806641e-13, 
    1.80658e-13, 1.806637e-13, 1.80666e-13, 1.806522e-13, 1.806121e-13, 
    1.805369e-13, 1.805133e-13, 1.803704e-13, 1.804902e-13, 1.802741e-13, 
    1.804631e-13, 1.800931e-13, 1.806198e-13, 1.804681e-13, 1.806651e-13, 
    1.806603e-13, 1.806419e-13, 1.80551e-13, 1.80609e-13, 1.805391e-13, 
    1.806561e-13, 1.806651e-13, 1.806624e-13, 1.806513e-13, 1.806626e-13, 
    1.80662e-13, 1.806662e-13, 1.806656e-13, 1.806512e-13, 1.806643e-13, 
    1.805931e-13, 1.805399e-13, 1.803047e-13, 1.800943e-13, 1.798253e-13, 
    1.796881e-13, 1.79644e-13, 1.796253e-13 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  8.152351, 8.16757, 8.16461, 8.17688, 8.170083, 8.178106, 8.155436, 
    8.168174, 8.160041, 8.153724, 8.200683, 8.177426, 8.224936, 8.210042, 
    8.249128, 8.222612, 8.25417, 8.248413, 8.265776, 8.260797, 8.283039, 
    8.268074, 8.294612, 8.279467, 8.281831, 8.26758, 8.182105, 8.197783, 
    8.181176, 8.18341, 8.182409, 8.170222, 8.164062, 8.151194, 8.153528, 
    8.162982, 8.184415, 8.177148, 8.195486, 8.195071, 8.215529, 8.206296, 
    8.242379, 8.230966, 8.261005, 8.253834, 8.260667, 8.258595, 8.260694, 
    8.25018, 8.254683, 8.245443, 8.208023, 8.21853, 8.187241, 8.168467, 
    8.155993, 8.147153, 8.148402, 8.150784, 8.163037, 8.174573, 8.183345, 
    8.189219, 8.195011, 8.212554, 8.221869, 8.244366, 8.240589, 8.246991, 
    8.253121, 8.263421, 8.261725, 8.266266, 8.246826, 8.259737, 8.23685, 
    8.244256, 8.196571, 8.179108, 8.171686, 8.165178, 8.149363, 8.160279, 
    8.155972, 8.166226, 8.172743, 8.169522, 8.189379, 8.181655, 8.222423, 
    8.204834, 8.252406, 8.241364, 8.255057, 8.248067, 8.260047, 8.249264, 
    8.267958, 8.272033, 8.269247, 8.279963, 8.248666, 8.260664, 8.169431, 
    8.169957, 8.172407, 8.161636, 8.160979, 8.151129, 8.159894, 8.163629, 
    8.17312, 8.178717, 8.184041, 8.195765, 8.208869, 8.227248, 8.24208, 
    8.250978, 8.245522, 8.250339, 8.244953, 8.242432, 8.270505, 8.254723, 
    8.27842, 8.277107, 8.266373, 8.277256, 8.170327, 8.1673, 8.156799, 
    8.165016, 8.150057, 8.158423, 8.163238, 8.181813, 8.185896, 8.18968, 
    8.197162, 8.206768, 8.223657, 8.239982, 8.253479, 8.25249, 8.252838, 
    8.255856, 8.248381, 8.257084, 8.258543, 8.254724, 8.276932, 8.270579, 
    8.27708, 8.272943, 8.168284, 8.173371, 8.170625, 8.175784, 8.172152, 
    8.188315, 8.19317, 8.215921, 8.206577, 8.221459, 8.208089, 8.210455, 
    8.221937, 8.208812, 8.239162, 8.218054, 8.255973, 8.234811, 8.257201, 
    8.253421, 8.259683, 8.265294, 8.272364, 8.285421, 8.282396, 8.293336, 
    8.180939, 8.187529, 8.186951, 8.193855, 8.198963, 8.210048, 8.227867, 
    8.221162, 8.23348, 8.235955, 8.217244, 8.228723, 8.191944, 8.197871, 
    8.194345, 8.181457, 8.222702, 8.201504, 8.242298, 8.229181, 8.264493, 
    8.247689, 8.28073, 8.294894, 8.308276, 8.323919, 8.191131, 8.186649, 
    8.194677, 8.205787, 8.216122, 8.229883, 8.231295, 8.233875, 8.242163, 
    8.2478, 8.234688, 8.249215, 8.199239, 8.224546, 8.184954, 8.196852, 
    8.205132, 8.201502, 8.220397, 8.224857, 8.244608, 8.233623, 8.291391, 
    8.266473, 8.335874, 8.316402, 8.185083, 8.191116, 8.212138, 8.202129, 
    8.230804, 8.23947, 8.245239, 8.252614, 8.253414, 8.25779, 8.250621, 
    8.257508, 8.229912, 8.243106, 8.209735, 8.217453, 8.213902, 8.210008, 
    8.222035, 8.234868, 8.235148, 8.240859, 8.252481, 8.230921, 8.2946, 
    8.256166, 8.197699, 8.20933, 8.210999, 8.206488, 8.237171, 8.226036, 
    8.257684, 8.249542, 8.262889, 8.256252, 8.255277, 8.246767, 8.241475, 
    8.226545, 8.215715, 8.207143, 8.209135, 8.218555, 8.235655, 8.253484, 
    8.249921, 8.261874, 8.228721, 8.243517, 8.236814, 8.251745, 8.220982, 
    8.247384, 8.214655, 8.21738, 8.225815, 8.24441, 8.24819, 8.252218, 
    8.249734, 8.236091, 8.234123, 8.225612, 8.223261, 8.216786, 8.211429, 
    8.216323, 8.221464, 8.236099, 8.250914, 8.265373, 8.268918, 8.285843, 
    8.272052, 8.294812, 8.27544, 8.30902, 8.248835, 8.274889, 8.226201, 
    8.231256, 8.241993, 8.263058, 8.251682, 8.264991, 8.234047, 8.218878, 
    8.214966, 8.207663, 8.215134, 8.214525, 8.221682, 8.219381, 8.236586, 
    8.227339, 8.25525, 8.264887, 8.292186, 8.308972, 8.326117, 8.333694, 
    8.336004, 8.336968 ;

 FGR =
  -324.559, -325.3203, -325.1727, -325.7857, -325.4464, -325.8472, -324.7141, 
    -325.3498, -324.9445, -324.6286, -326.9725, -325.8132, -328.1822, 
    -327.4428, -329.3127, -328.0661, -329.5625, -329.2789, -330.1368, 
    -329.8911, -330.9849, -330.2503, -331.5549, -330.8104, -330.9262, 
    -330.2257, -326.0483, -326.8278, -326.0017, -326.113, -326.0635, 
    -325.4528, -325.1437, -324.502, -324.6188, -325.0908, -326.1631, 
    -325.8003, -326.7181, -326.6974, -327.7161, -327.2568, -328.9802, 
    -328.4834, -329.9015, -329.5471, -329.8845, -329.7824, -329.8858, 
    -329.3662, -329.5887, -329.1321, -327.3425, -327.8649, -326.3049, 
    -325.363, -324.7417, -324.2995, -324.362, -324.4808, -325.0936, 
    -325.6713, -326.1108, -326.4046, -326.6944, -327.5652, -328.0299, 
    -329.0778, -328.892, -329.2079, -329.5119, -330.0203, -329.9368, 
    -330.1605, -329.2007, -329.838, -328.7755, -329.0733, -326.767, 
    -325.8985, -325.5241, -325.2008, -324.4099, -324.9557, -324.7404, 
    -325.254, -325.5795, -325.4188, -326.4127, -326.026, -328.0575, 
    -327.1831, -329.4764, -328.9302, -329.6076, -329.2622, -329.8535, 
    -329.3214, -330.2442, -330.4445, -330.3075, -330.8358, -329.2917, 
    -329.8839, -325.414, -325.4402, -325.5629, -325.0235, -324.9909, 
    -324.4985, -324.9372, -325.1235, -325.5989, -325.8788, -326.1453, 
    -326.7314, -327.3839, -328.2978, -328.9655, -329.4062, -329.1364, 
    -329.3745, -329.1081, -328.9835, -330.369, -329.5904, -330.7597, 
    -330.6953, -330.1655, -330.7025, -325.4587, -325.3078, -324.7822, 
    -325.1936, -324.445, -324.8632, -325.1032, -326.0328, -326.2385, 
    -326.4272, -326.8015, -327.2802, -328.1196, -328.8611, -329.5298, 
    -329.481, -329.4981, -329.6469, -329.2775, -329.7076, -329.7792, 
    -329.5911, -330.6866, -330.3737, -330.6939, -330.4903, -325.357, 
    -325.6111, -325.4737, -325.7316, -325.5495, -326.3578, -326.6002, 
    -327.7343, -327.2705, -328.0103, -327.3461, -327.4634, -328.0318, 
    -327.3824, -328.8196, -327.8397, -329.6527, -328.6712, -329.7134, 
    -329.5269, -329.8362, -330.1126, -330.4615, -331.1035, -330.955, 
    -331.493, -325.9902, -326.3191, -326.2913, -326.6363, -326.891, 
    -327.4438, -328.3291, -327.9966, -328.6083, -328.7307, -327.802, 
    -328.3711, -326.5401, -326.8351, -326.6604, -326.0155, -328.0717, 
    -327.0165, -328.9762, -328.3946, -330.0731, -329.2421, -330.8731, 
    -331.5675, -332.2264, -332.9903, -326.4999, -326.2763, -326.6777, 
    -327.23, -327.7456, -328.4292, -328.4998, -328.6275, -328.9701, -329.249, 
    -328.6668, -329.319, -326.9011, -328.1638, -326.1907, -326.784, -327.198, 
    -327.0176, -327.9589, -328.1803, -329.09, -328.6154, -331.3951, 
    -330.1694, -333.5759, -332.623, -326.1979, -326.4997, -327.5468, 
    -327.049, -328.4755, -328.8363, -329.1224, -329.4863, -329.5264, 
    -329.7422, -329.3885, -329.7287, -328.4307, -329.0165, -327.4285, 
    -327.8119, -327.6359, -327.442, -328.0402, -328.6755, -328.6909, 
    -328.9046, -329.4747, -328.4813, -331.5499, -329.6576, -326.8285, 
    -327.4062, -327.4909, -327.2667, -328.7909, -328.2384, -329.7372, 
    -329.3352, -329.9944, -329.6667, -329.6183, -329.1979, -328.9356, 
    -328.2634, -327.7253, -327.2995, -327.3986, -327.8664, -328.7148, 
    -329.5293, -329.3528, -329.9443, -328.3719, -329.0361, -328.7725, 
    -329.4438, -327.9874, -329.2235, -327.6733, -327.8087, -328.2274, 
    -329.0793, -329.2682, -329.4667, -329.3446, -328.7367, -328.6396, 
    -328.2177, -328.1003, -327.7794, -327.5128, -327.7559, -328.0109, 
    -328.7377, -329.4022, -330.1163, -330.2918, -331.1217, -330.4436, 
    -331.5601, -330.607, -332.2589, -329.2973, -330.5827, -328.2471, 
    -328.498, -328.96, -330.0006, -329.4408, -330.0964, -328.636, -327.8816, 
    -327.6887, -327.325, -327.697, -327.6668, -328.0227, -327.9085, 
    -328.7618, -328.3035, -329.6166, -330.0917, -331.4359, -332.2589, 
    -333.0998, -333.47, -333.5829, -333.63 ;

 FGR12 =
  -224.3942, -224.3558, -224.3631, -224.3327, -224.3492, -224.3296, 
    -224.3861, -224.3545, -224.3744, -224.3903, -224.2753, -224.3313, 
    -224.2157, -224.2509, -224.1633, -224.2217, -224.1515, -224.1644, 
    -224.1241, -224.1356, -224.0863, -224.1189, -224.0599, -224.0937, 
    -224.0886, -224.1201, -224.3193, -224.2825, -224.3217, -224.3164, 
    -224.3186, -224.3492, -224.3651, -224.3967, -224.3908, -224.3674, 
    -224.314, -224.3315, -224.2859, -224.2869, -224.2376, -224.2598, 
    -224.1784, -224.2006, -224.135, -224.1517, -224.136, -224.1406, 
    -224.1359, -224.1603, -224.1498, -224.1712, -224.2557, -224.2305, 
    -224.3067, -224.3545, -224.3848, -224.4071, -224.4039, -224.398, 
    -224.3672, -224.3379, -224.316, -224.3014, -224.2871, -224.246, 
    -224.2231, -224.1741, -224.1825, -224.168, -224.1533, -224.1297, 
    -224.1335, -224.1233, -224.1679, -224.1384, -224.1866, -224.1739, 
    -224.2856, -224.3267, -224.3463, -224.3617, -224.4016, -224.3741, 
    -224.385, -224.3587, -224.3426, -224.3504, -224.301, -224.3203, 
    -224.2217, -224.2637, -224.155, -224.1807, -224.1488, -224.1649, 
    -224.1376, -224.1622, -224.1193, -224.1104, -224.1165, -224.0921, 
    -224.1636, -224.1362, -224.3508, -224.3495, -224.3433, -224.3708, 
    -224.3723, -224.397, -224.3748, -224.3656, -224.3414, -224.3277, 
    -224.3145, -224.2854, -224.254, -224.2099, -224.1791, -224.1582, 
    -224.1708, -224.1597, -224.1722, -224.178, -224.1138, -224.1499, 
    -224.0956, -224.0985, -224.1232, -224.0981, -224.3486, -224.356, 
    -224.3827, -224.3618, -224.3997, -224.3787, -224.3669, -224.3204, 
    -224.3098, -224.3004, -224.2819, -224.2586, -224.2184, -224.1842, 
    -224.1524, -224.1546, -224.1539, -224.147, -224.1643, -224.1442, 
    -224.1411, -224.1496, -224.0989, -224.1133, -224.0985, -224.1078, 
    -224.3535, -224.3409, -224.3478, -224.3351, -224.3442, -224.3044, 
    -224.2925, -224.2372, -224.2592, -224.2237, -224.2554, -224.2499, 
    -224.2236, -224.2535, -224.1866, -224.2325, -224.1467, -224.1929, 
    -224.1439, -224.1525, -224.1381, -224.1255, -224.1093, -224.0803, 
    -224.0869, -224.0624, -224.3221, -224.3061, -224.307, -224.29, -224.2777, 
    -224.2506, -224.2081, -224.2239, -224.1946, -224.1889, -224.2332, 
    -224.2063, -224.295, -224.281, -224.289, -224.3211, -224.2209, -224.2721, 
    -224.1786, -224.205, -224.1273, -224.1665, -224.0906, -224.06, -224.0294, 
    -223.9965, -224.2968, -224.3078, -224.2879, -224.2616, -224.2362, 
    -224.2033, -224.1998, -224.1938, -224.1787, -224.1656, -224.1924, 
    -224.1622, -224.2787, -224.2162, -224.3124, -224.2835, -224.2629, 
    -224.2715, -224.2256, -224.215, -224.1735, -224.1942, -224.0679, 
    -224.1235, -223.9703, -224.0125, -224.3118, -224.2966, -224.246, 
    -224.2699, -224.2009, -224.1852, -224.1715, -224.1547, -224.1526, 
    -224.1427, -224.159, -224.1431, -224.2033, -224.1766, -224.2512, 
    -224.2329, -224.2412, -224.2506, -224.2217, -224.192, -224.1907, 
    -224.1822, -224.1574, -224.2007, -224.0621, -224.1486, -224.2805, 
    -224.2532, -224.2484, -224.2591, -224.1861, -224.2124, -224.1428, 
    -224.1615, -224.1307, -224.1461, -224.1483, -224.168, -224.1804, 
    -224.2114, -224.2372, -224.2575, -224.2527, -224.2304, -224.1901, 
    -224.1527, -224.1611, -224.1331, -224.206, -224.176, -224.1873, 
    -224.1565, -224.2245, -224.1688, -224.2394, -224.2329, -224.213, 
    -224.1743, -224.1647, -224.1556, -224.161, -224.189, -224.1933, 
    -224.2133, -224.2191, -224.2342, -224.2471, -224.2355, -224.2236, 
    -224.1886, -224.1587, -224.1254, -224.1171, -224.0805, -224.1112, 
    -224.0618, -224.1053, -224.0297, -224.1646, -224.105, -224.2118, 
    -224.1998, -224.1799, -224.1313, -224.1567, -224.1267, -224.1934, 
    -224.2301, -224.2387, -224.2564, -224.2383, -224.2397, -224.2225, 
    -224.228, -224.1875, -224.2091, -224.1486, -224.1268, -224.0652, 
    -224.0287, -223.9908, -223.9747, -223.9697, -223.9677 ;

 FGR_R =
  -324.559, -325.3203, -325.1727, -325.7857, -325.4464, -325.8472, -324.7141, 
    -325.3498, -324.9445, -324.6286, -326.9725, -325.8132, -328.1822, 
    -327.4428, -329.3127, -328.0661, -329.5625, -329.2789, -330.1368, 
    -329.8911, -330.9849, -330.2503, -331.5549, -330.8104, -330.9262, 
    -330.2257, -326.0483, -326.8278, -326.0017, -326.113, -326.0635, 
    -325.4528, -325.1437, -324.502, -324.6188, -325.0908, -326.1631, 
    -325.8003, -326.7181, -326.6974, -327.7161, -327.2568, -328.9802, 
    -328.4834, -329.9015, -329.5471, -329.8845, -329.7824, -329.8858, 
    -329.3662, -329.5887, -329.1321, -327.3425, -327.8649, -326.3049, 
    -325.363, -324.7417, -324.2995, -324.362, -324.4808, -325.0936, 
    -325.6713, -326.1108, -326.4046, -326.6944, -327.5652, -328.0299, 
    -329.0778, -328.892, -329.2079, -329.5119, -330.0203, -329.9368, 
    -330.1605, -329.2007, -329.838, -328.7755, -329.0733, -326.767, 
    -325.8985, -325.5241, -325.2008, -324.4099, -324.9557, -324.7404, 
    -325.254, -325.5795, -325.4188, -326.4127, -326.026, -328.0575, 
    -327.1831, -329.4764, -328.9302, -329.6076, -329.2622, -329.8535, 
    -329.3214, -330.2442, -330.4445, -330.3075, -330.8358, -329.2917, 
    -329.8839, -325.414, -325.4402, -325.5629, -325.0235, -324.9909, 
    -324.4985, -324.9372, -325.1235, -325.5989, -325.8788, -326.1453, 
    -326.7314, -327.3839, -328.2978, -328.9655, -329.4062, -329.1364, 
    -329.3745, -329.1081, -328.9835, -330.369, -329.5904, -330.7597, 
    -330.6953, -330.1655, -330.7025, -325.4587, -325.3078, -324.7822, 
    -325.1936, -324.445, -324.8632, -325.1032, -326.0328, -326.2385, 
    -326.4272, -326.8015, -327.2802, -328.1196, -328.8611, -329.5298, 
    -329.481, -329.4981, -329.6469, -329.2775, -329.7076, -329.7792, 
    -329.5911, -330.6866, -330.3737, -330.6939, -330.4903, -325.357, 
    -325.6111, -325.4737, -325.7316, -325.5495, -326.3578, -326.6002, 
    -327.7343, -327.2705, -328.0103, -327.3461, -327.4634, -328.0318, 
    -327.3824, -328.8196, -327.8397, -329.6527, -328.6712, -329.7134, 
    -329.5269, -329.8362, -330.1126, -330.4615, -331.1035, -330.955, 
    -331.493, -325.9902, -326.3191, -326.2913, -326.6363, -326.891, 
    -327.4438, -328.3291, -327.9966, -328.6083, -328.7307, -327.802, 
    -328.3711, -326.5401, -326.8351, -326.6604, -326.0155, -328.0717, 
    -327.0165, -328.9762, -328.3946, -330.0731, -329.2421, -330.8731, 
    -331.5675, -332.2264, -332.9903, -326.4999, -326.2763, -326.6777, 
    -327.23, -327.7456, -328.4292, -328.4998, -328.6275, -328.9701, -329.249, 
    -328.6668, -329.319, -326.9011, -328.1638, -326.1907, -326.784, -327.198, 
    -327.0176, -327.9589, -328.1803, -329.09, -328.6154, -331.3951, 
    -330.1694, -333.5759, -332.623, -326.1979, -326.4997, -327.5468, 
    -327.049, -328.4755, -328.8363, -329.1224, -329.4863, -329.5264, 
    -329.7422, -329.3885, -329.7287, -328.4307, -329.0165, -327.4285, 
    -327.8119, -327.6359, -327.442, -328.0402, -328.6755, -328.6909, 
    -328.9046, -329.4747, -328.4813, -331.5499, -329.6576, -326.8285, 
    -327.4062, -327.4909, -327.2667, -328.7909, -328.2384, -329.7372, 
    -329.3352, -329.9944, -329.6667, -329.6183, -329.1979, -328.9356, 
    -328.2634, -327.7253, -327.2995, -327.3986, -327.8664, -328.7148, 
    -329.5293, -329.3528, -329.9443, -328.3719, -329.0361, -328.7725, 
    -329.4438, -327.9874, -329.2235, -327.6733, -327.8087, -328.2274, 
    -329.0793, -329.2682, -329.4667, -329.3446, -328.7367, -328.6396, 
    -328.2177, -328.1003, -327.7794, -327.5128, -327.7559, -328.0109, 
    -328.7377, -329.4022, -330.1163, -330.2918, -331.1217, -330.4436, 
    -331.5601, -330.607, -332.2589, -329.2973, -330.5827, -328.2471, 
    -328.498, -328.96, -330.0006, -329.4408, -330.0964, -328.636, -327.8816, 
    -327.6887, -327.325, -327.697, -327.6668, -328.0227, -327.9085, 
    -328.7618, -328.3035, -329.6166, -330.0917, -331.4359, -332.2589, 
    -333.0998, -333.47, -333.5829, -333.63 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  74.77462, 74.82764, 74.81736, 74.86006, 74.83642, 74.86435, 74.78542, 
    74.82969, 74.80147, 74.77947, 74.94284, 74.86198, 75.02758, 74.97579, 
    75.10563, 75.01944, 75.12312, 75.10326, 75.16334, 75.14614, 75.22269, 
    75.17128, 75.26258, 75.21048, 75.21858, 75.16956, 74.87837, 74.93272, 
    74.87512, 74.88288, 74.87943, 74.83686, 74.81534, 74.77065, 74.77879, 
    74.81166, 74.88637, 74.86108, 74.92506, 74.92361, 74.99493, 74.96276, 
    75.08235, 75.0487, 75.14686, 75.12205, 75.14567, 75.13853, 75.14576, 
    75.10938, 75.12496, 75.09299, 74.96877, 75.00535, 74.89626, 74.8306, 
    74.78735, 74.75655, 74.7609, 74.76917, 74.81185, 74.85209, 74.88273, 
    74.90321, 74.9234, 74.98435, 75.01691, 75.08918, 75.07617, 75.09829, 
    75.11958, 75.15517, 75.14934, 75.16499, 75.09779, 75.14241, 75.06917, 
    75.08887, 74.92846, 74.86793, 74.84182, 74.81932, 74.76424, 74.80225, 
    74.78726, 74.82302, 74.84569, 74.8345, 74.90377, 74.87682, 75.01884, 
    74.9576, 75.1171, 75.07885, 75.12628, 75.1021, 75.1435, 75.10624, 
    75.17085, 75.18487, 75.17528, 75.21226, 75.10416, 75.14563, 74.83416, 
    74.83598, 74.84453, 74.80697, 74.8047, 74.77041, 74.80096, 74.81393, 
    74.84704, 74.86655, 74.88513, 74.92599, 74.97166, 75.03568, 75.08132, 
    75.11218, 75.09329, 75.10996, 75.09131, 75.08258, 75.17959, 75.12508, 
    75.20694, 75.20242, 75.16534, 75.20293, 74.83727, 74.82677, 74.79017, 
    74.81882, 74.76669, 74.79581, 74.81252, 74.87729, 74.89162, 74.90479, 
    74.93089, 74.96441, 75.0232, 75.07401, 75.12084, 75.11742, 75.11862, 
    75.12904, 75.10317, 75.13329, 75.13829, 75.12512, 75.20182, 75.17992, 
    75.20233, 75.18808, 74.83019, 74.84789, 74.83832, 74.85629, 74.84359, 
    74.89995, 74.91684, 74.9962, 74.96372, 75.01553, 74.96902, 74.97723, 
    75.01703, 74.97157, 75.0711, 75.00358, 75.12944, 75.06184, 75.13369, 
    75.12064, 75.1423, 75.16164, 75.18607, 75.231, 75.2206, 75.25826, 
    74.87432, 74.89725, 74.89531, 74.91936, 74.93715, 74.97587, 75.03788, 
    75.01458, 75.05745, 75.06602, 75.00095, 75.04082, 74.91265, 74.93324, 
    74.92104, 74.87608, 75.01984, 74.94593, 75.08207, 75.04247, 75.15887, 
    75.10069, 75.21487, 75.26346, 75.30957, 75.363, 74.90985, 74.89426, 
    74.92224, 74.96088, 74.997, 75.0449, 75.04984, 75.05879, 75.08164, 
    75.10117, 75.06154, 75.10608, 74.93785, 75.02629, 74.88829, 74.92966, 
    74.95864, 74.94601, 75.01194, 75.02745, 75.09003, 75.05795, 75.25139, 
    75.16561, 75.40396, 75.3373, 74.88879, 74.90984, 74.98307, 74.94821, 
    75.04814, 75.07227, 75.09231, 75.11779, 75.1206, 75.1357, 75.11095, 
    75.13477, 75.045, 75.08489, 74.97479, 75.00164, 74.98932, 74.97575, 
    75.01764, 75.06215, 75.06323, 75.07705, 75.11696, 75.04855, 75.26221, 
    75.12977, 74.93278, 74.97322, 74.97916, 74.96346, 75.07024, 75.03152, 
    75.13536, 75.10721, 75.15337, 75.13042, 75.12704, 75.0976, 75.07923, 
    75.03327, 74.99557, 74.96576, 74.9727, 75.00546, 75.0649, 75.1208, 
    75.10844, 75.14986, 75.04089, 75.08627, 75.06895, 75.11481, 75.01393, 
    75.09937, 74.99194, 75.00143, 75.03075, 75.08928, 75.10252, 75.11642, 
    75.10787, 75.06644, 75.05964, 75.03008, 75.02185, 74.99937, 74.9807, 
    74.99773, 75.01557, 75.06651, 75.1119, 75.1619, 75.17419, 75.23225, 
    75.1848, 75.26292, 75.19622, 75.31182, 75.10455, 75.19453, 75.03214, 
    75.04971, 75.08093, 75.15379, 75.1146, 75.1605, 75.05939, 75.00652, 
    74.99302, 74.96754, 74.9936, 74.99149, 75.01641, 75.00841, 75.06821, 
    75.03609, 75.12691, 75.16017, 75.25426, 75.31184, 75.37067, 75.39656, 
    75.40446, 75.40775 ;

 FIRA_R =
  74.77462, 74.82764, 74.81736, 74.86006, 74.83642, 74.86435, 74.78542, 
    74.82969, 74.80147, 74.77947, 74.94284, 74.86198, 75.02758, 74.97579, 
    75.10563, 75.01944, 75.12312, 75.10326, 75.16334, 75.14614, 75.22269, 
    75.17128, 75.26258, 75.21048, 75.21858, 75.16956, 74.87837, 74.93272, 
    74.87512, 74.88288, 74.87943, 74.83686, 74.81534, 74.77065, 74.77879, 
    74.81166, 74.88637, 74.86108, 74.92506, 74.92361, 74.99493, 74.96276, 
    75.08235, 75.0487, 75.14686, 75.12205, 75.14567, 75.13853, 75.14576, 
    75.10938, 75.12496, 75.09299, 74.96877, 75.00535, 74.89626, 74.8306, 
    74.78735, 74.75655, 74.7609, 74.76917, 74.81185, 74.85209, 74.88273, 
    74.90321, 74.9234, 74.98435, 75.01691, 75.08918, 75.07617, 75.09829, 
    75.11958, 75.15517, 75.14934, 75.16499, 75.09779, 75.14241, 75.06917, 
    75.08887, 74.92846, 74.86793, 74.84182, 74.81932, 74.76424, 74.80225, 
    74.78726, 74.82302, 74.84569, 74.8345, 74.90377, 74.87682, 75.01884, 
    74.9576, 75.1171, 75.07885, 75.12628, 75.1021, 75.1435, 75.10624, 
    75.17085, 75.18487, 75.17528, 75.21226, 75.10416, 75.14563, 74.83416, 
    74.83598, 74.84453, 74.80697, 74.8047, 74.77041, 74.80096, 74.81393, 
    74.84704, 74.86655, 74.88513, 74.92599, 74.97166, 75.03568, 75.08132, 
    75.11218, 75.09329, 75.10996, 75.09131, 75.08258, 75.17959, 75.12508, 
    75.20694, 75.20242, 75.16534, 75.20293, 74.83727, 74.82677, 74.79017, 
    74.81882, 74.76669, 74.79581, 74.81252, 74.87729, 74.89162, 74.90479, 
    74.93089, 74.96441, 75.0232, 75.07401, 75.12084, 75.11742, 75.11862, 
    75.12904, 75.10317, 75.13329, 75.13829, 75.12512, 75.20182, 75.17992, 
    75.20233, 75.18808, 74.83019, 74.84789, 74.83832, 74.85629, 74.84359, 
    74.89995, 74.91684, 74.9962, 74.96372, 75.01553, 74.96902, 74.97723, 
    75.01703, 74.97157, 75.0711, 75.00358, 75.12944, 75.06184, 75.13369, 
    75.12064, 75.1423, 75.16164, 75.18607, 75.231, 75.2206, 75.25826, 
    74.87432, 74.89725, 74.89531, 74.91936, 74.93715, 74.97587, 75.03788, 
    75.01458, 75.05745, 75.06602, 75.00095, 75.04082, 74.91265, 74.93324, 
    74.92104, 74.87608, 75.01984, 74.94593, 75.08207, 75.04247, 75.15887, 
    75.10069, 75.21487, 75.26346, 75.30957, 75.363, 74.90985, 74.89426, 
    74.92224, 74.96088, 74.997, 75.0449, 75.04984, 75.05879, 75.08164, 
    75.10117, 75.06154, 75.10608, 74.93785, 75.02629, 74.88829, 74.92966, 
    74.95864, 74.94601, 75.01194, 75.02745, 75.09003, 75.05795, 75.25139, 
    75.16561, 75.40396, 75.3373, 74.88879, 74.90984, 74.98307, 74.94821, 
    75.04814, 75.07227, 75.09231, 75.11779, 75.1206, 75.1357, 75.11095, 
    75.13477, 75.045, 75.08489, 74.97479, 75.00164, 74.98932, 74.97575, 
    75.01764, 75.06215, 75.06323, 75.07705, 75.11696, 75.04855, 75.26221, 
    75.12977, 74.93278, 74.97322, 74.97916, 74.96346, 75.07024, 75.03152, 
    75.13536, 75.10721, 75.15337, 75.13042, 75.12704, 75.0976, 75.07923, 
    75.03327, 74.99557, 74.96576, 74.9727, 75.00546, 75.0649, 75.1208, 
    75.10844, 75.14986, 75.04089, 75.08627, 75.06895, 75.11481, 75.01393, 
    75.09937, 74.99194, 75.00143, 75.03075, 75.08928, 75.10252, 75.11642, 
    75.10787, 75.06644, 75.05964, 75.03008, 75.02185, 74.99937, 74.9807, 
    74.99773, 75.01557, 75.06651, 75.1119, 75.1619, 75.17419, 75.23225, 
    75.1848, 75.26292, 75.19622, 75.31182, 75.10455, 75.19453, 75.03214, 
    75.04971, 75.08093, 75.15379, 75.1146, 75.1605, 75.05939, 75.00652, 
    74.99302, 74.96754, 74.9936, 74.99149, 75.01641, 75.00841, 75.06821, 
    75.03609, 75.12691, 75.16017, 75.25426, 75.31184, 75.37067, 75.39656, 
    75.40446, 75.40775 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  263.7356, 263.7886, 263.7783, 263.821, 263.7974, 263.8253, 263.7464, 
    263.7906, 263.7624, 263.7404, 263.9038, 263.8229, 263.9885, 263.9367, 
    264.0666, 263.9804, 264.084, 264.0642, 264.1243, 264.1071, 264.1836, 
    264.1322, 264.2235, 264.1714, 264.1795, 264.1305, 263.8393, 263.8936, 
    263.8361, 263.8438, 263.8404, 263.7978, 263.7763, 263.7316, 263.7397, 
    263.7726, 263.8473, 263.822, 263.886, 263.8846, 263.9559, 263.9237, 
    264.0433, 264.0096, 264.1078, 264.083, 264.1066, 264.0995, 264.1067, 
    264.0703, 264.0859, 264.0539, 263.9297, 263.9663, 263.8572, 263.7915, 
    263.7483, 263.7175, 263.7218, 263.7301, 263.7728, 263.813, 263.8437, 
    263.8641, 263.8843, 263.9453, 263.9778, 264.0501, 264.0371, 264.0592, 
    264.0805, 264.1161, 264.1103, 264.1259, 264.0587, 264.1034, 264.0301, 
    264.0498, 263.8894, 263.8289, 263.8028, 263.7802, 263.7252, 263.7632, 
    263.7482, 263.784, 263.8066, 263.7954, 263.8647, 263.8378, 263.9798, 
    263.9185, 264.078, 264.0398, 264.0872, 264.063, 264.1044, 264.0672, 
    264.1318, 264.1458, 264.1362, 264.1732, 264.0651, 264.1066, 263.7951, 
    263.7969, 263.8055, 263.7679, 263.7656, 263.7314, 263.7619, 263.7749, 
    263.808, 263.8275, 263.8461, 263.8869, 263.9326, 263.9966, 264.0423, 
    264.0731, 264.0542, 264.0709, 264.0522, 264.0435, 264.1405, 264.086, 
    264.1679, 264.1634, 264.1263, 264.1639, 263.7982, 263.7877, 263.7511, 
    263.7798, 263.7276, 263.7567, 263.7735, 263.8382, 263.8526, 263.8657, 
    263.8918, 263.9254, 263.9841, 264.0349, 264.0818, 264.0784, 264.0796, 
    264.09, 264.0641, 264.0942, 264.0992, 264.0861, 264.1628, 264.1408, 
    264.1633, 264.149, 263.7911, 263.8088, 263.7993, 263.8172, 263.8045, 
    263.8609, 263.8778, 263.9571, 263.9247, 263.9765, 263.93, 263.9382, 
    263.978, 263.9325, 264.032, 263.9645, 264.0904, 264.0228, 264.0946, 
    264.0816, 264.1032, 264.1226, 264.147, 264.1919, 264.1815, 264.2192, 
    263.8353, 263.8582, 263.8563, 263.8803, 263.8981, 263.9368, 263.9988, 
    263.9755, 264.0184, 264.0269, 263.9619, 264.0018, 263.8736, 263.8942, 
    263.882, 263.837, 263.9808, 263.9069, 264.043, 264.0034, 264.1198, 
    264.0616, 264.1758, 264.2244, 264.2705, 264.3239, 263.8708, 263.8552, 
    263.8832, 263.9218, 263.9579, 264.0058, 264.0108, 264.0197, 264.0426, 
    264.0621, 264.0225, 264.067, 263.8988, 263.9872, 263.8492, 263.8906, 
    263.9196, 263.907, 263.9729, 263.9884, 264.051, 264.0189, 264.2123, 
    264.1266, 264.3649, 264.2982, 263.8497, 263.8708, 263.944, 263.9091, 
    264.0091, 264.0332, 264.0533, 264.0787, 264.0815, 264.0966, 264.0719, 
    264.0957, 264.006, 264.0458, 263.9357, 263.9626, 263.9503, 263.9367, 
    263.9786, 264.0231, 264.0242, 264.038, 264.0779, 264.0095, 264.2231, 
    264.0907, 263.8937, 263.9341, 263.9401, 263.9244, 264.0312, 263.9925, 
    264.0963, 264.0681, 264.1143, 264.0914, 264.088, 264.0585, 264.0402, 
    263.9942, 263.9565, 263.9267, 263.9336, 263.9664, 264.0258, 264.0817, 
    264.0694, 264.1108, 264.0018, 264.0472, 264.0299, 264.0757, 263.9749, 
    264.0603, 263.9529, 263.9624, 263.9917, 264.0502, 264.0635, 264.0774, 
    264.0688, 264.0274, 264.0206, 263.991, 263.9828, 263.9603, 263.9417, 
    263.9586, 263.9765, 264.0274, 264.0728, 264.1228, 264.1351, 264.1932, 
    264.1457, 264.2239, 264.1572, 264.2728, 264.0655, 264.1555, 263.9931, 
    264.0107, 264.0419, 264.1147, 264.0755, 264.1214, 264.0203, 263.9675, 
    263.9539, 263.9285, 263.9545, 263.9524, 263.9774, 263.9694, 264.0291, 
    263.997, 264.0879, 264.1211, 264.2152, 264.2728, 264.3316, 264.3575, 
    264.3654, 264.3687 ;

 FIRE_R =
  263.7356, 263.7886, 263.7783, 263.821, 263.7974, 263.8253, 263.7464, 
    263.7906, 263.7624, 263.7404, 263.9038, 263.8229, 263.9885, 263.9367, 
    264.0666, 263.9804, 264.084, 264.0642, 264.1243, 264.1071, 264.1836, 
    264.1322, 264.2235, 264.1714, 264.1795, 264.1305, 263.8393, 263.8936, 
    263.8361, 263.8438, 263.8404, 263.7978, 263.7763, 263.7316, 263.7397, 
    263.7726, 263.8473, 263.822, 263.886, 263.8846, 263.9559, 263.9237, 
    264.0433, 264.0096, 264.1078, 264.083, 264.1066, 264.0995, 264.1067, 
    264.0703, 264.0859, 264.0539, 263.9297, 263.9663, 263.8572, 263.7915, 
    263.7483, 263.7175, 263.7218, 263.7301, 263.7728, 263.813, 263.8437, 
    263.8641, 263.8843, 263.9453, 263.9778, 264.0501, 264.0371, 264.0592, 
    264.0805, 264.1161, 264.1103, 264.1259, 264.0587, 264.1034, 264.0301, 
    264.0498, 263.8894, 263.8289, 263.8028, 263.7802, 263.7252, 263.7632, 
    263.7482, 263.784, 263.8066, 263.7954, 263.8647, 263.8378, 263.9798, 
    263.9185, 264.078, 264.0398, 264.0872, 264.063, 264.1044, 264.0672, 
    264.1318, 264.1458, 264.1362, 264.1732, 264.0651, 264.1066, 263.7951, 
    263.7969, 263.8055, 263.7679, 263.7656, 263.7314, 263.7619, 263.7749, 
    263.808, 263.8275, 263.8461, 263.8869, 263.9326, 263.9966, 264.0423, 
    264.0731, 264.0542, 264.0709, 264.0522, 264.0435, 264.1405, 264.086, 
    264.1679, 264.1634, 264.1263, 264.1639, 263.7982, 263.7877, 263.7511, 
    263.7798, 263.7276, 263.7567, 263.7735, 263.8382, 263.8526, 263.8657, 
    263.8918, 263.9254, 263.9841, 264.0349, 264.0818, 264.0784, 264.0796, 
    264.09, 264.0641, 264.0942, 264.0992, 264.0861, 264.1628, 264.1408, 
    264.1633, 264.149, 263.7911, 263.8088, 263.7993, 263.8172, 263.8045, 
    263.8609, 263.8778, 263.9571, 263.9247, 263.9765, 263.93, 263.9382, 
    263.978, 263.9325, 264.032, 263.9645, 264.0904, 264.0228, 264.0946, 
    264.0816, 264.1032, 264.1226, 264.147, 264.1919, 264.1815, 264.2192, 
    263.8353, 263.8582, 263.8563, 263.8803, 263.8981, 263.9368, 263.9988, 
    263.9755, 264.0184, 264.0269, 263.9619, 264.0018, 263.8736, 263.8942, 
    263.882, 263.837, 263.9808, 263.9069, 264.043, 264.0034, 264.1198, 
    264.0616, 264.1758, 264.2244, 264.2705, 264.3239, 263.8708, 263.8552, 
    263.8832, 263.9218, 263.9579, 264.0058, 264.0108, 264.0197, 264.0426, 
    264.0621, 264.0225, 264.067, 263.8988, 263.9872, 263.8492, 263.8906, 
    263.9196, 263.907, 263.9729, 263.9884, 264.051, 264.0189, 264.2123, 
    264.1266, 264.3649, 264.2982, 263.8497, 263.8708, 263.944, 263.9091, 
    264.0091, 264.0332, 264.0533, 264.0787, 264.0815, 264.0966, 264.0719, 
    264.0957, 264.006, 264.0458, 263.9357, 263.9626, 263.9503, 263.9367, 
    263.9786, 264.0231, 264.0242, 264.038, 264.0779, 264.0095, 264.2231, 
    264.0907, 263.8937, 263.9341, 263.9401, 263.9244, 264.0312, 263.9925, 
    264.0963, 264.0681, 264.1143, 264.0914, 264.088, 264.0585, 264.0402, 
    263.9942, 263.9565, 263.9267, 263.9336, 263.9664, 264.0258, 264.0817, 
    264.0694, 264.1108, 264.0018, 264.0472, 264.0299, 264.0757, 263.9749, 
    264.0603, 263.9529, 263.9624, 263.9917, 264.0502, 264.0635, 264.0774, 
    264.0688, 264.0274, 264.0206, 263.991, 263.9828, 263.9603, 263.9417, 
    263.9586, 263.9765, 264.0274, 264.0728, 264.1228, 264.1351, 264.1932, 
    264.1457, 264.2239, 264.1572, 264.2728, 264.0655, 264.1555, 263.9931, 
    264.0107, 264.0419, 264.1147, 264.0755, 264.1214, 264.0203, 263.9675, 
    263.9539, 263.9285, 263.9545, 263.9524, 263.9774, 263.9694, 264.0291, 
    263.997, 264.0879, 264.1211, 264.2152, 264.2728, 264.3316, 264.3575, 
    264.3654, 264.3687 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_R =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSDSND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSDSNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSDSNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSDSVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSDSVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSDSVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FSDSVILN =
  0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012 ;

 FSH =
  243.2853, 243.9773, 243.8432, 244.4004, 244.092, 244.4563, 243.4264, 
    244.0042, 243.6357, 243.3486, 245.4789, 244.4254, 246.5778, 245.9062, 
    247.6045, 246.4723, 247.8313, 247.5737, 248.353, 248.1298, 249.1232, 
    248.456, 249.6409, 248.9647, 249.0699, 248.4337, 244.639, 245.3474, 
    244.5967, 244.6978, 244.6528, 244.0977, 243.8168, 243.2336, 243.3398, 
    243.7688, 244.7433, 244.4137, 245.2477, 245.2289, 246.1544, 245.7372, 
    247.3024, 246.8514, 248.1392, 247.8173, 248.1238, 248.0311, 248.125, 
    247.653, 247.8551, 247.4404, 245.815, 246.2896, 244.8723, 244.0161, 
    243.4514, 243.0495, 243.1063, 243.2143, 243.7712, 244.2964, 244.6959, 
    244.9629, 245.2262, 246.0173, 246.4395, 247.391, 247.2223, 247.5092, 
    247.7854, 248.2471, 248.1713, 248.3744, 247.5027, 248.0815, 247.1167, 
    247.387, 245.2922, 244.5028, 244.1626, 243.8688, 243.1499, 243.646, 
    243.4503, 243.9171, 244.213, 244.0669, 244.9702, 244.6188, 246.4645, 
    245.6702, 247.7532, 247.257, 247.8723, 247.5586, 248.0956, 247.6123, 
    248.4505, 248.6323, 248.5079, 248.9877, 247.5854, 248.1232, 244.0625, 
    244.0863, 244.1978, 243.7076, 243.6779, 243.2304, 243.6291, 243.7984, 
    244.2305, 244.4849, 244.7272, 245.2599, 245.8526, 246.6828, 247.2891, 
    247.6893, 247.4443, 247.6606, 247.4186, 247.3054, 248.5638, 247.8567, 
    248.9187, 248.8601, 248.379, 248.8667, 244.1031, 243.966, 243.4883, 
    243.8622, 243.1817, 243.5619, 243.78, 244.6249, 244.8118, 244.9834, 
    245.3235, 245.7585, 246.521, 247.1943, 247.8017, 247.7573, 247.7728, 
    247.908, 247.5725, 247.9631, 248.0281, 247.8573, 248.8522, 248.568, 
    248.8589, 248.674, 244.0107, 244.2416, 244.1168, 244.3512, 244.1856, 
    244.9203, 245.1406, 246.1709, 245.7496, 246.4216, 245.8183, 245.9249, 
    246.4412, 245.8513, 247.1566, 246.2667, 247.9132, 247.022, 247.9684, 
    247.799, 248.08, 248.331, 248.6478, 249.2309, 249.0961, 249.5846, 
    244.5862, 244.8851, 244.8599, 245.1734, 245.4048, 245.9071, 246.7112, 
    246.4092, 246.9648, 247.076, 246.2325, 246.7494, 245.086, 245.354, 
    245.1953, 244.6092, 246.4774, 245.5189, 247.2988, 246.7707, 248.2951, 
    247.5403, 249.0216, 249.6523, 250.2507, 250.9444, 245.0494, 244.8462, 
    245.211, 245.7129, 246.1812, 246.8022, 246.8663, 246.9823, 247.2932, 
    247.5465, 247.0179, 247.6102, 245.414, 246.5611, 244.7684, 245.3076, 
    245.6838, 245.5199, 246.375, 246.5761, 247.4022, 246.9713, 249.4957, 
    248.3825, 251.4762, 250.6108, 244.7749, 245.0492, 246.0006, 245.5484, 
    246.8442, 247.1717, 247.4316, 247.7621, 247.7986, 247.9945, 247.6733, 
    247.9823, 246.8035, 247.3354, 245.8932, 246.2414, 246.0816, 245.9055, 
    246.4488, 247.0259, 247.0399, 247.2338, 247.7516, 246.8494, 249.6363, 
    247.9177, 245.348, 245.8728, 245.9498, 245.7462, 247.1306, 246.6288, 
    247.99, 247.6249, 248.2236, 247.9259, 247.882, 247.5002, 247.262, 
    246.6515, 246.1628, 245.7759, 245.866, 246.291, 247.0616, 247.8011, 
    247.6409, 248.1781, 246.7502, 247.3532, 247.114, 247.7235, 246.4008, 
    247.5234, 246.1156, 246.2386, 246.6189, 247.3924, 247.5641, 247.7443, 
    247.6334, 247.0814, 246.9933, 246.6101, 246.5034, 246.2119, 245.9697, 
    246.1906, 246.4222, 247.0824, 247.6857, 248.3343, 248.4937, 249.2474, 
    248.6315, 249.6456, 248.78, 250.2802, 247.5904, 248.7579, 246.6367, 
    246.8646, 247.2841, 248.2293, 247.7207, 248.3163, 246.9899, 246.3048, 
    246.1295, 245.7991, 246.1371, 246.1097, 246.4329, 246.3292, 247.1043, 
    246.688, 247.8805, 248.312, 249.5328, 250.2802, 251.0438, 251.3801, 
    251.4825, 251.5253 ;

 FSH_G =
  256.3885, 257.0815, 256.9472, 257.5051, 257.1963, 257.5611, 256.5297, 
    257.1084, 256.7394, 256.4519, 258.5851, 257.5302, 259.6856, 259.0131, 
    260.7138, 259.58, 260.9409, 260.683, 261.4634, 261.2399, 262.2347, 
    261.5665, 262.7531, 262.076, 262.1813, 261.5442, 257.7441, 258.4535, 
    257.7018, 257.803, 257.7579, 257.2021, 256.9207, 256.3367, 256.443, 
    256.8726, 257.8486, 257.5184, 258.3537, 258.3349, 259.2617, 258.8438, 
    260.4113, 259.9597, 261.2493, 260.9269, 261.2338, 261.141, 261.235, 
    260.7624, 260.9648, 260.5495, 258.9218, 259.397, 257.9777, 257.1203, 
    256.5548, 256.1523, 256.2092, 256.3173, 256.8751, 257.401, 257.8011, 
    258.0685, 258.3322, 259.1244, 259.5471, 260.5, 260.3311, 260.6184, 
    260.8949, 261.3573, 261.2814, 261.4848, 260.6118, 261.1915, 260.2254, 
    260.496, 258.3982, 257.6078, 257.267, 256.9728, 256.2528, 256.7497, 
    256.5537, 257.0212, 257.3175, 257.1712, 258.0758, 257.7239, 259.5722, 
    258.7768, 260.8627, 260.3658, 260.982, 260.6678, 261.2057, 260.7216, 
    261.561, 261.7431, 261.6185, 262.099, 260.6947, 261.2333, 257.1668, 
    257.1906, 257.3023, 256.8113, 256.7816, 256.3335, 256.7328, 256.9023, 
    257.3351, 257.5898, 257.8324, 258.3659, 258.9594, 259.7908, 260.398, 
    260.7988, 260.5534, 260.77, 260.5276, 260.4143, 261.6745, 260.9664, 
    262.0299, 261.9713, 261.4894, 261.9779, 257.2075, 257.0702, 256.5917, 
    256.9662, 256.2848, 256.6654, 256.8839, 257.73, 257.9172, 258.0891, 
    258.4296, 258.8652, 259.6288, 260.303, 260.9113, 260.8668, 260.8824, 
    261.0177, 260.6818, 261.0729, 261.138, 260.9669, 261.9633, 261.6787, 
    261.97, 261.7848, 257.115, 257.3462, 257.2212, 257.4559, 257.2901, 
    258.0258, 258.2464, 259.2782, 258.8563, 259.5293, 258.9251, 259.0318, 
    259.5488, 258.9581, 260.2653, 259.3741, 261.023, 260.1305, 261.0782, 
    260.9086, 261.19, 261.4413, 261.7586, 262.3425, 262.2076, 262.6968, 
    257.6913, 257.9906, 257.9653, 258.2794, 258.511, 259.014, 259.8193, 
    259.5169, 260.0732, 260.1846, 259.3399, 259.8575, 258.1918, 258.4602, 
    258.3012, 257.7143, 259.5851, 258.6252, 260.4077, 259.8789, 261.4054, 
    260.6495, 262.133, 262.7645, 263.3638, 264.0585, 258.1552, 257.9516, 
    258.317, 258.8195, 259.2886, 259.9104, 259.9745, 260.0907, 260.4021, 
    260.6558, 260.1264, 260.7195, 258.5202, 259.6689, 257.8737, 258.4137, 
    258.7904, 258.6263, 259.4826, 259.684, 260.5112, 260.0797, 262.6077, 
    261.493, 264.5911, 263.7245, 257.8803, 258.155, 259.1077, 258.6548, 
    259.9524, 260.2805, 260.5407, 260.8716, 260.9082, 261.1044, 260.7827, 
    261.0921, 259.9117, 260.4443, 259.0001, 259.3488, 259.1888, 259.0124, 
    259.5565, 260.1344, 260.1484, 260.3426, 260.8611, 259.9577, 262.7485, 
    261.0274, 258.4542, 258.9797, 259.0568, 258.8529, 260.2393, 259.7368, 
    261.0999, 260.7342, 261.3338, 261.0357, 260.9918, 260.6093, 260.3708, 
    259.7595, 259.2701, 258.8827, 258.9729, 259.3984, 260.1701, 260.9107, 
    260.7502, 261.2882, 259.8583, 260.4622, 260.2226, 260.833, 259.5085, 
    260.6326, 259.2228, 259.346, 259.7268, 260.5014, 260.6733, 260.8539, 
    260.7428, 260.19, 260.1017, 259.718, 259.6112, 259.3193, 259.0768, 
    259.2979, 259.5298, 260.1909, 260.7951, 261.4447, 261.6043, 262.3591, 
    261.7423, 262.7577, 261.8909, 263.3933, 260.6997, 261.8689, 259.7447, 
    259.9729, 260.3929, 261.3395, 260.8302, 261.4266, 260.0984, 259.4123, 
    259.2368, 258.9059, 259.2444, 259.2169, 259.5406, 259.4367, 260.213, 
    259.796, 260.9902, 261.4223, 262.6449, 263.3934, 264.1581, 264.4948, 
    264.5975, 264.6403 ;

 FSH_NODYNLNDUSE =
  243.2853, 243.9773, 243.8432, 244.4004, 244.092, 244.4563, 243.4264, 
    244.0042, 243.6357, 243.3486, 245.4789, 244.4254, 246.5778, 245.9062, 
    247.6045, 246.4723, 247.8313, 247.5737, 248.353, 248.1298, 249.1232, 
    248.456, 249.6409, 248.9647, 249.0699, 248.4337, 244.639, 245.3474, 
    244.5967, 244.6978, 244.6528, 244.0977, 243.8168, 243.2336, 243.3398, 
    243.7688, 244.7433, 244.4137, 245.2477, 245.2289, 246.1544, 245.7372, 
    247.3024, 246.8514, 248.1392, 247.8173, 248.1238, 248.0311, 248.125, 
    247.653, 247.8551, 247.4404, 245.815, 246.2896, 244.8723, 244.0161, 
    243.4514, 243.0495, 243.1063, 243.2143, 243.7712, 244.2964, 244.6959, 
    244.9629, 245.2262, 246.0173, 246.4395, 247.391, 247.2223, 247.5092, 
    247.7854, 248.2471, 248.1713, 248.3744, 247.5027, 248.0815, 247.1167, 
    247.387, 245.2922, 244.5028, 244.1626, 243.8688, 243.1499, 243.646, 
    243.4503, 243.9171, 244.213, 244.0669, 244.9702, 244.6188, 246.4645, 
    245.6702, 247.7532, 247.257, 247.8723, 247.5586, 248.0956, 247.6123, 
    248.4505, 248.6323, 248.5079, 248.9877, 247.5854, 248.1232, 244.0625, 
    244.0863, 244.1978, 243.7076, 243.6779, 243.2304, 243.6291, 243.7984, 
    244.2305, 244.4849, 244.7272, 245.2599, 245.8526, 246.6828, 247.2891, 
    247.6893, 247.4443, 247.6606, 247.4186, 247.3054, 248.5638, 247.8567, 
    248.9187, 248.8601, 248.379, 248.8667, 244.1031, 243.966, 243.4883, 
    243.8622, 243.1817, 243.5619, 243.78, 244.6249, 244.8118, 244.9834, 
    245.3235, 245.7585, 246.521, 247.1943, 247.8017, 247.7573, 247.7728, 
    247.908, 247.5725, 247.9631, 248.0281, 247.8573, 248.8522, 248.568, 
    248.8589, 248.674, 244.0107, 244.2416, 244.1168, 244.3512, 244.1856, 
    244.9203, 245.1406, 246.1709, 245.7496, 246.4216, 245.8183, 245.9249, 
    246.4412, 245.8513, 247.1566, 246.2667, 247.9132, 247.022, 247.9684, 
    247.799, 248.08, 248.331, 248.6478, 249.2309, 249.0961, 249.5846, 
    244.5862, 244.8851, 244.8599, 245.1734, 245.4048, 245.9071, 246.7112, 
    246.4092, 246.9648, 247.076, 246.2325, 246.7494, 245.086, 245.354, 
    245.1953, 244.6092, 246.4774, 245.5189, 247.2988, 246.7707, 248.2951, 
    247.5403, 249.0216, 249.6523, 250.2507, 250.9444, 245.0494, 244.8462, 
    245.211, 245.7129, 246.1812, 246.8022, 246.8663, 246.9823, 247.2932, 
    247.5465, 247.0179, 247.6102, 245.414, 246.5611, 244.7684, 245.3076, 
    245.6838, 245.5199, 246.375, 246.5761, 247.4022, 246.9713, 249.4957, 
    248.3825, 251.4762, 250.6108, 244.7749, 245.0492, 246.0006, 245.5484, 
    246.8442, 247.1717, 247.4316, 247.7621, 247.7986, 247.9945, 247.6733, 
    247.9823, 246.8035, 247.3354, 245.8932, 246.2414, 246.0816, 245.9055, 
    246.4488, 247.0259, 247.0399, 247.2338, 247.7516, 246.8494, 249.6363, 
    247.9177, 245.348, 245.8728, 245.9498, 245.7462, 247.1306, 246.6288, 
    247.99, 247.6249, 248.2236, 247.9259, 247.882, 247.5002, 247.262, 
    246.6515, 246.1628, 245.7759, 245.866, 246.291, 247.0616, 247.8011, 
    247.6409, 248.1781, 246.7502, 247.3532, 247.114, 247.7235, 246.4008, 
    247.5234, 246.1156, 246.2386, 246.6189, 247.3924, 247.5641, 247.7443, 
    247.6334, 247.0814, 246.9933, 246.6101, 246.5034, 246.2119, 245.9697, 
    246.1906, 246.4222, 247.0824, 247.6857, 248.3343, 248.4937, 249.2474, 
    248.6315, 249.6456, 248.78, 250.2802, 247.5904, 248.7579, 246.6367, 
    246.8646, 247.2841, 248.2293, 247.7207, 248.3163, 246.9899, 246.3048, 
    246.1295, 245.7991, 246.1371, 246.1097, 246.4329, 246.3292, 247.1043, 
    246.688, 247.8805, 248.312, 249.5328, 250.2802, 251.0438, 251.3801, 
    251.4825, 251.5253 ;

 FSH_R =
  243.2853, 243.9773, 243.8432, 244.4004, 244.092, 244.4563, 243.4264, 
    244.0042, 243.6357, 243.3486, 245.4789, 244.4254, 246.5778, 245.9062, 
    247.6045, 246.4723, 247.8313, 247.5737, 248.353, 248.1298, 249.1232, 
    248.456, 249.6409, 248.9647, 249.0699, 248.4337, 244.639, 245.3474, 
    244.5967, 244.6978, 244.6528, 244.0977, 243.8168, 243.2336, 243.3398, 
    243.7688, 244.7433, 244.4137, 245.2477, 245.2289, 246.1544, 245.7372, 
    247.3024, 246.8514, 248.1392, 247.8173, 248.1238, 248.0311, 248.125, 
    247.653, 247.8551, 247.4404, 245.815, 246.2896, 244.8723, 244.0161, 
    243.4514, 243.0495, 243.1063, 243.2143, 243.7712, 244.2964, 244.6959, 
    244.9629, 245.2262, 246.0173, 246.4395, 247.391, 247.2223, 247.5092, 
    247.7854, 248.2471, 248.1713, 248.3744, 247.5027, 248.0815, 247.1167, 
    247.387, 245.2922, 244.5028, 244.1626, 243.8688, 243.1499, 243.646, 
    243.4503, 243.9171, 244.213, 244.0669, 244.9702, 244.6188, 246.4645, 
    245.6702, 247.7532, 247.257, 247.8723, 247.5586, 248.0956, 247.6123, 
    248.4505, 248.6323, 248.5079, 248.9877, 247.5854, 248.1232, 244.0625, 
    244.0863, 244.1978, 243.7076, 243.6779, 243.2304, 243.6291, 243.7984, 
    244.2305, 244.4849, 244.7272, 245.2599, 245.8526, 246.6828, 247.2891, 
    247.6893, 247.4443, 247.6606, 247.4186, 247.3054, 248.5638, 247.8567, 
    248.9187, 248.8601, 248.379, 248.8667, 244.1031, 243.966, 243.4883, 
    243.8622, 243.1817, 243.5619, 243.78, 244.6249, 244.8118, 244.9834, 
    245.3235, 245.7585, 246.521, 247.1943, 247.8017, 247.7573, 247.7728, 
    247.908, 247.5725, 247.9631, 248.0281, 247.8573, 248.8522, 248.568, 
    248.8589, 248.674, 244.0107, 244.2416, 244.1168, 244.3512, 244.1856, 
    244.9203, 245.1406, 246.1709, 245.7496, 246.4216, 245.8183, 245.9249, 
    246.4412, 245.8513, 247.1566, 246.2667, 247.9132, 247.022, 247.9684, 
    247.799, 248.08, 248.331, 248.6478, 249.2309, 249.0961, 249.5846, 
    244.5862, 244.8851, 244.8599, 245.1734, 245.4048, 245.9071, 246.7112, 
    246.4092, 246.9648, 247.076, 246.2325, 246.7494, 245.086, 245.354, 
    245.1953, 244.6092, 246.4774, 245.5189, 247.2988, 246.7707, 248.2951, 
    247.5403, 249.0216, 249.6523, 250.2507, 250.9444, 245.0494, 244.8462, 
    245.211, 245.7129, 246.1812, 246.8022, 246.8663, 246.9823, 247.2932, 
    247.5465, 247.0179, 247.6102, 245.414, 246.5611, 244.7684, 245.3076, 
    245.6838, 245.5199, 246.375, 246.5761, 247.4022, 246.9713, 249.4957, 
    248.3825, 251.4762, 250.6108, 244.7749, 245.0492, 246.0006, 245.5484, 
    246.8442, 247.1717, 247.4316, 247.7621, 247.7986, 247.9945, 247.6733, 
    247.9823, 246.8035, 247.3354, 245.8932, 246.2414, 246.0816, 245.9055, 
    246.4488, 247.0259, 247.0399, 247.2338, 247.7516, 246.8494, 249.6363, 
    247.9177, 245.348, 245.8728, 245.9498, 245.7462, 247.1306, 246.6288, 
    247.99, 247.6249, 248.2236, 247.9259, 247.882, 247.5002, 247.262, 
    246.6515, 246.1628, 245.7759, 245.866, 246.291, 247.0616, 247.8011, 
    247.6409, 248.1781, 246.7502, 247.3532, 247.114, 247.7235, 246.4008, 
    247.5234, 246.1156, 246.2386, 246.6189, 247.3924, 247.5641, 247.7443, 
    247.6334, 247.0814, 246.9933, 246.6101, 246.5034, 246.2119, 245.9697, 
    246.1906, 246.4222, 247.0824, 247.6857, 248.3343, 248.4937, 249.2474, 
    248.6315, 249.6456, 248.78, 250.2802, 247.5904, 248.7579, 246.6367, 
    246.8646, 247.2841, 248.2293, 247.7207, 248.3163, 246.9899, 246.3048, 
    246.1295, 245.7991, 246.1371, 246.1097, 246.4329, 246.3292, 247.1043, 
    246.688, 247.8805, 248.312, 249.5328, 250.2802, 251.0438, 251.3801, 
    251.4825, 251.5253 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -13.10316, -13.10416, -13.10397, -13.10477, -13.10433, -13.10485, 
    -13.10337, -13.10419, -13.10368, -13.10326, -13.10628, -13.1048, 
    -13.10787, -13.10693, -13.1093, -13.10771, -13.10963, -13.10928, 
    -13.11039, -13.11007, -13.11147, -13.11054, -13.11223, -13.11126, 
    -13.1114, -13.11051, -13.10512, -13.10609, -13.10506, -13.1052, 
    -13.10514, -13.10433, -13.10392, -13.1031, -13.10325, -13.10386, 
    -13.10526, -13.1048, -13.10601, -13.10598, -13.10728, -13.1067, 
    -13.10889, -13.10828, -13.11009, -13.10963, -13.11006, -13.10993, 
    -13.11007, -13.10939, -13.10968, -13.10909, -13.1068, -13.10747, 
    -13.10545, -13.10419, -13.10341, -13.10283, -13.10291, -13.10307, 
    -13.10386, -13.10463, -13.10521, -13.10559, -13.10598, -13.10706, 
    -13.10767, -13.10901, -13.10878, -13.10918, -13.10958, -13.11024, 
    -13.11013, -13.11042, -13.10918, -13.11, -13.10866, -13.10901, -13.10601, 
    -13.10493, -13.10441, -13.10401, -13.10298, -13.10368, -13.1034, 
    -13.10408, -13.10451, -13.1043, -13.10561, -13.10509, -13.10771, 
    -13.10659, -13.10953, -13.10883, -13.10971, -13.10926, -13.11002, 
    -13.10934, -13.11053, -13.11078, -13.11061, -13.1113, -13.1093, 
    -13.11006, -13.10429, -13.10433, -13.10449, -13.10377, -13.10373, 
    -13.10309, -13.10367, -13.1039, -13.10454, -13.1049, -13.10525, 
    -13.10602, -13.10685, -13.10802, -13.10887, -13.10945, -13.1091, 
    -13.10941, -13.10906, -13.1089, -13.11068, -13.10968, -13.1112, 
    -13.11112, -13.11042, -13.11113, -13.10435, -13.10416, -13.10346, 
    -13.10401, -13.10302, -13.10357, -13.10387, -13.10509, -13.10538, 
    -13.10562, -13.10611, -13.10673, -13.1078, -13.10873, -13.10961, 
    -13.10954, -13.10957, -13.10976, -13.10928, -13.10983, -13.10992, 
    -13.10968, -13.11111, -13.1107, -13.11112, -13.11085, -13.10422, 
    -13.10455, -13.10437, -13.1047, -13.10446, -13.10551, -13.10583, 
    -13.10729, -13.10671, -13.10765, -13.10681, -13.10696, -13.10766, 
    -13.10686, -13.10867, -13.10742, -13.10976, -13.10848, -13.10984, 
    -13.1096, -13.11, -13.11036, -13.11081, -13.11164, -13.11145, -13.11216, 
    -13.10505, -13.10547, -13.10545, -13.1059, -13.10622, -13.10694, 
    -13.10807, -13.10765, -13.10844, -13.10859, -13.1074, -13.10812, 
    -13.10576, -13.10614, -13.10593, -13.10507, -13.10773, -13.10637, 
    -13.10888, -13.10816, -13.11031, -13.10922, -13.11135, -13.11223, 
    -13.11312, -13.1141, -13.10572, -13.10543, -13.10596, -13.10665, 
    -13.10732, -13.1082, -13.1083, -13.10846, -13.10888, -13.10924, -13.1085, 
    -13.10933, -13.1062, -13.10785, -13.10531, -13.10607, -13.10661, 
    -13.10639, -13.1076, -13.10789, -13.10903, -13.10845, -13.112, -13.11041, 
    -13.1149, -13.11363, -13.10532, -13.10572, -13.10706, -13.10643, 
    -13.10827, -13.10871, -13.10908, -13.10954, -13.1096, -13.10988, 
    -13.10942, -13.10986, -13.1082, -13.10894, -13.10692, -13.10741, 
    -13.10719, -13.10694, -13.10771, -13.10851, -13.10854, -13.10879, 
    -13.10947, -13.10827, -13.11217, -13.10971, -13.10615, -13.10687, 
    -13.107, -13.10671, -13.10867, -13.10796, -13.10987, -13.10935, 
    -13.11021, -13.10978, -13.10972, -13.10918, -13.10884, -13.10799, 
    -13.1073, -13.10676, -13.10688, -13.10748, -13.10856, -13.1096, 
    -13.10936, -13.11014, -13.10813, -13.10896, -13.10864, -13.10949, 
    -13.10763, -13.10915, -13.10724, -13.10741, -13.10794, -13.109, 
    -13.10927, -13.10952, -13.10937, -13.10859, -13.10847, -13.10793, 
    -13.10778, -13.10737, -13.10703, -13.10734, -13.10766, -13.1086, 
    -13.10943, -13.11036, -13.11059, -13.11163, -13.11076, -13.11218, 
    -13.11093, -13.11312, -13.10927, -13.11093, -13.10797, -13.1083, 
    -13.10885, -13.11019, -13.10949, -13.11032, -13.10847, -13.10749, 
    -13.10726, -13.10679, -13.10727, -13.10723, -13.10769, -13.10754, 
    -13.10863, -13.10805, -13.10971, -13.11032, -13.11207, -13.11315, 
    -13.11427, -13.11476, -13.11491, -13.11498 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531 ;

 FSRND =
  0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151 ;

 FSRNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSRNI =
  0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505 ;

 FSRVD =
  0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803 ;

 FSRVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSRVI =
  0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  2.809604e-14, 2.822128e-14, 2.819686e-14, 2.829796e-14, 2.824182e-14, 
    2.830801e-14, 2.812127e-14, 2.822611e-14, 2.815912e-14, 2.810706e-14, 
    2.849423e-14, 2.830228e-14, 2.869358e-14, 2.857098e-14, 2.88789e-14, 
    2.867447e-14, 2.892011e-14, 2.887287e-14, 2.901481e-14, 2.897409e-14, 
    2.915586e-14, 2.903352e-14, 2.925002e-14, 2.912656e-14, 2.914586e-14, 
    2.902938e-14, 2.8341e-14, 2.847052e-14, 2.83333e-14, 2.835176e-14, 
    2.834343e-14, 2.82429e-14, 2.81923e-14, 2.80862e-14, 2.810541e-14, 
    2.81833e-14, 2.835988e-14, 2.829983e-14, 2.845097e-14, 2.844756e-14, 
    2.861602e-14, 2.854003e-14, 2.882342e-14, 2.874277e-14, 2.897576e-14, 
    2.891711e-14, 2.897297e-14, 2.895598e-14, 2.897312e-14, 2.888716e-14, 
    2.892394e-14, 2.88483e-14, 2.855456e-14, 2.864098e-14, 2.838328e-14, 
    2.822859e-14, 2.812577e-14, 2.805293e-14, 2.806317e-14, 2.808282e-14, 
    2.81837e-14, 2.827855e-14, 2.835091e-14, 2.83993e-14, 2.8447e-14, 
    2.859172e-14, 2.86682e-14, 2.88397e-14, 2.880867e-14, 2.886115e-14, 
    2.891125e-14, 2.899544e-14, 2.898155e-14, 2.901864e-14, 2.885959e-14, 
    2.896528e-14, 2.87908e-14, 2.88385e-14, 2.846044e-14, 2.831612e-14, 
    2.8255e-14, 2.820134e-14, 2.807108e-14, 2.816101e-14, 2.812553e-14, 
    2.820981e-14, 2.826342e-14, 2.823685e-14, 2.84006e-14, 2.833688e-14, 
    2.86727e-14, 2.852796e-14, 2.890543e-14, 2.881498e-14, 2.892703e-14, 
    2.886982e-14, 2.896783e-14, 2.887958e-14, 2.90324e-14, 2.906573e-14, 
    2.90429e-14, 2.913032e-14, 2.887454e-14, 2.897274e-14, 2.823626e-14, 
    2.82406e-14, 2.826071e-14, 2.817215e-14, 2.816671e-14, 2.808554e-14, 
    2.815768e-14, 2.818845e-14, 2.826645e-14, 2.831263e-14, 2.835653e-14, 
    2.845316e-14, 2.856115e-14, 2.871222e-14, 2.882081e-14, 2.889362e-14, 
    2.884892e-14, 2.888834e-14, 2.884423e-14, 2.882352e-14, 2.905318e-14, 
    2.89242e-14, 2.911768e-14, 2.910696e-14, 2.901934e-14, 2.91081e-14, 
    2.824358e-14, 2.821864e-14, 2.813227e-14, 2.819981e-14, 2.807665e-14, 
    2.814559e-14, 2.818523e-14, 2.833823e-14, 2.837179e-14, 2.840301e-14, 
    2.846461e-14, 2.854373e-14, 2.868267e-14, 2.88036e-14, 2.891405e-14, 
    2.890591e-14, 2.890875e-14, 2.893342e-14, 2.887225e-14, 2.894341e-14, 
    2.895535e-14, 2.892409e-14, 2.910545e-14, 2.905361e-14, 2.910663e-14, 
    2.907283e-14, 2.82267e-14, 2.826856e-14, 2.824589e-14, 2.828848e-14, 
    2.825844e-14, 2.839187e-14, 2.843186e-14, 2.861918e-14, 2.854218e-14, 
    2.866464e-14, 2.855455e-14, 2.857406e-14, 2.866864e-14, 2.856042e-14, 
    2.879689e-14, 2.863656e-14, 2.893435e-14, 2.877422e-14, 2.894435e-14, 
    2.891337e-14, 2.896455e-14, 2.901045e-14, 2.906811e-14, 2.917472e-14, 
    2.914996e-14, 2.923912e-14, 2.833099e-14, 2.838535e-14, 2.838051e-14, 
    2.843739e-14, 2.847947e-14, 2.857074e-14, 2.871724e-14, 2.866207e-14, 
    2.876322e-14, 2.878356e-14, 2.862977e-14, 2.872418e-14, 2.842148e-14, 
    2.847035e-14, 2.844119e-14, 2.833492e-14, 2.867462e-14, 2.850018e-14, 
    2.882232e-14, 2.872769e-14, 2.900383e-14, 2.886648e-14, 2.913636e-14, 
    2.925198e-14, 2.936063e-14, 2.948788e-14, 2.841497e-14, 2.837797e-14, 
    2.844409e-14, 2.853575e-14, 2.862067e-14, 2.873376e-14, 2.874528e-14, 
    2.876645e-14, 2.882132e-14, 2.886751e-14, 2.877314e-14, 2.887902e-14, 
    2.848174e-14, 2.868974e-14, 2.836371e-14, 2.846187e-14, 2.852998e-14, 
    2.850004e-14, 2.865544e-14, 2.869207e-14, 2.884114e-14, 2.876403e-14, 
    2.92234e-14, 2.902002e-14, 2.958466e-14, 2.942673e-14, 2.836504e-14, 
    2.841472e-14, 2.858792e-14, 2.850547e-14, 2.874122e-14, 2.879934e-14, 
    2.88465e-14, 2.890694e-14, 2.891339e-14, 2.894921e-14, 2.889047e-14, 
    2.894683e-14, 2.873374e-14, 2.882891e-14, 2.856779e-14, 2.863129e-14, 
    2.860203e-14, 2.856995e-14, 2.866884e-14, 2.877435e-14, 2.877651e-14, 
    2.881033e-14, 2.890587e-14, 2.874172e-14, 2.924969e-14, 2.893589e-14, 
    2.846894e-14, 2.856483e-14, 2.857843e-14, 2.854128e-14, 2.879344e-14, 
    2.870203e-14, 2.894833e-14, 2.888167e-14, 2.899079e-14, 2.893655e-14, 
    2.892852e-14, 2.885887e-14, 2.881548e-14, 2.870603e-14, 2.861695e-14, 
    2.854637e-14, 2.856272e-14, 2.864028e-14, 2.878072e-14, 2.89137e-14, 
    2.888454e-14, 2.898217e-14, 2.872361e-14, 2.883201e-14, 2.879007e-14, 
    2.889929e-14, 2.866052e-14, 2.886447e-14, 2.860843e-14, 2.86308e-14, 
    2.870014e-14, 2.883978e-14, 2.887054e-14, 2.890357e-14, 2.888313e-14, 
    2.878446e-14, 2.876824e-14, 2.869827e-14, 2.867897e-14, 2.86257e-14, 
    2.858157e-14, 2.862186e-14, 2.866412e-14, 2.878428e-14, 2.889263e-14, 
    2.90108e-14, 2.903971e-14, 2.917806e-14, 2.906547e-14, 2.925133e-14, 
    2.90934e-14, 2.936673e-14, 2.887613e-14, 2.908913e-14, 2.870328e-14, 
    2.874475e-14, 2.881992e-14, 2.899227e-14, 2.889908e-14, 2.900801e-14, 
    2.876758e-14, 2.864303e-14, 2.861071e-14, 2.855063e-14, 2.861204e-14, 
    2.860704e-14, 2.866584e-14, 2.864689e-14, 2.87882e-14, 2.871227e-14, 
    2.8928e-14, 2.900684e-14, 2.922951e-14, 2.936615e-14, 2.950526e-14, 
    2.95667e-14, 2.95854e-14, 2.95932e-14 ;

 F_DENIT_vr =
  1.604313e-12, 1.611464e-12, 1.61007e-12, 1.615843e-12, 1.612637e-12, 
    1.616417e-12, 1.605754e-12, 1.61174e-12, 1.607915e-12, 1.604942e-12, 
    1.62705e-12, 1.616089e-12, 1.638433e-12, 1.631433e-12, 1.649015e-12, 
    1.637342e-12, 1.651368e-12, 1.648671e-12, 1.656776e-12, 1.654451e-12, 
    1.66483e-12, 1.657844e-12, 1.670206e-12, 1.663157e-12, 1.664259e-12, 
    1.657607e-12, 1.618301e-12, 1.625696e-12, 1.617861e-12, 1.618915e-12, 
    1.618439e-12, 1.612698e-12, 1.60981e-12, 1.603751e-12, 1.604848e-12, 
    1.609295e-12, 1.619378e-12, 1.615949e-12, 1.62458e-12, 1.624385e-12, 
    1.634004e-12, 1.629665e-12, 1.645847e-12, 1.641242e-12, 1.654546e-12, 
    1.651197e-12, 1.654386e-12, 1.653416e-12, 1.654395e-12, 1.649487e-12, 
    1.651587e-12, 1.647268e-12, 1.630495e-12, 1.635429e-12, 1.620715e-12, 
    1.611882e-12, 1.606011e-12, 1.601851e-12, 1.602436e-12, 1.603558e-12, 
    1.609318e-12, 1.614734e-12, 1.618866e-12, 1.62163e-12, 1.624353e-12, 
    1.632617e-12, 1.636984e-12, 1.646777e-12, 1.645005e-12, 1.648001e-12, 
    1.650862e-12, 1.655669e-12, 1.654877e-12, 1.656994e-12, 1.647913e-12, 
    1.653948e-12, 1.643984e-12, 1.646708e-12, 1.62512e-12, 1.61688e-12, 
    1.61339e-12, 1.610325e-12, 1.602888e-12, 1.608023e-12, 1.605997e-12, 
    1.610809e-12, 1.613871e-12, 1.612353e-12, 1.621704e-12, 1.618065e-12, 
    1.637241e-12, 1.628976e-12, 1.65053e-12, 1.645365e-12, 1.651763e-12, 
    1.648497e-12, 1.654093e-12, 1.649054e-12, 1.65778e-12, 1.659683e-12, 
    1.65838e-12, 1.663372e-12, 1.648766e-12, 1.654373e-12, 1.61232e-12, 
    1.612567e-12, 1.613716e-12, 1.608659e-12, 1.608348e-12, 1.603713e-12, 
    1.607833e-12, 1.609589e-12, 1.614044e-12, 1.61668e-12, 1.619187e-12, 
    1.624705e-12, 1.630871e-12, 1.639497e-12, 1.645698e-12, 1.649855e-12, 
    1.647303e-12, 1.649554e-12, 1.647035e-12, 1.645853e-12, 1.658967e-12, 
    1.651601e-12, 1.662649e-12, 1.662038e-12, 1.657034e-12, 1.662102e-12, 
    1.612738e-12, 1.611314e-12, 1.606382e-12, 1.610239e-12, 1.603206e-12, 
    1.607142e-12, 1.609406e-12, 1.618142e-12, 1.620058e-12, 1.621841e-12, 
    1.625359e-12, 1.629876e-12, 1.63781e-12, 1.644715e-12, 1.651022e-12, 
    1.650557e-12, 1.65072e-12, 1.652128e-12, 1.648635e-12, 1.652699e-12, 
    1.653381e-12, 1.651595e-12, 1.661952e-12, 1.658991e-12, 1.662019e-12, 
    1.660089e-12, 1.611774e-12, 1.614164e-12, 1.61287e-12, 1.615301e-12, 
    1.613586e-12, 1.621205e-12, 1.623489e-12, 1.634185e-12, 1.629788e-12, 
    1.636781e-12, 1.630494e-12, 1.631608e-12, 1.637009e-12, 1.630829e-12, 
    1.644332e-12, 1.635177e-12, 1.652182e-12, 1.643037e-12, 1.652752e-12, 
    1.650983e-12, 1.653905e-12, 1.656526e-12, 1.659819e-12, 1.665907e-12, 
    1.664493e-12, 1.669584e-12, 1.617729e-12, 1.620833e-12, 1.620556e-12, 
    1.623804e-12, 1.626207e-12, 1.631419e-12, 1.639784e-12, 1.636634e-12, 
    1.64241e-12, 1.643571e-12, 1.634789e-12, 1.640181e-12, 1.622896e-12, 
    1.625686e-12, 1.624021e-12, 1.617953e-12, 1.637351e-12, 1.62739e-12, 
    1.645784e-12, 1.640381e-12, 1.656149e-12, 1.648306e-12, 1.663716e-12, 
    1.670318e-12, 1.676522e-12, 1.683788e-12, 1.622524e-12, 1.620411e-12, 
    1.624187e-12, 1.629421e-12, 1.63427e-12, 1.640728e-12, 1.641385e-12, 
    1.642594e-12, 1.645727e-12, 1.648365e-12, 1.642976e-12, 1.649022e-12, 
    1.626337e-12, 1.638214e-12, 1.619597e-12, 1.625202e-12, 1.629091e-12, 
    1.627382e-12, 1.636255e-12, 1.638347e-12, 1.646859e-12, 1.642456e-12, 
    1.668686e-12, 1.657073e-12, 1.689315e-12, 1.680297e-12, 1.619673e-12, 
    1.62251e-12, 1.6324e-12, 1.627692e-12, 1.641153e-12, 1.644472e-12, 
    1.647165e-12, 1.650616e-12, 1.650984e-12, 1.65303e-12, 1.649676e-12, 
    1.652894e-12, 1.640726e-12, 1.64616e-12, 1.63125e-12, 1.634876e-12, 
    1.633206e-12, 1.631374e-12, 1.63702e-12, 1.643045e-12, 1.643169e-12, 
    1.6451e-12, 1.650555e-12, 1.641182e-12, 1.670187e-12, 1.652269e-12, 
    1.625606e-12, 1.631082e-12, 1.631858e-12, 1.629737e-12, 1.644135e-12, 
    1.638915e-12, 1.652979e-12, 1.649173e-12, 1.655404e-12, 1.652307e-12, 
    1.651848e-12, 1.647871e-12, 1.645394e-12, 1.639144e-12, 1.634058e-12, 
    1.630027e-12, 1.630961e-12, 1.635389e-12, 1.643409e-12, 1.651002e-12, 
    1.649337e-12, 1.654912e-12, 1.640148e-12, 1.646338e-12, 1.643943e-12, 
    1.65018e-12, 1.636545e-12, 1.648191e-12, 1.633571e-12, 1.634849e-12, 
    1.638808e-12, 1.646782e-12, 1.648538e-12, 1.650424e-12, 1.649256e-12, 
    1.643623e-12, 1.642696e-12, 1.638701e-12, 1.637599e-12, 1.634557e-12, 
    1.632037e-12, 1.634338e-12, 1.636751e-12, 1.643612e-12, 1.649799e-12, 
    1.656547e-12, 1.658197e-12, 1.666097e-12, 1.659669e-12, 1.670281e-12, 
    1.661263e-12, 1.676871e-12, 1.648857e-12, 1.66102e-12, 1.638987e-12, 
    1.641355e-12, 1.645647e-12, 1.655489e-12, 1.650168e-12, 1.656387e-12, 
    1.642659e-12, 1.635546e-12, 1.633701e-12, 1.630271e-12, 1.633777e-12, 
    1.633492e-12, 1.636849e-12, 1.635767e-12, 1.643836e-12, 1.6395e-12, 
    1.651819e-12, 1.65632e-12, 1.669035e-12, 1.676838e-12, 1.684781e-12, 
    1.688289e-12, 1.689357e-12, 1.689802e-12,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  7.549451e-16, 7.557162e-16, 7.555651e-16, 7.561827e-16, 7.558394e-16, 
    7.562421e-16, 7.55098e-16, 7.557428e-16, 7.553305e-16, 7.550081e-16, 
    7.573603e-16, 7.562047e-16, 7.585288e-16, 7.578091e-16, 7.595942e-16, 
    7.58417e-16, 7.598275e-16, 7.595569e-16, 7.603594e-16, 7.601295e-16, 
    7.611465e-16, 7.60463e-16, 7.616621e-16, 7.609819e-16, 7.610887e-16, 
    7.604374e-16, 7.564418e-16, 7.572232e-16, 7.563943e-16, 7.565065e-16, 
    7.564549e-16, 7.558443e-16, 7.555358e-16, 7.548784e-16, 7.549968e-16, 
    7.554782e-16, 7.565519e-16, 7.56187e-16, 7.570955e-16, 7.570752e-16, 
    7.580716e-16, 7.57624e-16, 7.592736e-16, 7.588079e-16, 7.601383e-16, 
    7.598059e-16, 7.601218e-16, 7.600249e-16, 7.601212e-16, 7.596344e-16, 
    7.598422e-16, 7.594114e-16, 7.577162e-16, 7.582236e-16, 7.56695e-16, 
    7.557588e-16, 7.55124e-16, 7.546718e-16, 7.547345e-16, 7.548572e-16, 
    7.554796e-16, 7.560574e-16, 7.564951e-16, 7.567857e-16, 7.570704e-16, 
    7.579316e-16, 7.583773e-16, 7.593666e-16, 7.591872e-16, 7.594879e-16, 
    7.59772e-16, 7.602474e-16, 7.601687e-16, 7.603769e-16, 7.594754e-16, 
    7.600764e-16, 7.590796e-16, 7.59354e-16, 7.57161e-16, 7.56288e-16, 
    7.55919e-16, 7.555884e-16, 7.547835e-16, 7.553404e-16, 7.551208e-16, 
    7.556375e-16, 7.559649e-16, 7.558017e-16, 7.567929e-16, 7.564086e-16, 
    7.584026e-16, 7.575517e-16, 7.597398e-16, 7.592224e-16, 7.598607e-16, 
    7.595353e-16, 7.60091e-16, 7.5959e-16, 7.604527e-16, 7.6064e-16, 
    7.605109e-16, 7.609976e-16, 7.595582e-16, 7.601159e-16, 7.558014e-16, 
    7.55828e-16, 7.559497e-16, 7.554082e-16, 7.553742e-16, 7.548714e-16, 
    7.553167e-16, 7.555064e-16, 7.559816e-16, 7.562616e-16, 7.565263e-16, 
    7.571061e-16, 7.577471e-16, 7.5863e-16, 7.592553e-16, 7.596701e-16, 
    7.594148e-16, 7.596391e-16, 7.593872e-16, 7.592675e-16, 7.605685e-16, 
    7.598421e-16, 7.60926e-16, 7.608664e-16, 7.603771e-16, 7.608713e-16, 
    7.558452e-16, 7.556917e-16, 7.551613e-16, 7.555755e-16, 7.548151e-16, 
    7.552424e-16, 7.554863e-16, 7.564171e-16, 7.566175e-16, 7.568057e-16, 
    7.571731e-16, 7.57642e-16, 7.584575e-16, 7.591559e-16, 7.597856e-16, 
    7.597385e-16, 7.597545e-16, 7.59894e-16, 7.59546e-16, 7.599495e-16, 
    7.600169e-16, 7.598394e-16, 7.608566e-16, 7.605676e-16, 7.608625e-16, 
    7.606733e-16, 7.557404e-16, 7.559952e-16, 7.558564e-16, 7.561161e-16, 
    7.559324e-16, 7.567407e-16, 7.5698e-16, 7.580884e-16, 7.576331e-16, 
    7.58353e-16, 7.577049e-16, 7.578205e-16, 7.583769e-16, 7.577378e-16, 
    7.591168e-16, 7.581868e-16, 7.598987e-16, 7.589857e-16, 7.599542e-16, 
    7.597775e-16, 7.600665e-16, 7.603257e-16, 7.606472e-16, 7.612399e-16, 
    7.611016e-16, 7.615924e-16, 7.563733e-16, 7.56701e-16, 7.566706e-16, 
    7.570111e-16, 7.572617e-16, 7.578019e-16, 7.586582e-16, 7.58336e-16, 
    7.589221e-16, 7.590398e-16, 7.581453e-16, 7.586966e-16, 7.569123e-16, 
    7.572044e-16, 7.570289e-16, 7.563898e-16, 7.584064e-16, 7.573797e-16, 
    7.59258e-16, 7.587117e-16, 7.602871e-16, 7.595103e-16, 7.610259e-16, 
    7.616647e-16, 7.622521e-16, 7.629364e-16, 7.568776e-16, 7.566542e-16, 
    7.570499e-16, 7.575965e-16, 7.580943e-16, 7.587532e-16, 7.588186e-16, 
    7.589405e-16, 7.592549e-16, 7.595194e-16, 7.589788e-16, 7.595835e-16, 
    7.572739e-16, 7.584938e-16, 7.565624e-16, 7.571522e-16, 7.575547e-16, 
    7.573767e-16, 7.582903e-16, 7.585031e-16, 7.593635e-16, 7.589194e-16, 
    7.61507e-16, 7.603772e-16, 7.634466e-16, 7.626081e-16, 7.565759e-16, 
    7.568735e-16, 7.579023e-16, 7.574145e-16, 7.587943e-16, 7.5913e-16, 
    7.593987e-16, 7.597443e-16, 7.597791e-16, 7.599826e-16, 7.596477e-16, 
    7.599677e-16, 7.587476e-16, 7.592954e-16, 7.577768e-16, 7.581497e-16, 
    7.579772e-16, 7.577878e-16, 7.583668e-16, 7.589803e-16, 7.589905e-16, 
    7.59185e-16, 7.597357e-16, 7.587877e-16, 7.616522e-16, 7.599034e-16, 
    7.571968e-16, 7.577665e-16, 7.578443e-16, 7.576248e-16, 7.590946e-16, 
    7.585663e-16, 7.599773e-16, 7.595979e-16, 7.602152e-16, 7.599092e-16, 
    7.598627e-16, 7.594663e-16, 7.59217e-16, 7.585858e-16, 7.580648e-16, 
    7.576486e-16, 7.577441e-16, 7.582006e-16, 7.590152e-16, 7.597752e-16, 
    7.59609e-16, 7.601602e-16, 7.58682e-16, 7.593075e-16, 7.590658e-16, 
    7.596898e-16, 7.583251e-16, 7.595071e-16, 7.580191e-16, 7.581496e-16, 
    7.585538e-16, 7.593609e-16, 7.595334e-16, 7.597223e-16, 7.596041e-16, 
    7.590403e-16, 7.589456e-16, 7.585392e-16, 7.584268e-16, 7.581149e-16, 
    7.578548e-16, 7.580918e-16, 7.583386e-16, 7.590345e-16, 7.596545e-16, 
    7.603217e-16, 7.604829e-16, 7.612547e-16, 7.606289e-16, 7.61659e-16, 
    7.607874e-16, 7.622833e-16, 7.5957e-16, 7.60771e-16, 7.585716e-16, 
    7.588112e-16, 7.592457e-16, 7.602247e-16, 7.596949e-16, 7.603122e-16, 
    7.589413e-16, 7.582184e-16, 7.580268e-16, 7.576735e-16, 7.580336e-16, 
    7.580043e-16, 7.583475e-16, 7.58236e-16, 7.590556e-16, 7.586164e-16, 
    7.598534e-16, 7.602991e-16, 7.615344e-16, 7.622781e-16, 7.630216e-16, 
    7.633464e-16, 7.634447e-16, 7.634852e-16 ;

 F_N2O_NIT =
  2.408731e-14, 2.429515e-14, 2.425467e-14, 2.442284e-14, 2.432947e-14, 
    2.44397e-14, 2.412936e-14, 2.430341e-14, 2.419222e-14, 2.410595e-14, 
    2.475091e-14, 2.443034e-14, 2.508615e-14, 2.488003e-14, 2.539948e-14, 
    2.505402e-14, 2.546943e-14, 2.538947e-14, 2.56305e-14, 2.556132e-14, 
    2.587092e-14, 2.566245e-14, 2.603216e-14, 2.582105e-14, 2.585401e-14, 
    2.565558e-14, 2.449469e-14, 2.47109e-14, 2.448191e-14, 2.451267e-14, 
    2.449886e-14, 2.433139e-14, 2.424723e-14, 2.407143e-14, 2.410329e-14, 
    2.423243e-14, 2.452649e-14, 2.442646e-14, 2.467895e-14, 2.467323e-14, 
    2.495588e-14, 2.482823e-14, 2.530578e-14, 2.516957e-14, 2.556421e-14, 
    2.546466e-14, 2.555952e-14, 2.553073e-14, 2.555989e-14, 2.541398e-14, 
    2.547644e-14, 2.534823e-14, 2.485214e-14, 2.499743e-14, 2.45654e-14, 
    2.43075e-14, 2.413697e-14, 2.401634e-14, 2.403337e-14, 2.406586e-14, 
    2.423318e-14, 2.439104e-14, 2.45117e-14, 2.459258e-14, 2.46724e-14, 
    2.491487e-14, 2.504369e-14, 2.533337e-14, 2.528095e-14, 2.536977e-14, 
    2.545476e-14, 2.559779e-14, 2.557422e-14, 2.563734e-14, 2.536741e-14, 
    2.554664e-14, 2.525111e-14, 2.533176e-14, 2.469418e-14, 2.445343e-14, 
    2.435149e-14, 2.426243e-14, 2.404647e-14, 2.41955e-14, 2.413669e-14, 
    2.42767e-14, 2.436589e-14, 2.432175e-14, 2.459479e-14, 2.448845e-14, 
    2.505133e-14, 2.480807e-14, 2.544484e-14, 2.52917e-14, 2.548161e-14, 
    2.538461e-14, 2.555093e-14, 2.540121e-14, 2.566084e-14, 2.571756e-14, 
    2.567879e-14, 2.582786e-14, 2.539291e-14, 2.55595e-14, 2.432053e-14, 
    2.432773e-14, 2.436126e-14, 2.421403e-14, 2.420504e-14, 2.407054e-14, 
    2.419019e-14, 2.424124e-14, 2.437106e-14, 2.444802e-14, 2.452129e-14, 
    2.468281e-14, 2.486383e-14, 2.511811e-14, 2.530161e-14, 2.5425e-14, 
    2.53493e-14, 2.541612e-14, 2.534142e-14, 2.530644e-14, 2.569629e-14, 
    2.547701e-14, 2.580639e-14, 2.57881e-14, 2.563882e-14, 2.579015e-14, 
    2.433278e-14, 2.429138e-14, 2.414795e-14, 2.426016e-14, 2.405592e-14, 
    2.417013e-14, 2.423593e-14, 2.449067e-14, 2.454682e-14, 2.459895e-14, 
    2.470207e-14, 2.483474e-14, 2.506836e-14, 2.527255e-14, 2.54597e-14, 
    2.544596e-14, 2.545079e-14, 2.549269e-14, 2.538897e-14, 2.550973e-14, 
    2.553003e-14, 2.547697e-14, 2.578565e-14, 2.569726e-14, 2.57877e-14, 
    2.573013e-14, 2.430483e-14, 2.437451e-14, 2.433684e-14, 2.44077e-14, 
    2.435777e-14, 2.458021e-14, 2.46471e-14, 2.496135e-14, 2.483212e-14, 
    2.503795e-14, 2.485298e-14, 2.488571e-14, 2.504468e-14, 2.486295e-14, 
    2.526127e-14, 2.499087e-14, 2.549432e-14, 2.522301e-14, 2.551136e-14, 
    2.545887e-14, 2.55458e-14, 2.562379e-14, 2.572208e-14, 2.590396e-14, 
    2.586178e-14, 2.601426e-14, 2.447859e-14, 2.456934e-14, 2.456133e-14, 
    2.465646e-14, 2.472694e-14, 2.488005e-14, 2.512664e-14, 2.503376e-14, 
    2.52044e-14, 2.523873e-14, 2.497953e-14, 2.513851e-14, 2.463014e-14, 
    2.471191e-14, 2.46632e-14, 2.448571e-14, 2.505513e-14, 2.476206e-14, 
    2.530462e-14, 2.514481e-14, 2.561266e-14, 2.537943e-14, 2.583857e-14, 
    2.603616e-14, 2.622282e-14, 2.644184e-14, 2.461893e-14, 2.455718e-14, 
    2.466778e-14, 2.482124e-14, 2.496405e-14, 2.515458e-14, 2.517411e-14, 
    2.520989e-14, 2.530272e-14, 2.538091e-14, 2.522121e-14, 2.540052e-14, 
    2.47309e-14, 2.508065e-14, 2.453383e-14, 2.469784e-14, 2.481214e-14, 
    2.476196e-14, 2.502312e-14, 2.508488e-14, 2.533666e-14, 2.520634e-14, 
    2.598732e-14, 2.564027e-14, 2.660922e-14, 2.633657e-14, 2.453563e-14, 
    2.46187e-14, 2.490898e-14, 2.477065e-14, 2.516731e-14, 2.526545e-14, 
    2.534537e-14, 2.544773e-14, 2.545879e-14, 2.551955e-14, 2.542001e-14, 
    2.551561e-14, 2.515495e-14, 2.531579e-14, 2.487568e-14, 2.498243e-14, 
    2.493329e-14, 2.487944e-14, 2.504581e-14, 2.52237e-14, 2.522749e-14, 
    2.528467e-14, 2.544618e-14, 2.516888e-14, 2.603229e-14, 2.54973e-14, 
    2.470946e-14, 2.48702e-14, 2.48932e-14, 2.483084e-14, 2.52556e-14, 
    2.510126e-14, 2.551807e-14, 2.540506e-14, 2.559035e-14, 2.549819e-14, 
    2.548464e-14, 2.536656e-14, 2.529318e-14, 2.510831e-14, 2.495839e-14, 
    2.483984e-14, 2.486738e-14, 2.499769e-14, 2.523459e-14, 2.545976e-14, 
    2.541035e-14, 2.557621e-14, 2.513839e-14, 2.53215e-14, 2.525064e-14, 
    2.54356e-14, 2.503129e-14, 2.537544e-14, 2.494371e-14, 2.49814e-14, 
    2.509819e-14, 2.533399e-14, 2.538629e-14, 2.544222e-14, 2.54077e-14, 
    2.524064e-14, 2.521331e-14, 2.509533e-14, 2.506281e-14, 2.497317e-14, 
    2.489907e-14, 2.496676e-14, 2.503795e-14, 2.524068e-14, 2.542411e-14, 
    2.562487e-14, 2.567413e-14, 2.590999e-14, 2.571791e-14, 2.603528e-14, 
    2.576534e-14, 2.623353e-14, 2.539544e-14, 2.575746e-14, 2.510351e-14, 
    2.517354e-14, 2.530047e-14, 2.559282e-14, 2.543476e-14, 2.561965e-14, 
    2.521224e-14, 2.50022e-14, 2.4948e-14, 2.484704e-14, 2.49503e-14, 
    2.494189e-14, 2.504089e-14, 2.500905e-14, 2.524742e-14, 2.511923e-14, 
    2.548427e-14, 2.561816e-14, 2.599823e-14, 2.623265e-14, 2.64724e-14, 
    2.65786e-14, 2.661096e-14, 2.66245e-14 ;

 F_NIT =
  4.014551e-11, 4.049193e-11, 4.042445e-11, 4.070474e-11, 4.054912e-11, 
    4.073283e-11, 4.021559e-11, 4.050569e-11, 4.032037e-11, 4.017659e-11, 
    4.125151e-11, 4.071723e-11, 4.181026e-11, 4.146671e-11, 4.233246e-11, 
    4.17567e-11, 4.244905e-11, 4.231578e-11, 4.27175e-11, 4.260221e-11, 
    4.31182e-11, 4.277076e-11, 4.338693e-11, 4.303508e-11, 4.309002e-11, 
    4.27593e-11, 4.082448e-11, 4.118483e-11, 4.080318e-11, 4.085445e-11, 
    4.083144e-11, 4.055232e-11, 4.041205e-11, 4.011905e-11, 4.017215e-11, 
    4.038738e-11, 4.087749e-11, 4.071076e-11, 4.113158e-11, 4.112206e-11, 
    4.159313e-11, 4.138039e-11, 4.21763e-11, 4.194928e-11, 4.260701e-11, 
    4.24411e-11, 4.25992e-11, 4.255122e-11, 4.259982e-11, 4.235663e-11, 
    4.246073e-11, 4.224705e-11, 4.142024e-11, 4.166238e-11, 4.094233e-11, 
    4.05125e-11, 4.022828e-11, 4.002723e-11, 4.005561e-11, 4.010976e-11, 
    4.038864e-11, 4.065173e-11, 4.085283e-11, 4.098763e-11, 4.112067e-11, 
    4.152479e-11, 4.173948e-11, 4.222228e-11, 4.213492e-11, 4.228295e-11, 
    4.24246e-11, 4.266299e-11, 4.26237e-11, 4.272889e-11, 4.227901e-11, 
    4.257773e-11, 4.208518e-11, 4.22196e-11, 4.115696e-11, 4.075572e-11, 
    4.058582e-11, 4.043738e-11, 4.007744e-11, 4.032583e-11, 4.022781e-11, 
    4.046117e-11, 4.060982e-11, 4.053626e-11, 4.099131e-11, 4.081408e-11, 
    4.175221e-11, 4.134678e-11, 4.240807e-11, 4.215283e-11, 4.246935e-11, 
    4.230769e-11, 4.258488e-11, 4.233536e-11, 4.276807e-11, 4.28626e-11, 
    4.279798e-11, 4.304643e-11, 4.232152e-11, 4.259916e-11, 4.053422e-11, 
    4.054622e-11, 4.06021e-11, 4.035672e-11, 4.034173e-11, 4.011757e-11, 
    4.031698e-11, 4.040206e-11, 4.061843e-11, 4.07467e-11, 4.086882e-11, 
    4.113801e-11, 4.143972e-11, 4.186351e-11, 4.216935e-11, 4.2375e-11, 
    4.224883e-11, 4.236021e-11, 4.22357e-11, 4.217741e-11, 4.282716e-11, 
    4.246168e-11, 4.301064e-11, 4.298017e-11, 4.273137e-11, 4.298359e-11, 
    4.055463e-11, 4.048563e-11, 4.024659e-11, 4.043359e-11, 4.009319e-11, 
    4.028355e-11, 4.039321e-11, 4.081778e-11, 4.091136e-11, 4.099825e-11, 
    4.117012e-11, 4.139123e-11, 4.178061e-11, 4.212092e-11, 4.243283e-11, 
    4.240993e-11, 4.241799e-11, 4.248782e-11, 4.231495e-11, 4.251622e-11, 
    4.255005e-11, 4.246162e-11, 4.297608e-11, 4.282877e-11, 4.297951e-11, 
    4.288355e-11, 4.050804e-11, 4.062419e-11, 4.05614e-11, 4.06795e-11, 
    4.059628e-11, 4.096701e-11, 4.10785e-11, 4.160226e-11, 4.138687e-11, 
    4.172991e-11, 4.142164e-11, 4.147618e-11, 4.174113e-11, 4.143826e-11, 
    4.210211e-11, 4.165145e-11, 4.249052e-11, 4.203836e-11, 4.251894e-11, 
    4.243145e-11, 4.257633e-11, 4.270632e-11, 4.287013e-11, 4.317326e-11, 
    4.310296e-11, 4.33571e-11, 4.079765e-11, 4.094889e-11, 4.093556e-11, 
    4.10941e-11, 4.121157e-11, 4.146675e-11, 4.187774e-11, 4.172293e-11, 
    4.200734e-11, 4.206455e-11, 4.163255e-11, 4.189752e-11, 4.105023e-11, 
    4.118651e-11, 4.110533e-11, 4.080952e-11, 4.175855e-11, 4.127009e-11, 
    4.217436e-11, 4.190802e-11, 4.268777e-11, 4.229906e-11, 4.306429e-11, 
    4.339361e-11, 4.370469e-11, 4.406973e-11, 4.103155e-11, 4.092864e-11, 
    4.111297e-11, 4.136873e-11, 4.160675e-11, 4.192429e-11, 4.195684e-11, 
    4.201649e-11, 4.217119e-11, 4.230151e-11, 4.203536e-11, 4.23342e-11, 
    4.121816e-11, 4.180109e-11, 4.088972e-11, 4.116307e-11, 4.135357e-11, 
    4.126994e-11, 4.170521e-11, 4.180813e-11, 4.222776e-11, 4.201057e-11, 
    4.33122e-11, 4.273379e-11, 4.434871e-11, 4.389429e-11, 4.089271e-11, 
    4.103117e-11, 4.151497e-11, 4.128441e-11, 4.194552e-11, 4.210908e-11, 
    4.224228e-11, 4.241289e-11, 4.243132e-11, 4.253259e-11, 4.236669e-11, 
    4.252602e-11, 4.192493e-11, 4.219299e-11, 4.145947e-11, 4.163739e-11, 
    4.155548e-11, 4.146574e-11, 4.174302e-11, 4.20395e-11, 4.204583e-11, 
    4.214112e-11, 4.24103e-11, 4.194813e-11, 4.338715e-11, 4.24955e-11, 
    4.118243e-11, 4.145034e-11, 4.148866e-11, 4.138473e-11, 4.209266e-11, 
    4.183543e-11, 4.253012e-11, 4.234177e-11, 4.265058e-11, 4.249698e-11, 
    4.24744e-11, 4.22776e-11, 4.215531e-11, 4.184718e-11, 4.159732e-11, 
    4.139974e-11, 4.144563e-11, 4.166282e-11, 4.205765e-11, 4.243294e-11, 
    4.235058e-11, 4.262701e-11, 4.189732e-11, 4.22025e-11, 4.208441e-11, 
    4.239267e-11, 4.171881e-11, 4.22924e-11, 4.157284e-11, 4.163567e-11, 
    4.183032e-11, 4.222332e-11, 4.231049e-11, 4.240371e-11, 4.234616e-11, 
    4.206773e-11, 4.202219e-11, 4.182556e-11, 4.177135e-11, 4.162195e-11, 
    4.149846e-11, 4.161127e-11, 4.172991e-11, 4.206781e-11, 4.237352e-11, 
    4.270813e-11, 4.279021e-11, 4.318331e-11, 4.286318e-11, 4.339213e-11, 
    4.294223e-11, 4.372255e-11, 4.232573e-11, 4.29291e-11, 4.183919e-11, 
    4.19559e-11, 4.216745e-11, 4.26547e-11, 4.239127e-11, 4.269943e-11, 
    4.20204e-11, 4.167033e-11, 4.157999e-11, 4.141174e-11, 4.158383e-11, 
    4.156982e-11, 4.173482e-11, 4.168175e-11, 4.207904e-11, 4.186539e-11, 
    4.247378e-11, 4.269693e-11, 4.333038e-11, 4.372109e-11, 4.412066e-11, 
    4.429766e-11, 4.435161e-11, 4.437416e-11 ;

 F_NIT_vr =
  2.347564e-10, 2.357934e-10, 2.355912e-10, 2.364283e-10, 2.359636e-10, 
    2.365114e-10, 2.349653e-10, 2.35833e-10, 2.352787e-10, 2.348476e-10, 
    2.380524e-10, 2.364637e-10, 2.397047e-10, 2.386894e-10, 2.412401e-10, 
    2.39546e-10, 2.415818e-10, 2.411906e-10, 2.423672e-10, 2.420296e-10, 
    2.435355e-10, 2.425222e-10, 2.443165e-10, 2.43293e-10, 2.434528e-10, 
    2.424876e-10, 2.367849e-10, 2.378563e-10, 2.36721e-10, 2.368738e-10, 
    2.368049e-10, 2.359722e-10, 2.355528e-10, 2.346749e-10, 2.348339e-10, 
    2.354785e-10, 2.369407e-10, 2.364436e-10, 2.376955e-10, 2.376673e-10, 
    2.390624e-10, 2.384329e-10, 2.407807e-10, 2.401126e-10, 2.420434e-10, 
    2.415571e-10, 2.420201e-10, 2.418792e-10, 2.420212e-10, 2.413087e-10, 
    2.416134e-10, 2.409866e-10, 2.385536e-10, 2.392694e-10, 2.371349e-10, 
    2.35853e-10, 2.350024e-10, 2.343994e-10, 2.344842e-10, 2.346467e-10, 
    2.354818e-10, 2.362674e-10, 2.368667e-10, 2.372675e-10, 2.376625e-10, 
    2.388601e-10, 2.394942e-10, 2.409153e-10, 2.406585e-10, 2.41093e-10, 
    2.415085e-10, 2.422062e-10, 2.420911e-10, 2.423984e-10, 2.410802e-10, 
    2.41956e-10, 2.405103e-10, 2.409054e-10, 2.377725e-10, 2.365787e-10, 
    2.360717e-10, 2.356279e-10, 2.345495e-10, 2.35294e-10, 2.350001e-10, 
    2.356982e-10, 2.361421e-10, 2.359221e-10, 2.372782e-10, 2.367503e-10, 
    2.395314e-10, 2.383326e-10, 2.414603e-10, 2.407106e-10, 2.416393e-10, 
    2.411652e-10, 2.419772e-10, 2.41246e-10, 2.425124e-10, 2.427885e-10, 
    2.425994e-10, 2.433242e-10, 2.412039e-10, 2.420177e-10, 2.359173e-10, 
    2.359532e-10, 2.361198e-10, 2.35386e-10, 2.353411e-10, 2.346691e-10, 
    2.352664e-10, 2.35521e-10, 2.361672e-10, 2.365494e-10, 2.369129e-10, 
    2.377133e-10, 2.386074e-10, 2.398589e-10, 2.407589e-10, 2.413624e-10, 
    2.40992e-10, 2.413185e-10, 2.40953e-10, 2.407813e-10, 2.426844e-10, 
    2.416153e-10, 2.432193e-10, 2.431305e-10, 2.424038e-10, 2.431398e-10, 
    2.359779e-10, 2.357714e-10, 2.350561e-10, 2.356154e-10, 2.345956e-10, 
    2.351662e-10, 2.354941e-10, 2.36761e-10, 2.370394e-10, 2.372978e-10, 
    2.378081e-10, 2.384633e-10, 2.396142e-10, 2.40616e-10, 2.415317e-10, 
    2.414642e-10, 2.414877e-10, 2.41692e-10, 2.41185e-10, 2.417747e-10, 
    2.418735e-10, 2.416145e-10, 2.431179e-10, 2.426881e-10, 2.431276e-10, 
    2.428474e-10, 2.358381e-10, 2.361846e-10, 2.359969e-10, 2.363494e-10, 
    2.361005e-10, 2.372052e-10, 2.375363e-10, 2.390879e-10, 2.384504e-10, 
    2.394647e-10, 2.385529e-10, 2.387144e-10, 2.39497e-10, 2.386015e-10, 
    2.4056e-10, 2.392314e-10, 2.416997e-10, 2.403717e-10, 2.417825e-10, 
    2.415257e-10, 2.419498e-10, 2.423302e-10, 2.428082e-10, 2.436917e-10, 
    2.434865e-10, 2.442258e-10, 2.367016e-10, 2.371514e-10, 2.371117e-10, 
    2.375826e-10, 2.37931e-10, 2.386872e-10, 2.399007e-10, 2.394438e-10, 
    2.402818e-10, 2.404502e-10, 2.391761e-10, 2.39958e-10, 2.374504e-10, 
    2.378547e-10, 2.376137e-10, 2.367334e-10, 2.39547e-10, 2.381018e-10, 
    2.407709e-10, 2.399869e-10, 2.422752e-10, 2.411365e-10, 2.433737e-10, 
    2.443316e-10, 2.452334e-10, 2.46288e-10, 2.37397e-10, 2.370906e-10, 
    2.376382e-10, 2.383969e-10, 2.391006e-10, 2.400376e-10, 2.401332e-10, 
    2.403084e-10, 2.40763e-10, 2.411458e-10, 2.403634e-10, 2.412411e-10, 
    2.379484e-10, 2.396724e-10, 2.369717e-10, 2.377843e-10, 2.383488e-10, 
    2.381009e-10, 2.393885e-10, 2.396918e-10, 2.409265e-10, 2.40288e-10, 
    2.440944e-10, 2.424087e-10, 2.470914e-10, 2.45781e-10, 2.369834e-10, 
    2.373949e-10, 2.388291e-10, 2.381464e-10, 2.400995e-10, 2.405808e-10, 
    2.409717e-10, 2.414724e-10, 2.415259e-10, 2.418227e-10, 2.41336e-10, 
    2.41803e-10, 2.40037e-10, 2.408256e-10, 2.386624e-10, 2.391881e-10, 
    2.389459e-10, 2.386801e-10, 2.394993e-10, 2.40373e-10, 2.403913e-10, 
    2.406711e-10, 2.414612e-10, 2.401029e-10, 2.443113e-10, 2.417101e-10, 
    2.378439e-10, 2.386375e-10, 2.387506e-10, 2.38443e-10, 2.40532e-10, 
    2.397745e-10, 2.418155e-10, 2.41263e-10, 2.421674e-10, 2.417178e-10, 
    2.416511e-10, 2.41074e-10, 2.407142e-10, 2.398073e-10, 2.390692e-10, 
    2.384848e-10, 2.386202e-10, 2.392624e-10, 2.404258e-10, 2.415278e-10, 
    2.41286e-10, 2.420956e-10, 2.399528e-10, 2.408507e-10, 2.405031e-10, 
    2.414084e-10, 2.394306e-10, 2.41119e-10, 2.389992e-10, 2.391845e-10, 
    2.397587e-10, 2.409153e-10, 2.411708e-10, 2.414443e-10, 2.41275e-10, 
    2.404571e-10, 2.403228e-10, 2.397432e-10, 2.39583e-10, 2.391419e-10, 
    2.387763e-10, 2.391099e-10, 2.394598e-10, 2.404556e-10, 2.413531e-10, 
    2.423326e-10, 2.425724e-10, 2.43718e-10, 2.427849e-10, 2.443246e-10, 
    2.43015e-10, 2.452822e-10, 2.412162e-10, 2.429815e-10, 2.397849e-10, 
    2.401285e-10, 2.407506e-10, 2.421789e-10, 2.414071e-10, 2.423095e-10, 
    2.403174e-10, 2.392849e-10, 2.390177e-10, 2.3852e-10, 2.390286e-10, 
    2.389873e-10, 2.394744e-10, 2.393173e-10, 2.404879e-10, 2.398589e-10, 
    2.416463e-10, 2.422995e-10, 2.441455e-10, 2.452783e-10, 2.464327e-10, 
    2.469423e-10, 2.470975e-10, 2.471621e-10,
  1.335097e-10, 1.345181e-10, 1.343218e-10, 1.351368e-10, 1.346845e-10, 
    1.352185e-10, 1.337139e-10, 1.345582e-10, 1.34019e-10, 1.336004e-10, 
    1.367235e-10, 1.351732e-10, 1.383408e-10, 1.37347e-10, 1.398483e-10, 
    1.381859e-10, 1.401844e-10, 1.398003e-10, 1.409575e-10, 1.406256e-10, 
    1.421095e-10, 1.411108e-10, 1.428809e-10, 1.418708e-10, 1.420286e-10, 
    1.410779e-10, 1.354847e-10, 1.365301e-10, 1.354229e-10, 1.355717e-10, 
    1.355049e-10, 1.346938e-10, 1.342858e-10, 1.334327e-10, 1.335874e-10, 
    1.342141e-10, 1.356387e-10, 1.351545e-10, 1.363761e-10, 1.363484e-10, 
    1.37713e-10, 1.370971e-10, 1.39398e-10, 1.387427e-10, 1.406395e-10, 
    1.401616e-10, 1.40617e-10, 1.404789e-10, 1.406188e-10, 1.399181e-10, 
    1.402182e-10, 1.396022e-10, 1.372124e-10, 1.379132e-10, 1.358269e-10, 
    1.34578e-10, 1.337509e-10, 1.331651e-10, 1.332479e-10, 1.334057e-10, 
    1.342177e-10, 1.34983e-10, 1.355672e-10, 1.359585e-10, 1.363445e-10, 
    1.375151e-10, 1.381362e-10, 1.395306e-10, 1.392786e-10, 1.397056e-10, 
    1.40114e-10, 1.408007e-10, 1.406876e-10, 1.409904e-10, 1.396944e-10, 
    1.405552e-10, 1.391352e-10, 1.39523e-10, 1.364493e-10, 1.352851e-10, 
    1.347912e-10, 1.343596e-10, 1.333115e-10, 1.340349e-10, 1.337496e-10, 
    1.344289e-10, 1.348611e-10, 1.346473e-10, 1.359692e-10, 1.354547e-10, 
    1.381731e-10, 1.369998e-10, 1.400664e-10, 1.393303e-10, 1.40243e-10, 
    1.39777e-10, 1.405758e-10, 1.398568e-10, 1.411031e-10, 1.41375e-10, 
    1.411892e-10, 1.419035e-10, 1.39817e-10, 1.40617e-10, 1.346413e-10, 
    1.346762e-10, 1.348387e-10, 1.341249e-10, 1.340813e-10, 1.334285e-10, 
    1.340093e-10, 1.342569e-10, 1.348862e-10, 1.35259e-10, 1.356137e-10, 
    1.363947e-10, 1.37269e-10, 1.384949e-10, 1.39378e-10, 1.399711e-10, 
    1.396073e-10, 1.399285e-10, 1.395695e-10, 1.394013e-10, 1.412731e-10, 
    1.40221e-10, 1.418007e-10, 1.417131e-10, 1.409976e-10, 1.41723e-10, 
    1.347007e-10, 1.345e-10, 1.338043e-10, 1.343486e-10, 1.333575e-10, 
    1.339119e-10, 1.342311e-10, 1.354654e-10, 1.357372e-10, 1.359893e-10, 
    1.364879e-10, 1.371286e-10, 1.382553e-10, 1.392382e-10, 1.401378e-10, 
    1.400719e-10, 1.400951e-10, 1.402963e-10, 1.39798e-10, 1.403782e-10, 
    1.404756e-10, 1.402209e-10, 1.417014e-10, 1.412779e-10, 1.417113e-10, 
    1.414354e-10, 1.345652e-10, 1.349029e-10, 1.347204e-10, 1.350637e-10, 
    1.348218e-10, 1.358986e-10, 1.362221e-10, 1.377394e-10, 1.37116e-10, 
    1.381087e-10, 1.372167e-10, 1.373746e-10, 1.381411e-10, 1.372649e-10, 
    1.39184e-10, 1.378818e-10, 1.403041e-10, 1.389999e-10, 1.40386e-10, 
    1.401339e-10, 1.405513e-10, 1.409255e-10, 1.413968e-10, 1.422679e-10, 
    1.42066e-10, 1.427956e-10, 1.35407e-10, 1.358461e-10, 1.358074e-10, 
    1.362674e-10, 1.36608e-10, 1.373473e-10, 1.38536e-10, 1.380886e-10, 
    1.389104e-10, 1.390756e-10, 1.378272e-10, 1.385932e-10, 1.361402e-10, 
    1.365354e-10, 1.363001e-10, 1.354416e-10, 1.381916e-10, 1.367778e-10, 
    1.393926e-10, 1.386237e-10, 1.408722e-10, 1.397523e-10, 1.419549e-10, 
    1.429002e-10, 1.43792e-10, 1.448365e-10, 1.360859e-10, 1.357874e-10, 
    1.363222e-10, 1.370634e-10, 1.377525e-10, 1.386705e-10, 1.387646e-10, 
    1.389368e-10, 1.393834e-10, 1.397593e-10, 1.389913e-10, 1.398536e-10, 
    1.366271e-10, 1.383146e-10, 1.356745e-10, 1.364675e-10, 1.370197e-10, 
    1.367774e-10, 1.380375e-10, 1.383351e-10, 1.395467e-10, 1.389199e-10, 
    1.426667e-10, 1.410046e-10, 1.456336e-10, 1.443347e-10, 1.356831e-10, 
    1.360849e-10, 1.374869e-10, 1.368192e-10, 1.387319e-10, 1.392041e-10, 
    1.395885e-10, 1.400804e-10, 1.401335e-10, 1.404253e-10, 1.399473e-10, 
    1.404064e-10, 1.386725e-10, 1.394464e-10, 1.373264e-10, 1.378413e-10, 
    1.376043e-10, 1.373446e-10, 1.381469e-10, 1.390034e-10, 1.390217e-10, 
    1.392968e-10, 1.400729e-10, 1.387397e-10, 1.428816e-10, 1.403184e-10, 
    1.365236e-10, 1.372998e-10, 1.374108e-10, 1.371099e-10, 1.391568e-10, 
    1.384138e-10, 1.404182e-10, 1.398754e-10, 1.407651e-10, 1.403228e-10, 
    1.402577e-10, 1.396904e-10, 1.393377e-10, 1.384479e-10, 1.377254e-10, 
    1.371535e-10, 1.372864e-10, 1.379149e-10, 1.390559e-10, 1.401383e-10, 
    1.399009e-10, 1.406974e-10, 1.385929e-10, 1.394739e-10, 1.391332e-10, 
    1.400224e-10, 1.380767e-10, 1.397328e-10, 1.376545e-10, 1.378363e-10, 
    1.383991e-10, 1.395337e-10, 1.397853e-10, 1.40054e-10, 1.398881e-10, 
    1.390849e-10, 1.389534e-10, 1.383854e-10, 1.382287e-10, 1.377967e-10, 
    1.374393e-10, 1.377658e-10, 1.38109e-10, 1.390852e-10, 1.399671e-10, 
    1.409309e-10, 1.411671e-10, 1.422968e-10, 1.413769e-10, 1.428959e-10, 
    1.41604e-10, 1.438431e-10, 1.39829e-10, 1.415662e-10, 1.384247e-10, 
    1.38762e-10, 1.393726e-10, 1.407769e-10, 1.400182e-10, 1.409057e-10, 
    1.389483e-10, 1.379366e-10, 1.376753e-10, 1.371882e-10, 1.376864e-10, 
    1.376459e-10, 1.381232e-10, 1.379697e-10, 1.391177e-10, 1.385006e-10, 
    1.402561e-10, 1.408987e-10, 1.42719e-10, 1.43839e-10, 1.449823e-10, 
    1.45488e-10, 1.456421e-10, 1.457065e-10,
  1.248478e-10, 1.259514e-10, 1.257365e-10, 1.26629e-10, 1.261336e-10, 
    1.267185e-10, 1.250712e-10, 1.259953e-10, 1.25405e-10, 1.24947e-10, 
    1.283686e-10, 1.266689e-10, 1.301443e-10, 1.290529e-10, 1.31802e-10, 
    1.299742e-10, 1.321718e-10, 1.317491e-10, 1.330231e-10, 1.326576e-10, 
    1.342925e-10, 1.331919e-10, 1.351434e-10, 1.340294e-10, 1.342034e-10, 
    1.331557e-10, 1.270102e-10, 1.281564e-10, 1.269424e-10, 1.271056e-10, 
    1.270324e-10, 1.261438e-10, 1.25697e-10, 1.247636e-10, 1.249329e-10, 
    1.256186e-10, 1.27179e-10, 1.266484e-10, 1.279875e-10, 1.279572e-10, 
    1.294547e-10, 1.287786e-10, 1.313066e-10, 1.30586e-10, 1.326728e-10, 
    1.321467e-10, 1.326481e-10, 1.32496e-10, 1.326501e-10, 1.318788e-10, 
    1.32209e-10, 1.315312e-10, 1.289051e-10, 1.296746e-10, 1.273853e-10, 
    1.260169e-10, 1.251117e-10, 1.244709e-10, 1.245614e-10, 1.24734e-10, 
    1.256226e-10, 1.264605e-10, 1.271006e-10, 1.275296e-10, 1.279528e-10, 
    1.292374e-10, 1.299196e-10, 1.314525e-10, 1.311753e-10, 1.31645e-10, 
    1.320944e-10, 1.328503e-10, 1.327258e-10, 1.330593e-10, 1.316326e-10, 
    1.325801e-10, 1.310176e-10, 1.314441e-10, 1.280678e-10, 1.267915e-10, 
    1.262505e-10, 1.257778e-10, 1.24631e-10, 1.254225e-10, 1.251102e-10, 
    1.258537e-10, 1.26327e-10, 1.260928e-10, 1.275413e-10, 1.269773e-10, 
    1.299601e-10, 1.286718e-10, 1.32042e-10, 1.312322e-10, 1.322364e-10, 
    1.317236e-10, 1.326027e-10, 1.318114e-10, 1.331835e-10, 1.33483e-10, 
    1.332783e-10, 1.340655e-10, 1.317676e-10, 1.326481e-10, 1.260863e-10, 
    1.261245e-10, 1.263024e-10, 1.255209e-10, 1.254732e-10, 1.24759e-10, 
    1.253944e-10, 1.256654e-10, 1.263545e-10, 1.267629e-10, 1.271516e-10, 
    1.28008e-10, 1.289672e-10, 1.303137e-10, 1.312846e-10, 1.319371e-10, 
    1.315369e-10, 1.318902e-10, 1.314952e-10, 1.313103e-10, 1.333707e-10, 
    1.322121e-10, 1.339521e-10, 1.338556e-10, 1.330672e-10, 1.338665e-10, 
    1.261513e-10, 1.259316e-10, 1.251701e-10, 1.257659e-10, 1.246813e-10, 
    1.252879e-10, 1.256372e-10, 1.269891e-10, 1.27287e-10, 1.275634e-10, 
    1.281101e-10, 1.288132e-10, 1.300504e-10, 1.311309e-10, 1.321206e-10, 
    1.32048e-10, 1.320735e-10, 1.32295e-10, 1.317467e-10, 1.323851e-10, 
    1.324924e-10, 1.32212e-10, 1.338427e-10, 1.33376e-10, 1.338536e-10, 
    1.335496e-10, 1.26003e-10, 1.263728e-10, 1.261729e-10, 1.265489e-10, 
    1.26284e-10, 1.274639e-10, 1.278186e-10, 1.294837e-10, 1.287993e-10, 
    1.298893e-10, 1.289099e-10, 1.290832e-10, 1.299249e-10, 1.289627e-10, 
    1.310712e-10, 1.296401e-10, 1.323036e-10, 1.308688e-10, 1.323937e-10, 
    1.321163e-10, 1.325758e-10, 1.329879e-10, 1.335071e-10, 1.344672e-10, 
    1.342446e-10, 1.350492e-10, 1.26925e-10, 1.274063e-10, 1.273639e-10, 
    1.278683e-10, 1.282419e-10, 1.290532e-10, 1.303589e-10, 1.298672e-10, 
    1.307704e-10, 1.30952e-10, 1.295802e-10, 1.304217e-10, 1.277288e-10, 
    1.281623e-10, 1.279042e-10, 1.26963e-10, 1.299804e-10, 1.284281e-10, 
    1.313007e-10, 1.304552e-10, 1.329291e-10, 1.316963e-10, 1.341222e-10, 
    1.351647e-10, 1.361491e-10, 1.37303e-10, 1.276693e-10, 1.273419e-10, 
    1.279284e-10, 1.287416e-10, 1.294981e-10, 1.305067e-10, 1.306101e-10, 
    1.307995e-10, 1.312906e-10, 1.31704e-10, 1.308594e-10, 1.318078e-10, 
    1.282629e-10, 1.301156e-10, 1.272182e-10, 1.280878e-10, 1.286936e-10, 
    1.284277e-10, 1.298111e-10, 1.301381e-10, 1.314702e-10, 1.307809e-10, 
    1.349071e-10, 1.330749e-10, 1.381844e-10, 1.367485e-10, 1.272276e-10, 
    1.276682e-10, 1.292065e-10, 1.284736e-10, 1.305742e-10, 1.310934e-10, 
    1.315161e-10, 1.320574e-10, 1.321158e-10, 1.32437e-10, 1.319109e-10, 
    1.324162e-10, 1.305089e-10, 1.313598e-10, 1.290303e-10, 1.295956e-10, 
    1.293354e-10, 1.290502e-10, 1.299313e-10, 1.308726e-10, 1.308928e-10, 
    1.311953e-10, 1.320491e-10, 1.305827e-10, 1.351442e-10, 1.323194e-10, 
    1.281493e-10, 1.29001e-10, 1.291229e-10, 1.287926e-10, 1.310413e-10, 
    1.302246e-10, 1.324292e-10, 1.318319e-10, 1.328112e-10, 1.323241e-10, 
    1.322526e-10, 1.316283e-10, 1.312402e-10, 1.30262e-10, 1.294684e-10, 
    1.288405e-10, 1.289863e-10, 1.296765e-10, 1.309303e-10, 1.321211e-10, 
    1.318599e-10, 1.327366e-10, 1.304214e-10, 1.313901e-10, 1.310153e-10, 
    1.319935e-10, 1.298542e-10, 1.316749e-10, 1.293905e-10, 1.295901e-10, 
    1.302084e-10, 1.314559e-10, 1.317326e-10, 1.320283e-10, 1.318458e-10, 
    1.309622e-10, 1.308177e-10, 1.301934e-10, 1.300212e-10, 1.295466e-10, 
    1.291543e-10, 1.295127e-10, 1.298896e-10, 1.309626e-10, 1.319327e-10, 
    1.329937e-10, 1.332539e-10, 1.344991e-10, 1.334851e-10, 1.3516e-10, 
    1.337354e-10, 1.362055e-10, 1.317808e-10, 1.336937e-10, 1.302366e-10, 
    1.306072e-10, 1.312787e-10, 1.328242e-10, 1.319889e-10, 1.32966e-10, 
    1.308121e-10, 1.297003e-10, 1.294133e-10, 1.288786e-10, 1.294256e-10, 
    1.29381e-10, 1.299053e-10, 1.297367e-10, 1.309983e-10, 1.3032e-10, 
    1.322507e-10, 1.329583e-10, 1.349648e-10, 1.36201e-10, 1.374642e-10, 
    1.380233e-10, 1.381937e-10, 1.38265e-10,
  1.280645e-10, 1.292799e-10, 1.290432e-10, 1.300266e-10, 1.294806e-10, 
    1.301252e-10, 1.283104e-10, 1.293282e-10, 1.286781e-10, 1.281737e-10, 
    1.319453e-10, 1.300705e-10, 1.339062e-10, 1.327006e-10, 1.35739e-10, 
    1.337183e-10, 1.361483e-10, 1.356805e-10, 1.370906e-10, 1.366859e-10, 
    1.384971e-10, 1.372776e-10, 1.394404e-10, 1.382054e-10, 1.383982e-10, 
    1.372374e-10, 1.304468e-10, 1.317112e-10, 1.30372e-10, 1.305519e-10, 
    1.304712e-10, 1.294919e-10, 1.289997e-10, 1.279718e-10, 1.281581e-10, 
    1.289132e-10, 1.306329e-10, 1.300479e-10, 1.315246e-10, 1.314911e-10, 
    1.331443e-10, 1.323977e-10, 1.35191e-10, 1.343943e-10, 1.367028e-10, 
    1.361205e-10, 1.366754e-10, 1.36507e-10, 1.366776e-10, 1.35824e-10, 
    1.361894e-10, 1.354395e-10, 1.325374e-10, 1.333872e-10, 1.308604e-10, 
    1.293522e-10, 1.28355e-10, 1.276497e-10, 1.277493e-10, 1.279393e-10, 
    1.289177e-10, 1.298408e-10, 1.305464e-10, 1.310194e-10, 1.314863e-10, 
    1.329044e-10, 1.336579e-10, 1.353524e-10, 1.350458e-10, 1.355654e-10, 
    1.360626e-10, 1.368993e-10, 1.367614e-10, 1.371307e-10, 1.355517e-10, 
    1.366001e-10, 1.348714e-10, 1.353432e-10, 1.316134e-10, 1.302056e-10, 
    1.296094e-10, 1.290886e-10, 1.278259e-10, 1.286973e-10, 1.283534e-10, 
    1.291722e-10, 1.296937e-10, 1.294357e-10, 1.310324e-10, 1.304105e-10, 
    1.337026e-10, 1.322798e-10, 1.360046e-10, 1.351087e-10, 1.362197e-10, 
    1.356523e-10, 1.366252e-10, 1.357494e-10, 1.372682e-10, 1.376e-10, 
    1.373733e-10, 1.382454e-10, 1.357009e-10, 1.366754e-10, 1.294284e-10, 
    1.294705e-10, 1.296666e-10, 1.288057e-10, 1.287531e-10, 1.279667e-10, 
    1.286663e-10, 1.289648e-10, 1.29724e-10, 1.301741e-10, 1.306026e-10, 
    1.315472e-10, 1.32606e-10, 1.340933e-10, 1.351667e-10, 1.358886e-10, 
    1.354457e-10, 1.358366e-10, 1.353997e-10, 1.351951e-10, 1.374757e-10, 
    1.361928e-10, 1.381198e-10, 1.380128e-10, 1.371395e-10, 1.380248e-10, 
    1.295001e-10, 1.29258e-10, 1.284193e-10, 1.290754e-10, 1.278812e-10, 
    1.28549e-10, 1.289338e-10, 1.304235e-10, 1.307519e-10, 1.310568e-10, 
    1.316599e-10, 1.324359e-10, 1.338023e-10, 1.349968e-10, 1.360915e-10, 
    1.360112e-10, 1.360395e-10, 1.362846e-10, 1.356778e-10, 1.363843e-10, 
    1.365031e-10, 1.361927e-10, 1.379985e-10, 1.374814e-10, 1.380105e-10, 
    1.376737e-10, 1.293367e-10, 1.297442e-10, 1.295239e-10, 1.299383e-10, 
    1.296463e-10, 1.309471e-10, 1.313384e-10, 1.331764e-10, 1.324206e-10, 
    1.336244e-10, 1.325426e-10, 1.32734e-10, 1.336638e-10, 1.32601e-10, 
    1.349308e-10, 1.333491e-10, 1.362941e-10, 1.347071e-10, 1.363939e-10, 
    1.360868e-10, 1.365954e-10, 1.370516e-10, 1.376266e-10, 1.386907e-10, 
    1.384439e-10, 1.39336e-10, 1.303529e-10, 1.308836e-10, 1.308368e-10, 
    1.313931e-10, 1.318053e-10, 1.327009e-10, 1.341432e-10, 1.336e-10, 
    1.345981e-10, 1.347989e-10, 1.332828e-10, 1.342127e-10, 1.312393e-10, 
    1.317175e-10, 1.314327e-10, 1.303947e-10, 1.337251e-10, 1.320109e-10, 
    1.351845e-10, 1.342497e-10, 1.369865e-10, 1.356222e-10, 1.383082e-10, 
    1.394641e-10, 1.405562e-10, 1.418376e-10, 1.311736e-10, 1.308125e-10, 
    1.314594e-10, 1.323569e-10, 1.331922e-10, 1.343066e-10, 1.344209e-10, 
    1.346303e-10, 1.351733e-10, 1.356306e-10, 1.346965e-10, 1.357454e-10, 
    1.318286e-10, 1.338744e-10, 1.306761e-10, 1.316353e-10, 1.323039e-10, 
    1.320104e-10, 1.335379e-10, 1.338992e-10, 1.35372e-10, 1.346097e-10, 
    1.391784e-10, 1.371481e-10, 1.428169e-10, 1.412217e-10, 1.306865e-10, 
    1.311724e-10, 1.328701e-10, 1.32061e-10, 1.343812e-10, 1.349553e-10, 
    1.354228e-10, 1.360216e-10, 1.360863e-10, 1.364418e-10, 1.358595e-10, 
    1.364187e-10, 1.34309e-10, 1.352499e-10, 1.326755e-10, 1.332999e-10, 
    1.330125e-10, 1.326976e-10, 1.336707e-10, 1.347112e-10, 1.347334e-10, 
    1.350679e-10, 1.360127e-10, 1.343906e-10, 1.394415e-10, 1.363118e-10, 
    1.317032e-10, 1.326433e-10, 1.327778e-10, 1.324131e-10, 1.348977e-10, 
    1.339949e-10, 1.364331e-10, 1.35772e-10, 1.368559e-10, 1.363168e-10, 
    1.362376e-10, 1.355468e-10, 1.351177e-10, 1.340362e-10, 1.331593e-10, 
    1.32466e-10, 1.32627e-10, 1.333892e-10, 1.34775e-10, 1.360922e-10, 
    1.358031e-10, 1.367734e-10, 1.342123e-10, 1.352834e-10, 1.34869e-10, 
    1.359509e-10, 1.335855e-10, 1.355986e-10, 1.330733e-10, 1.332938e-10, 
    1.33977e-10, 1.353562e-10, 1.356623e-10, 1.359894e-10, 1.357875e-10, 
    1.348102e-10, 1.346504e-10, 1.339603e-10, 1.337701e-10, 1.332458e-10, 
    1.328124e-10, 1.332083e-10, 1.336247e-10, 1.348106e-10, 1.358836e-10, 
    1.370581e-10, 1.373463e-10, 1.387261e-10, 1.376024e-10, 1.394591e-10, 
    1.378798e-10, 1.40619e-10, 1.357157e-10, 1.378335e-10, 1.340081e-10, 
    1.344177e-10, 1.351602e-10, 1.368704e-10, 1.359458e-10, 1.370274e-10, 
    1.346442e-10, 1.334156e-10, 1.330986e-10, 1.325081e-10, 1.331121e-10, 
    1.330629e-10, 1.33642e-10, 1.334558e-10, 1.348501e-10, 1.341003e-10, 
    1.362356e-10, 1.370189e-10, 1.392424e-10, 1.406139e-10, 1.420165e-10, 
    1.426379e-10, 1.428273e-10, 1.429065e-10,
  1.381445e-10, 1.394321e-10, 1.391812e-10, 1.402237e-10, 1.396448e-10, 
    1.403282e-10, 1.38405e-10, 1.394834e-10, 1.387944e-10, 1.382601e-10, 
    1.422596e-10, 1.402703e-10, 1.443425e-10, 1.430614e-10, 1.462921e-10, 
    1.441428e-10, 1.467276e-10, 1.462297e-10, 1.477311e-10, 1.473001e-10, 
    1.492303e-10, 1.479303e-10, 1.502365e-10, 1.489192e-10, 1.491249e-10, 
    1.478875e-10, 1.406692e-10, 1.42011e-10, 1.4059e-10, 1.407808e-10, 
    1.406951e-10, 1.396568e-10, 1.391352e-10, 1.380463e-10, 1.382436e-10, 
    1.390436e-10, 1.408667e-10, 1.402462e-10, 1.418127e-10, 1.417772e-10, 
    1.435327e-10, 1.427397e-10, 1.457088e-10, 1.448613e-10, 1.47318e-10, 
    1.46698e-10, 1.472889e-10, 1.471096e-10, 1.472912e-10, 1.463824e-10, 
    1.467714e-10, 1.459732e-10, 1.42888e-10, 1.437908e-10, 1.411079e-10, 
    1.395088e-10, 1.384522e-10, 1.377052e-10, 1.378107e-10, 1.380119e-10, 
    1.390482e-10, 1.400266e-10, 1.407749e-10, 1.412767e-10, 1.417721e-10, 
    1.432781e-10, 1.440786e-10, 1.458806e-10, 1.455543e-10, 1.461072e-10, 
    1.466364e-10, 1.475274e-10, 1.473805e-10, 1.477738e-10, 1.460925e-10, 
    1.472087e-10, 1.453687e-10, 1.458707e-10, 1.419073e-10, 1.404134e-10, 
    1.397815e-10, 1.392294e-10, 1.378918e-10, 1.388148e-10, 1.384505e-10, 
    1.393179e-10, 1.398708e-10, 1.395972e-10, 1.412904e-10, 1.406308e-10, 
    1.441261e-10, 1.426145e-10, 1.465746e-10, 1.456213e-10, 1.468036e-10, 
    1.461996e-10, 1.472355e-10, 1.46303e-10, 1.479204e-10, 1.48274e-10, 
    1.480323e-10, 1.489618e-10, 1.462514e-10, 1.472889e-10, 1.395895e-10, 
    1.396341e-10, 1.39842e-10, 1.389296e-10, 1.388739e-10, 1.380409e-10, 
    1.387819e-10, 1.390982e-10, 1.399028e-10, 1.4038e-10, 1.408345e-10, 
    1.418368e-10, 1.429609e-10, 1.445414e-10, 1.45683e-10, 1.464511e-10, 
    1.459798e-10, 1.463958e-10, 1.459308e-10, 1.457131e-10, 1.481414e-10, 
    1.467751e-10, 1.488279e-10, 1.487138e-10, 1.477832e-10, 1.487267e-10, 
    1.396654e-10, 1.394089e-10, 1.385203e-10, 1.392154e-10, 1.379504e-10, 
    1.386577e-10, 1.390654e-10, 1.406446e-10, 1.409929e-10, 1.413163e-10, 
    1.419564e-10, 1.427802e-10, 1.442321e-10, 1.455022e-10, 1.466672e-10, 
    1.465816e-10, 1.466117e-10, 1.468727e-10, 1.462268e-10, 1.469789e-10, 
    1.471054e-10, 1.467749e-10, 1.486986e-10, 1.481475e-10, 1.487114e-10, 
    1.483525e-10, 1.394922e-10, 1.399242e-10, 1.396907e-10, 1.4013e-10, 
    1.398205e-10, 1.412001e-10, 1.416152e-10, 1.435669e-10, 1.42764e-10, 
    1.44043e-10, 1.428936e-10, 1.430969e-10, 1.44085e-10, 1.429556e-10, 
    1.454321e-10, 1.437505e-10, 1.468829e-10, 1.451941e-10, 1.469891e-10, 
    1.466621e-10, 1.472036e-10, 1.476896e-10, 1.483023e-10, 1.494367e-10, 
    1.491735e-10, 1.50125e-10, 1.405696e-10, 1.411326e-10, 1.410829e-10, 
    1.416733e-10, 1.421108e-10, 1.430617e-10, 1.445945e-10, 1.440169e-10, 
    1.450781e-10, 1.452917e-10, 1.436799e-10, 1.446684e-10, 1.4151e-10, 
    1.420176e-10, 1.417152e-10, 1.40614e-10, 1.4415e-10, 1.423291e-10, 
    1.457019e-10, 1.447076e-10, 1.476203e-10, 1.461676e-10, 1.490288e-10, 
    1.502619e-10, 1.514275e-10, 1.527967e-10, 1.414403e-10, 1.410572e-10, 
    1.417435e-10, 1.426964e-10, 1.435837e-10, 1.447682e-10, 1.448897e-10, 
    1.451123e-10, 1.456899e-10, 1.461766e-10, 1.451828e-10, 1.462988e-10, 
    1.421357e-10, 1.443086e-10, 1.409125e-10, 1.419304e-10, 1.426401e-10, 
    1.423285e-10, 1.43951e-10, 1.44335e-10, 1.459014e-10, 1.450904e-10, 
    1.49957e-10, 1.477925e-10, 1.538438e-10, 1.521385e-10, 1.409235e-10, 
    1.414389e-10, 1.432415e-10, 1.423822e-10, 1.448474e-10, 1.45458e-10, 
    1.459554e-10, 1.465927e-10, 1.466616e-10, 1.470401e-10, 1.464202e-10, 
    1.470155e-10, 1.447707e-10, 1.457714e-10, 1.430348e-10, 1.436981e-10, 
    1.433927e-10, 1.430582e-10, 1.440921e-10, 1.451985e-10, 1.452221e-10, 
    1.455779e-10, 1.465835e-10, 1.448575e-10, 1.50238e-10, 1.469019e-10, 
    1.420023e-10, 1.430007e-10, 1.431435e-10, 1.42756e-10, 1.453967e-10, 
    1.444367e-10, 1.470308e-10, 1.463271e-10, 1.474812e-10, 1.46907e-10, 
    1.468227e-10, 1.460874e-10, 1.456308e-10, 1.444807e-10, 1.435488e-10, 
    1.428122e-10, 1.429833e-10, 1.43793e-10, 1.452663e-10, 1.466679e-10, 
    1.463602e-10, 1.473933e-10, 1.446679e-10, 1.458072e-10, 1.453662e-10, 
    1.465175e-10, 1.440016e-10, 1.461428e-10, 1.434573e-10, 1.436916e-10, 
    1.444177e-10, 1.458847e-10, 1.462103e-10, 1.465585e-10, 1.463435e-10, 
    1.453038e-10, 1.451338e-10, 1.444e-10, 1.441978e-10, 1.436406e-10, 
    1.431802e-10, 1.436008e-10, 1.440433e-10, 1.453042e-10, 1.464459e-10, 
    1.476965e-10, 1.480035e-10, 1.494746e-10, 1.482766e-10, 1.502567e-10, 
    1.485725e-10, 1.514948e-10, 1.462672e-10, 1.485229e-10, 1.444507e-10, 
    1.448863e-10, 1.456761e-10, 1.474967e-10, 1.465121e-10, 1.476639e-10, 
    1.451271e-10, 1.438211e-10, 1.434841e-10, 1.428569e-10, 1.434985e-10, 
    1.434462e-10, 1.440616e-10, 1.438637e-10, 1.453461e-10, 1.445487e-10, 
    1.468206e-10, 1.476548e-10, 1.500252e-10, 1.514892e-10, 1.529879e-10, 
    1.536523e-10, 1.538548e-10, 1.539396e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24531.83, 24551.72, 24547.82, 24564.11, 24555.04, 24565.75, 24535.83, 
    24552.52, 24541.83, 24533.61, 24596.43, 24564.84, 24630.29, 24609.35, 
    24662.39, 24627, 24669.66, 24661.35, 24686.58, 24679.28, 24712.32, 
    24689.96, 24729.92, 24706.94, 24710.5, 24689.24, 24571.13, 24592.46, 
    24569.88, 24572.89, 24571.54, 24555.23, 24547.11, 24530.33, 24533.36, 
    24545.69, 24574.25, 24564.46, 24589.29, 24588.73, 24617.01, 24604.15, 
    24652.72, 24638.81, 24679.58, 24669.16, 24679.09, 24676.07, 24679.13, 
    24663.9, 24670.39, 24657.09, 24606.55, 24621.23, 24578.08, 24552.92, 
    24536.56, 24525.12, 24526.73, 24529.8, 24545.76, 24561.01, 24572.8, 
    24580.76, 24588.64, 24612.87, 24625.95, 24655.56, 24650.17, 24659.32, 
    24668.13, 24683.12, 24680.64, 24687.3, 24659.07, 24677.74, 24647.12, 
    24655.4, 24590.8, 24567.09, 24557.17, 24548.57, 24527.97, 24542.15, 
    24536.53, 24549.95, 24558.57, 24554.29, 24580.98, 24570.52, 24626.73, 
    24602.14, 24667.1, 24651.28, 24670.93, 24660.85, 24678.19, 24662.57, 
    24689.79, 24695.83, 24691.7, 24707.67, 24661.71, 24679.09, 24554.18, 
    24554.87, 24558.12, 24543.93, 24543.06, 24530.25, 24541.64, 24546.54, 
    24559.07, 24566.56, 24573.74, 24589.68, 24607.73, 24633.57, 24652.29, 
    24665.04, 24657.2, 24664.12, 24656.39, 24652.79, 24693.57, 24670.46, 
    24705.36, 24703.39, 24687.46, 24703.61, 24555.36, 24551.36, 24537.61, 
    24548.35, 24528.86, 24539.72, 24546.03, 24570.74, 24576.25, 24581.4, 
    24591.58, 24604.81, 24628.47, 24649.31, 24668.65, 24667.22, 24667.72, 
    24672.09, 24661.31, 24673.87, 24676, 24670.45, 24703.13, 24693.67, 
    24703.35, 24697.18, 24552.66, 24559.41, 24555.75, 24562.63, 24557.78, 
    24579.54, 24586.15, 24617.57, 24604.54, 24625.36, 24606.64, 24609.93, 
    24626.05, 24607.64, 24648.16, 24620.57, 24672.26, 24644.25, 24674.04, 
    24668.56, 24677.65, 24685.87, 24696.32, 24715.91, 24711.34, 24727.96, 
    24569.55, 24578.47, 24577.68, 24587.07, 24594.05, 24609.36, 24634.45, 
    24624.93, 24642.35, 24645.86, 24619.42, 24635.67, 24584.48, 24592.56, 
    24587.74, 24570.26, 24627.12, 24597.55, 24652.61, 24636.31, 24684.7, 
    24660.32, 24708.83, 24730.37, 24751.07, 24775.73, 24583.37, 24577.27, 
    24588.19, 24603.46, 24617.84, 24637.29, 24639.27, 24642.91, 24652.41, 
    24660.47, 24644.07, 24662.5, 24594.45, 24629.73, 24574.98, 24591.17, 
    24602.55, 24597.54, 24623.85, 24630.16, 24655.91, 24642.55, 24725.01, 
    24687.62, 24794.71, 24763.9, 24575.15, 24583.35, 24612.28, 24598.4, 
    24638.58, 24648.59, 24656.8, 24667.41, 24668.56, 24674.9, 24664.53, 
    24674.49, 24637.33, 24653.76, 24608.92, 24619.71, 24614.73, 24609.3, 
    24626.17, 24644.32, 24644.71, 24650.56, 24667.25, 24638.75, 24729.95, 
    24672.58, 24592.32, 24608.37, 24610.68, 24604.42, 24647.58, 24631.84, 
    24674.75, 24662.97, 24682.34, 24672.67, 24671.25, 24658.99, 24651.43, 
    24632.57, 24617.28, 24605.32, 24608.09, 24621.27, 24645.44, 24668.66, 
    24663.53, 24680.85, 24635.66, 24654.35, 24647.08, 24666.15, 24624.68, 
    24659.91, 24615.79, 24619.61, 24631.53, 24655.63, 24661.03, 24666.83, 
    24663.25, 24646.05, 24643.27, 24631.24, 24627.91, 24618.77, 24611.28, 
    24618.12, 24625.37, 24646.06, 24664.96, 24685.99, 24691.21, 24716.57, 
    24695.88, 24730.28, 24700.96, 24752.28, 24661.98, 24700.11, 24632.07, 
    24639.22, 24652.18, 24682.6, 24666.06, 24685.44, 24643.16, 24621.72, 
    24616.22, 24606.05, 24616.46, 24615.6, 24625.67, 24622.42, 24646.75, 
    24633.69, 24671.22, 24685.28, 24726.2, 24752.18, 24779.18, 24791.21, 
    24794.91, 24796.46 ;

 GC_ICE1 =
  17605.62, 17637.39, 17631.16, 17657.16, 17642.68, 17659.79, 17612.01, 
    17638.66, 17621.59, 17608.45, 17708.78, 17658.33, 17762.79, 17729.39, 
    17813.91, 17757.55, 17825.48, 17812.26, 17852.39, 17840.79, 17893.36, 
    17857.79, 17921.35, 17884.79, 17890.45, 17856.63, 17668.38, 17702.43, 
    17666.38, 17671.2, 17669.03, 17642.98, 17630.02, 17603.22, 17608.05, 
    17627.75, 17673.37, 17657.73, 17697.38, 17696.48, 17741.61, 17721.09, 
    17798.52, 17776.38, 17841.27, 17824.69, 17840.48, 17835.68, 17840.55, 
    17816.31, 17826.64, 17805.48, 17724.92, 17748.34, 17679.48, 17639.3, 
    17613.17, 17594.89, 17597.46, 17602.38, 17627.87, 17652.22, 17671.05, 
    17683.77, 17696.35, 17735, 17755.87, 17803.04, 17794.46, 17809.02, 
    17823.05, 17846.9, 17842.95, 17853.55, 17808.63, 17838.33, 17789.6, 
    17802.78, 17699.79, 17661.93, 17646.09, 17632.36, 17599.44, 17622.1, 
    17613.13, 17634.55, 17648.32, 17641.5, 17684.12, 17667.41, 17757.11, 
    17717.88, 17821.41, 17796.22, 17827.5, 17811.46, 17839.05, 17814.2, 
    17857.52, 17867.12, 17860.55, 17885.96, 17812.83, 17840.49, 17641.3, 
    17642.42, 17647.6, 17624.93, 17623.56, 17603.09, 17621.29, 17629.1, 
    17649.12, 17661.09, 17672.56, 17697.99, 17726.8, 17768.03, 17797.84, 
    17818.13, 17805.65, 17816.66, 17804.36, 17798.63, 17863.52, 17826.74, 
    17882.28, 17879.15, 17853.8, 17879.5, 17643.2, 17636.81, 17614.84, 
    17632.01, 17600.87, 17618.22, 17628.29, 17667.76, 17676.56, 17684.78, 
    17701.04, 17722.14, 17759.89, 17793.1, 17823.87, 17821.59, 17822.39, 
    17829.35, 17812.18, 17832.18, 17835.56, 17826.74, 17878.73, 17863.68, 
    17879.08, 17869.26, 17638.88, 17649.66, 17643.83, 17654.81, 17647.07, 
    17681.82, 17692.36, 17742.5, 17721.72, 17754.93, 17725.06, 17730.31, 
    17756.03, 17726.66, 17791.26, 17747.29, 17829.62, 17785.04, 17832.45, 
    17823.73, 17838.2, 17851.28, 17867.9, 17899.07, 17891.79, 17918.23, 
    17665.87, 17680.11, 17678.85, 17693.84, 17704.97, 17729.4, 17769.43, 
    17754.25, 17782.02, 17787.59, 17745.44, 17771.37, 17689.7, 17702.6, 
    17694.9, 17666.99, 17757.74, 17710.55, 17798.34, 17772.39, 17849.4, 
    17810.62, 17887.81, 17922.06, 17954.98, 17994.13, 17687.93, 17678.2, 
    17695.62, 17719.98, 17742.94, 17773.96, 17777.11, 17782.91, 17798.02, 
    17810.85, 17784.75, 17814.09, 17705.61, 17761.9, 17674.53, 17700.38, 
    17718.53, 17710.54, 17752.52, 17762.59, 17803.59, 17782.34, 17913.54, 
    17854.05, 18024.22, 17975.37, 17674.81, 17687.9, 17734.05, 17711.91, 
    17776.02, 17791.94, 17805.01, 17821.89, 17823.72, 17833.82, 17817.31, 
    17833.16, 17774.03, 17800.16, 17728.7, 17745.92, 17737.97, 17729.31, 
    17756.22, 17785.15, 17785.77, 17795.08, 17821.65, 17776.28, 17921.39, 
    17830.13, 17702.21, 17727.82, 17731.51, 17721.51, 17790.33, 17765.27, 
    17833.57, 17814.84, 17845.65, 17830.26, 17828.01, 17808.5, 17796.47, 
    17766.43, 17742.03, 17722.96, 17727.37, 17748.39, 17786.92, 17823.89, 
    17815.72, 17843.29, 17771.36, 17801.11, 17789.54, 17819.89, 17753.85, 
    17809.96, 17739.65, 17745.75, 17764.77, 17803.15, 17811.74, 17820.98, 
    17815.28, 17787.9, 17783.47, 17764.3, 17758.99, 17744.42, 17732.46, 
    17743.38, 17754.94, 17787.91, 17817.99, 17851.46, 17859.77, 17900.12, 
    17867.2, 17921.92, 17875.28, 17956.9, 17813.25, 17873.92, 17765.64, 
    17777.03, 17797.66, 17846.07, 17819.75, 17850.58, 17783.29, 17749.13, 
    17740.35, 17724.11, 17740.72, 17739.36, 17755.42, 17750.24, 17789.01, 
    17768.22, 17827.96, 17850.33, 17915.44, 17956.74, 17999.61, 18018.69, 
    18024.54, 18026.99 ;

 GC_LIQ1 =
  5232.783, 5234.812, 5234.414, 5236.075, 5235.15, 5236.243, 5233.19, 
    5234.893, 5233.803, 5232.963, 5239.384, 5236.15, 5242.863, 5240.711, 
    5246.213, 5242.525, 5246.975, 5246.105, 5248.749, 5247.983, 5251.45, 
    5249.104, 5253.299, 5250.884, 5251.258, 5249.027, 5236.792, 5238.976, 
    5236.664, 5236.972, 5236.833, 5235.169, 5234.341, 5232.629, 5232.938, 
    5234.196, 5237.111, 5236.111, 5238.65, 5238.592, 5241.499, 5240.177, 
    5245.201, 5243.746, 5248.015, 5246.923, 5247.963, 5247.647, 5247.968, 
    5246.371, 5247.052, 5245.659, 5240.423, 5241.932, 5237.501, 5234.934, 
    5233.265, 5232.098, 5232.262, 5232.576, 5234.204, 5235.759, 5236.962, 
    5237.775, 5238.583, 5241.073, 5242.417, 5245.499, 5244.935, 5245.892, 
    5246.815, 5248.386, 5248.126, 5248.825, 5245.866, 5247.822, 5244.615, 
    5245.481, 5238.805, 5236.38, 5235.368, 5234.49, 5232.388, 5233.835, 
    5233.262, 5234.63, 5235.51, 5235.074, 5237.798, 5236.73, 5242.498, 
    5239.97, 5246.707, 5245.05, 5247.108, 5246.052, 5247.869, 5246.232, 
    5249.086, 5249.719, 5249.286, 5250.961, 5246.143, 5247.964, 5235.062, 
    5235.133, 5235.464, 5234.016, 5233.928, 5232.621, 5233.783, 5234.283, 
    5235.562, 5236.326, 5237.059, 5238.689, 5240.544, 5243.201, 5245.157, 
    5246.491, 5245.67, 5246.395, 5245.585, 5245.208, 5249.481, 5247.058, 
    5250.718, 5250.512, 5248.841, 5250.535, 5235.183, 5234.775, 5233.372, 
    5234.468, 5232.479, 5233.587, 5234.23, 5236.752, 5237.315, 5237.84, 
    5238.886, 5240.245, 5242.676, 5244.845, 5246.869, 5246.719, 5246.772, 
    5247.229, 5246.1, 5247.417, 5247.64, 5247.058, 5250.484, 5249.492, 
    5250.508, 5249.86, 5234.907, 5235.596, 5235.223, 5235.925, 5235.43, 
    5237.651, 5238.327, 5241.556, 5240.217, 5242.357, 5240.433, 5240.771, 
    5242.428, 5240.536, 5244.724, 5241.864, 5247.248, 5244.315, 5247.435, 
    5246.86, 5247.813, 5248.675, 5249.77, 5251.827, 5251.346, 5253.093, 
    5236.631, 5237.542, 5237.461, 5238.422, 5239.139, 5240.712, 5243.291, 
    5242.313, 5244.116, 5244.483, 5241.746, 5243.417, 5238.155, 5238.986, 
    5238.491, 5236.703, 5242.538, 5239.499, 5245.189, 5243.484, 5248.551, 
    5245.997, 5251.083, 5253.346, 5255.528, 5258.146, 5238.042, 5237.419, 
    5238.537, 5240.105, 5241.584, 5243.587, 5243.794, 5244.175, 5245.168, 
    5246.012, 5244.296, 5246.225, 5239.18, 5242.806, 5237.185, 5238.843, 
    5240.012, 5239.498, 5242.202, 5242.851, 5245.535, 5244.137, 5252.783, 
    5248.858, 5260.191, 5256.88, 5237.203, 5238.04, 5241.012, 5239.586, 
    5243.722, 5244.769, 5245.628, 5246.739, 5246.859, 5247.524, 5246.437, 
    5247.481, 5243.591, 5245.31, 5240.667, 5241.776, 5241.265, 5240.706, 
    5242.44, 5244.323, 5244.363, 5244.975, 5246.723, 5243.739, 5253.302, 
    5247.281, 5238.961, 5240.611, 5240.848, 5240.204, 5244.663, 5243.023, 
    5247.508, 5246.274, 5248.304, 5247.29, 5247.142, 5245.857, 5245.066, 
    5243.098, 5241.526, 5240.297, 5240.582, 5241.936, 5244.439, 5246.87, 
    5246.332, 5248.148, 5243.416, 5245.372, 5244.611, 5246.607, 5242.287, 
    5245.954, 5241.373, 5241.765, 5242.991, 5245.506, 5246.071, 5246.679, 
    5246.303, 5244.503, 5244.212, 5242.961, 5242.619, 5241.68, 5240.91, 
    5241.613, 5242.357, 5244.504, 5246.482, 5248.687, 5249.234, 5251.896, 
    5249.724, 5253.337, 5250.257, 5255.655, 5246.17, 5250.167, 5243.047, 
    5243.789, 5245.145, 5248.332, 5246.598, 5248.629, 5244.2, 5241.983, 
    5241.417, 5240.372, 5241.441, 5241.354, 5242.388, 5242.055, 5244.576, 
    5243.213, 5247.138, 5248.613, 5252.908, 5255.645, 5258.517, 5259.814, 
    5260.213, 5260.38 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.956448e-09, 8.995829e-09, 8.988173e-09, 9.019937e-09, 9.002316e-09, 
    9.023116e-09, 8.964432e-09, 8.997393e-09, 8.976351e-09, 8.959993e-09, 
    9.081578e-09, 9.021353e-09, 9.144131e-09, 9.105723e-09, 9.202203e-09, 
    9.138154e-09, 9.215118e-09, 9.200354e-09, 9.244784e-09, 9.232056e-09, 
    9.288887e-09, 9.250659e-09, 9.318345e-09, 9.279757e-09, 9.285794e-09, 
    9.249399e-09, 9.033473e-09, 9.074081e-09, 9.031067e-09, 9.036857e-09, 
    9.034259e-09, 9.00268e-09, 8.986768e-09, 8.953438e-09, 8.959488e-09, 
    8.983968e-09, 9.039462e-09, 9.020623e-09, 9.068097e-09, 9.067025e-09, 
    9.119877e-09, 9.096047e-09, 9.184878e-09, 9.159631e-09, 9.232587e-09, 
    9.21424e-09, 9.231726e-09, 9.226423e-09, 9.231795e-09, 9.204886e-09, 
    9.216415e-09, 9.192736e-09, 9.100511e-09, 9.127616e-09, 9.046775e-09, 
    8.998167e-09, 8.965878e-09, 8.942965e-09, 8.946205e-09, 8.95238e-09, 
    8.984111e-09, 9.013944e-09, 9.036679e-09, 9.051886e-09, 9.066871e-09, 
    9.112229e-09, 9.136234e-09, 9.189984e-09, 9.180282e-09, 9.196716e-09, 
    9.212415e-09, 9.238772e-09, 9.234433e-09, 9.246046e-09, 9.196282e-09, 
    9.229355e-09, 9.174758e-09, 9.189691e-09, 9.070948e-09, 9.025705e-09, 
    9.006478e-09, 8.989645e-09, 8.948695e-09, 8.976975e-09, 8.965827e-09, 
    8.992347e-09, 9.009199e-09, 9.000864e-09, 9.052303e-09, 9.032305e-09, 
    9.137657e-09, 9.092279e-09, 9.210583e-09, 9.182274e-09, 9.217369e-09, 
    9.199461e-09, 9.230146e-09, 9.202529e-09, 9.250367e-09, 9.260784e-09, 
    9.253665e-09, 9.281009e-09, 9.200998e-09, 9.231726e-09, 9.00063e-09, 
    9.00199e-09, 9.008323e-09, 8.980487e-09, 8.978783e-09, 8.953272e-09, 
    8.975971e-09, 8.985638e-09, 9.010176e-09, 9.02469e-09, 9.038487e-09, 
    9.068823e-09, 9.102703e-09, 9.150076e-09, 9.184109e-09, 9.206922e-09, 
    9.192934e-09, 9.205284e-09, 9.191478e-09, 9.185007e-09, 9.256881e-09, 
    9.216523e-09, 9.277076e-09, 9.273725e-09, 9.246322e-09, 9.274102e-09, 
    9.002945e-09, 8.995122e-09, 8.967964e-09, 8.989217e-09, 8.950494e-09, 
    8.972171e-09, 8.984634e-09, 9.032724e-09, 9.043289e-09, 9.053086e-09, 
    9.072435e-09, 9.097267e-09, 9.140829e-09, 9.178729e-09, 9.213328e-09, 
    9.210792e-09, 9.211685e-09, 9.219415e-09, 9.200269e-09, 9.222558e-09, 
    9.226299e-09, 9.216517e-09, 9.273276e-09, 9.257061e-09, 9.273654e-09, 
    9.263096e-09, 8.997665e-09, 9.010827e-09, 9.003715e-09, 9.017089e-09, 
    9.007668e-09, 9.049564e-09, 9.062125e-09, 9.120901e-09, 9.096778e-09, 
    9.135169e-09, 9.100678e-09, 9.10679e-09, 9.136422e-09, 9.102542e-09, 
    9.17664e-09, 9.126405e-09, 9.219715e-09, 9.169552e-09, 9.222858e-09, 
    9.213178e-09, 9.229205e-09, 9.24356e-09, 9.261618e-09, 9.294939e-09, 
    9.287223e-09, 9.315088e-09, 9.030448e-09, 9.047521e-09, 9.046017e-09, 
    9.063883e-09, 9.077096e-09, 9.105732e-09, 9.151662e-09, 9.13439e-09, 
    9.166097e-09, 9.172463e-09, 9.124292e-09, 9.153869e-09, 9.058946e-09, 
    9.074284e-09, 9.065151e-09, 9.031796e-09, 9.138371e-09, 9.083678e-09, 
    9.184672e-09, 9.155043e-09, 9.241513e-09, 9.19851e-09, 9.282975e-09, 
    9.319085e-09, 9.353066e-09, 9.392782e-09, 9.056838e-09, 9.045237e-09, 
    9.066008e-09, 9.094744e-09, 9.121405e-09, 9.15685e-09, 9.160477e-09, 
    9.167117e-09, 9.184316e-09, 9.198778e-09, 9.169217e-09, 9.202403e-09, 
    9.077842e-09, 9.143118e-09, 9.040853e-09, 9.071648e-09, 9.09305e-09, 
    9.083661e-09, 9.132416e-09, 9.143907e-09, 9.190603e-09, 9.166464e-09, 
    9.310174e-09, 9.246593e-09, 9.423018e-09, 9.373716e-09, 9.041185e-09, 
    9.056797e-09, 9.111135e-09, 9.085281e-09, 9.159216e-09, 9.177414e-09, 
    9.192209e-09, 9.211121e-09, 9.213162e-09, 9.224367e-09, 9.206006e-09, 
    9.223642e-09, 9.156926e-09, 9.186739e-09, 9.104923e-09, 9.124837e-09, 
    9.115675e-09, 9.105627e-09, 9.136641e-09, 9.169683e-09, 9.170388e-09, 
    9.180982e-09, 9.210841e-09, 9.159516e-09, 9.318383e-09, 9.220273e-09, 
    9.073822e-09, 9.103895e-09, 9.10819e-09, 9.09654e-09, 9.175591e-09, 
    9.146948e-09, 9.224094e-09, 9.203244e-09, 9.237406e-09, 9.220431e-09, 
    9.217933e-09, 9.19613e-09, 9.182556e-09, 9.148262e-09, 9.120358e-09, 
    9.09823e-09, 9.103375e-09, 9.127682e-09, 9.171703e-09, 9.213347e-09, 
    9.204226e-09, 9.23481e-09, 9.153855e-09, 9.187802e-09, 9.174682e-09, 
    9.208891e-09, 9.133932e-09, 9.197768e-09, 9.117614e-09, 9.124642e-09, 
    9.14638e-09, 9.190105e-09, 9.199777e-09, 9.210106e-09, 9.203732e-09, 
    9.172821e-09, 9.167756e-09, 9.145851e-09, 9.139804e-09, 9.123112e-09, 
    9.109293e-09, 9.121919e-09, 9.135179e-09, 9.172834e-09, 9.206768e-09, 
    9.243765e-09, 9.252818e-09, 9.296047e-09, 9.260859e-09, 9.318929e-09, 
    9.269561e-09, 9.355018e-09, 9.201465e-09, 9.268106e-09, 9.147368e-09, 
    9.160376e-09, 9.183903e-09, 9.237863e-09, 9.208731e-09, 9.242799e-09, 
    9.167557e-09, 9.128521e-09, 9.11842e-09, 9.099575e-09, 9.118851e-09, 
    9.117283e-09, 9.135727e-09, 9.1298e-09, 9.174084e-09, 9.150297e-09, 
    9.217871e-09, 9.24253e-09, 9.312169e-09, 9.354859e-09, 9.398312e-09, 
    9.417497e-09, 9.423337e-09, 9.425777e-09 ;

 H2OCAN =
  0.05992912, 0.05991415, 0.059917, 0.05990504, 0.05991157, 0.05990382, 
    0.05992595, 0.05991368, 0.05992144, 0.05992759, 0.05988215, 0.05990448, 
    0.05985782, 0.0598722, 0.05983553, 0.05986024, 0.05983046, 0.05983594, 
    0.05981864, 0.05982359, 0.05980198, 0.05981635, 0.05979019, 0.05980526, 
    0.05980302, 0.05981687, 0.05989969, 0.059885, 0.05990063, 0.05989852, 
    0.0598994, 0.05991154, 0.05991784, 0.05993005, 0.05992778, 0.05991869, 
    0.05989756, 0.05990455, 0.0598863, 0.05988671, 0.05986678, 0.05987578, 
    0.0598419, 0.0598515, 0.05982338, 0.05983054, 0.05982377, 0.05982578, 
    0.05982374, 0.05983421, 0.05982975, 0.05983884, 0.05987415, 0.05986391, 
    0.05989467, 0.05991368, 0.05992547, 0.05993403, 0.05993283, 0.05993059, 
    0.05991865, 0.0599071, 0.05989837, 0.05989255, 0.05988677, 0.05987026, 
    0.05986082, 0.05984011, 0.0598436, 0.05983748, 0.05983123, 0.05982107, 
    0.0598227, 0.05981828, 0.05983745, 0.05982482, 0.05984564, 0.05984, 
    0.05988625, 0.05990262, 0.05991045, 0.05991649, 0.05993192, 0.05992133, 
    0.05992553, 0.0599153, 0.05990893, 0.05991204, 0.05989239, 0.05990009, 
    0.05986026, 0.05987737, 0.05983196, 0.05984286, 0.0598293, 0.05983618, 
    0.05982446, 0.05983501, 0.05981654, 0.05981262, 0.05981532, 0.05980457, 
    0.05983562, 0.05982387, 0.05991217, 0.05991167, 0.05990922, 0.05992002, 
    0.05992062, 0.05993016, 0.05992158, 0.059918, 0.05990847, 0.05990302, 
    0.05989776, 0.05988613, 0.05987347, 0.05985539, 0.05984217, 0.0598333, 
    0.05983867, 0.05983394, 0.05983927, 0.05984172, 0.05981416, 0.05982977, 
    0.05980612, 0.0598074, 0.05981821, 0.05980725, 0.0599113, 0.05991422, 
    0.05992465, 0.05991649, 0.05993119, 0.0599231, 0.05991852, 0.05990016, 
    0.05989585, 0.05989219, 0.0598847, 0.05987532, 0.05985888, 0.05984434, 
    0.05983082, 0.05983179, 0.05983146, 0.05982854, 0.05983591, 0.05982732, 
    0.05982598, 0.05982964, 0.05980758, 0.05981389, 0.05980743, 0.05981151, 
    0.05991324, 0.05990829, 0.05991099, 0.05990597, 0.05990959, 0.05989377, 
    0.05988901, 0.05986665, 0.05987556, 0.05986108, 0.05987401, 0.05987179, 
    0.05986105, 0.05987325, 0.05984535, 0.05986468, 0.05982843, 0.0598483, 
    0.0598272, 0.05983088, 0.05982468, 0.05981922, 0.05981213, 0.05979931, 
    0.05980225, 0.05979131, 0.05990079, 0.05989442, 0.05989479, 0.05988797, 
    0.05988301, 0.05987206, 0.05985465, 0.05986114, 0.059849, 0.05984662, 
    0.05986495, 0.0598539, 0.05989, 0.05988435, 0.05988755, 0.0599004, 
    0.05985992, 0.05988075, 0.05984199, 0.05985332, 0.05982002, 0.05983685, 
    0.0598039, 0.05979019, 0.05977627, 0.05976099, 0.05989072, 0.05989508, 
    0.0598871, 0.05987654, 0.05986618, 0.05985266, 0.05985117, 0.05984869, 
    0.059842, 0.05983646, 0.05984809, 0.05983504, 0.05988344, 0.05985801, 
    0.05989691, 0.05988539, 0.05987707, 0.05988052, 0.05986183, 0.05985749, 
    0.05983981, 0.05984886, 0.05979376, 0.05981834, 0.05974861, 0.05976845, 
    0.05989665, 0.05989065, 0.05987021, 0.05987987, 0.05985165, 0.05984475, 
    0.05983895, 0.05983184, 0.05983092, 0.05982667, 0.05983366, 0.05982687, 
    0.05985263, 0.05984113, 0.05987231, 0.05986486, 0.05986822, 0.05987205, 
    0.05986025, 0.05984796, 0.05984738, 0.05984348, 0.05983301, 0.05985153, 
    0.05979116, 0.05982921, 0.05988414, 0.05987313, 0.05987118, 0.05987551, 
    0.05984545, 0.05985642, 0.05982672, 0.05983473, 0.05982152, 0.05982812, 
    0.0598291, 0.05983748, 0.05984275, 0.05985598, 0.0598666, 0.05987484, 
    0.05987291, 0.05986384, 0.05984713, 0.05983098, 0.05983458, 0.05982252, 
    0.05985372, 0.05984086, 0.05984595, 0.0598326, 0.05986138, 0.05983787, 
    0.05986748, 0.05986483, 0.05985663, 0.0598402, 0.05983607, 0.05983223, 
    0.05983453, 0.05984665, 0.05984848, 0.05985675, 0.05985919, 0.05986538, 
    0.05987065, 0.05986591, 0.059861, 0.05984651, 0.05983354, 0.05981919, 
    0.05981554, 0.05979943, 0.05981299, 0.05979101, 0.05981039, 0.05977641, 
    0.05983603, 0.0598103, 0.05985615, 0.05985118, 0.05984252, 0.05982178, 
    0.05983266, 0.05981978, 0.05984853, 0.05986368, 0.0598672, 0.0598744, 
    0.05986704, 0.05986762, 0.05986058, 0.05986282, 0.05984602, 0.05985505, 
    0.05982922, 0.0598198, 0.05979257, 0.05977592, 0.05975832, 0.05975068, 
    0.05974833, 0.05974736 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  3.78638, 3.799462, 3.796917, 3.807488, 3.801623, 3.808548, 3.789031, 
    3.799981, 3.792989, 3.787558, 3.828065, 3.807961, 3.849054, 3.836164, 
    3.868615, 3.847044, 3.872977, 3.867995, 3.883013, 3.878706, 3.897955, 
    3.885002, 3.907969, 3.894861, 3.896908, 3.884574, 3.812004, 3.825556, 
    3.811201, 3.813131, 3.812266, 3.801743, 3.796446, 3.785384, 3.787391, 
    3.795518, 3.813999, 3.80772, 3.823569, 3.82321, 3.840912, 3.832923, 
    3.862776, 3.854273, 3.878886, 3.872684, 3.878594, 3.876801, 3.878617, 
    3.869525, 3.873418, 3.865426, 3.834417, 3.843509, 3.816442, 3.800234, 
    3.78951, 3.781912, 3.782985, 3.785031, 3.795565, 3.805495, 3.813075, 
    3.818151, 3.823159, 3.838338, 3.8464, 3.864495, 3.861228, 3.866766, 
    3.872067, 3.880976, 3.879509, 3.883438, 3.866622, 3.87779, 3.859367, 
    3.864399, 3.824507, 3.809414, 3.803001, 3.797406, 3.78381, 3.793194, 
    3.789492, 3.798307, 3.803914, 3.801141, 3.81829, 3.811615, 3.846879, 
    3.831658, 3.871449, 3.861898, 3.873741, 3.867695, 3.878058, 3.868731, 
    3.884902, 3.888428, 3.886018, 3.895288, 3.868214, 3.878592, 3.801062, 
    3.801514, 3.803623, 3.794361, 3.793795, 3.785328, 3.792863, 3.796074, 
    3.80424, 3.809075, 3.813677, 3.82381, 3.83515, 3.851055, 3.862517, 
    3.870214, 3.865494, 3.86966, 3.865002, 3.862821, 3.887105, 3.873454, 
    3.893954, 3.892817, 3.883531, 3.892946, 3.801832, 3.79923, 3.790203, 
    3.797266, 3.784407, 3.791599, 3.795738, 3.811751, 3.81528, 3.81855, 
    3.825019, 3.833331, 3.847947, 3.860702, 3.872377, 3.871521, 3.871822, 
    3.874432, 3.867967, 3.875494, 3.876757, 3.873453, 3.892665, 3.887169, 
    3.892793, 3.889215, 3.800076, 3.804457, 3.802089, 3.806542, 3.803403, 
    3.817371, 3.821566, 3.841252, 3.833167, 3.846045, 3.834474, 3.836522, 
    3.84646, 3.8351, 3.859995, 3.843098, 3.874533, 3.857605, 3.875596, 
    3.872326, 3.877742, 3.882597, 3.888713, 3.900014, 3.897395, 3.906863, 
    3.810996, 3.81669, 3.816191, 3.822159, 3.826577, 3.836169, 3.851591, 
    3.845786, 3.85645, 3.858593, 3.842396, 3.852332, 3.820507, 3.825632, 
    3.822582, 3.811443, 3.84712, 3.828776, 3.862706, 3.852729, 3.881904, 
    3.867371, 3.895954, 3.908216, 3.919795, 3.933347, 3.819804, 3.815931, 
    3.82287, 3.832482, 3.841425, 3.853336, 3.854558, 3.856792, 3.862588, 
    3.867465, 3.857497, 3.868688, 3.826816, 3.848716, 3.814465, 3.82475, 
    3.831916, 3.828774, 3.845124, 3.848985, 3.864704, 3.856573, 3.905185, 
    3.883619, 3.943696, 3.926835, 3.814578, 3.819792, 3.837978, 3.829317, 
    3.854134, 3.86026, 3.865249, 3.871629, 3.87232, 3.876105, 3.869904, 
    3.875861, 3.853361, 3.863404, 3.835898, 3.842577, 3.839504, 3.836134, 
    3.846543, 3.857653, 3.857894, 3.861461, 3.87152, 3.854234, 3.907968, 
    3.874708, 3.825483, 3.835548, 3.836992, 3.833089, 3.859646, 3.850006, 
    3.876014, 3.868972, 3.880516, 3.874776, 3.873932, 3.866571, 3.861993, 
    3.850447, 3.841073, 3.833655, 3.835379, 3.843532, 3.858334, 3.872381, 
    3.8693, 3.879637, 3.85233, 3.86376, 3.859338, 3.870878, 3.845631, 
    3.86711, 3.840155, 3.842513, 3.849815, 3.864533, 3.867802, 3.871287, 
    3.869137, 3.858711, 3.857007, 3.849638, 3.847604, 3.842, 3.837364, 
    3.841599, 3.846049, 3.858717, 3.870159, 3.882665, 3.885732, 3.900383, 
    3.888448, 3.908153, 3.891387, 3.920448, 3.868363, 3.890903, 3.850149, 
    3.854524, 3.862444, 3.880664, 3.870823, 3.882336, 3.856941, 3.843811, 
    3.840425, 3.834105, 3.840569, 3.840044, 3.846236, 3.844246, 3.859138, 
    3.851133, 3.873909, 3.882246, 3.905869, 3.920402, 3.935244, 3.941808, 
    3.943807, 3.944643,
  3.296503, 3.30925, 3.306771, 3.31707, 3.311357, 3.318104, 3.299088, 
    3.309754, 3.302943, 3.297653, 3.336786, 3.317532, 3.356738, 3.344494, 
    3.375332, 3.354825, 3.379481, 3.374749, 3.389031, 3.384935, 3.403237, 
    3.390923, 3.412769, 3.400298, 3.402243, 3.390516, 3.321474, 3.334403, 
    3.320692, 3.322572, 3.32173, 3.311472, 3.306307, 3.295536, 3.29749, 
    3.305406, 3.323417, 3.3173, 3.332532, 3.332192, 3.349006, 3.341416, 
    3.369786, 3.361705, 3.385106, 3.379208, 3.384827, 3.383124, 3.38485, 
    3.376202, 3.379905, 3.372306, 3.342835, 3.351472, 3.325761, 3.309997, 
    3.299553, 3.292152, 3.293198, 3.29519, 3.305452, 3.315131, 3.32252, 
    3.327387, 3.332143, 3.34655, 3.354217, 3.371417, 3.368316, 3.373577, 
    3.378622, 3.387093, 3.385699, 3.389433, 3.373444, 3.384061, 3.366548, 
    3.37133, 3.333406, 3.318951, 3.312694, 3.307246, 3.294001, 3.303142, 
    3.299536, 3.308126, 3.31359, 3.310888, 3.327518, 3.321096, 3.354671, 
    3.340212, 3.378033, 3.368953, 3.380213, 3.374465, 3.384317, 3.375449, 
    3.390827, 3.394179, 3.391887, 3.400707, 3.374958, 3.384825, 3.310811, 
    3.311252, 3.313307, 3.304278, 3.303728, 3.29548, 3.302821, 3.305948, 
    3.313909, 3.31862, 3.323106, 3.33276, 3.343529, 3.358643, 3.36954, 
    3.376859, 3.372372, 3.376333, 3.371904, 3.369831, 3.39292, 3.379937, 
    3.399438, 3.398358, 3.389521, 3.398479, 3.311561, 3.309026, 3.300229, 
    3.307112, 3.294584, 3.301589, 3.30562, 3.321226, 3.32466, 3.327764, 
    3.333909, 3.341804, 3.35569, 3.367813, 3.378917, 3.378103, 3.378389, 
    3.38087, 3.374723, 3.38188, 3.383079, 3.379939, 3.398213, 3.392985, 
    3.398335, 3.39493, 3.309851, 3.314119, 3.311812, 3.31615, 3.313091, 
    3.32664, 3.330624, 3.349324, 3.341647, 3.353881, 3.342891, 3.344834, 
    3.354268, 3.343486, 3.367138, 3.351076, 3.380966, 3.364861, 3.381977, 
    3.378868, 3.384019, 3.388634, 3.394453, 3.405201, 3.402711, 3.41172, 
    3.320493, 3.325996, 3.325526, 3.331193, 3.335387, 3.344501, 3.359154, 
    3.35364, 3.363775, 3.36581, 3.350418, 3.359856, 3.329622, 3.334485, 
    3.331593, 3.320927, 3.354902, 3.337472, 3.36972, 3.360236, 3.387975, 
    3.374151, 3.40134, 3.413, 3.42403, 3.436924, 3.328955, 3.325279, 
    3.331869, 3.340993, 3.349494, 3.360813, 3.361976, 3.364099, 3.369609, 
    3.374246, 3.364764, 3.375409, 3.335603, 3.356421, 3.323874, 3.333647, 
    3.340457, 3.337474, 3.353011, 3.356679, 3.371617, 3.363892, 3.410114, 
    3.389601, 3.446787, 3.430727, 3.323985, 3.328945, 3.346216, 3.337991, 
    3.361573, 3.367395, 3.37214, 3.378203, 3.378862, 3.38246, 3.376565, 
    3.382229, 3.360837, 3.370384, 3.344245, 3.350589, 3.347671, 3.344469, 
    3.354359, 3.364912, 3.365147, 3.368535, 3.378081, 3.361669, 3.412752, 
    3.381116, 3.334351, 3.343904, 3.345282, 3.341575, 3.366811, 3.357648, 
    3.382374, 3.375679, 3.386656, 3.381197, 3.380394, 3.373396, 3.369043, 
    3.358066, 3.349159, 3.342114, 3.343752, 3.351494, 3.365561, 3.378918, 
    3.375987, 3.385821, 3.359858, 3.37072, 3.366516, 3.37749, 3.353491, 
    3.373891, 3.348289, 3.35053, 3.357467, 3.371452, 3.374566, 3.377877, 
    3.375836, 3.36592, 3.364302, 3.3573, 3.355364, 3.350043, 3.345637, 
    3.34966, 3.353886, 3.365928, 3.376805, 3.388698, 3.391618, 3.405543, 
    3.394191, 3.412927, 3.396974, 3.424637, 3.37509, 3.396524, 3.357786, 
    3.361944, 3.369467, 3.38679, 3.377438, 3.388381, 3.364239, 3.351757, 
    3.348545, 3.34254, 3.348683, 3.348183, 3.354068, 3.352176, 3.366329, 
    3.358721, 3.380371, 3.388297, 3.410772, 3.424601, 3.438739, 3.44499, 
    3.446895, 3.447692,
  3.020753, 3.034852, 3.032108, 3.043507, 3.03718, 3.04465, 3.023607, 
    3.035413, 3.027873, 3.02202, 3.065719, 3.044017, 3.088386, 3.074456, 
    3.109537, 3.086215, 3.114164, 3.108863, 3.124689, 3.120171, 3.140379, 
    3.126776, 3.150894, 3.137127, 3.139277, 3.126328, 3.048376, 3.063011, 
    3.04751, 3.049594, 3.048659, 3.03731, 3.031603, 3.019677, 3.02184, 
    3.030601, 3.050531, 3.043755, 3.060854, 3.060467, 3.079584, 3.070954, 
    3.103217, 3.094022, 3.120359, 3.113855, 3.120053, 3.118173, 3.120078, 
    3.110517, 3.114625, 3.106083, 3.072569, 3.082391, 3.053165, 3.03569, 
    3.024125, 3.015937, 3.017094, 3.019299, 3.030652, 3.041355, 3.04953, 
    3.055007, 3.060412, 3.076811, 3.085518, 3.105078, 3.101542, 3.107534, 
    3.113208, 3.122553, 3.121014, 3.125136, 3.107377, 3.119212, 3.099529, 
    3.104972, 3.06188, 3.045582, 3.038672, 3.032635, 3.017983, 3.028096, 
    3.024106, 3.033604, 3.039651, 3.036659, 3.055157, 3.047956, 3.086035, 
    3.06959, 3.11256, 3.102268, 3.114963, 3.108537, 3.119492, 3.109657, 
    3.126672, 3.130374, 3.127843, 3.137573, 3.109098, 3.120053, 3.036575, 
    3.037063, 3.039336, 3.029353, 3.028743, 3.019618, 3.027737, 3.031199, 
    3.040002, 3.045217, 3.050181, 3.061116, 3.073362, 3.090547, 3.102936, 
    3.111261, 3.106155, 3.110663, 3.105624, 3.103264, 3.128986, 3.114663, 
    3.136173, 3.13498, 3.125234, 3.135114, 3.037406, 3.0346, 3.024871, 
    3.032482, 3.018625, 3.026376, 3.030839, 3.048106, 3.05191, 3.055439, 
    3.06242, 3.071395, 3.087187, 3.100975, 3.113532, 3.112634, 3.11295, 
    3.115688, 3.108832, 3.116802, 3.118128, 3.114662, 3.13482, 3.129051, 
    3.134954, 3.131197, 3.035511, 3.040236, 3.037682, 3.042485, 3.039101, 
    3.054169, 3.058698, 3.079955, 3.071218, 3.085132, 3.07263, 3.074842, 
    3.085585, 3.073305, 3.100214, 3.081951, 3.115794, 3.097631, 3.116909, 
    3.113479, 3.11916, 3.124254, 3.130671, 3.142538, 3.139787, 3.149731, 
    3.047288, 3.053434, 3.052893, 3.059333, 3.064103, 3.07446, 3.091124, 
    3.08485, 3.096375, 3.098693, 3.081186, 3.091926, 3.057552, 3.063086, 
    3.059791, 3.047772, 3.086294, 3.06648, 3.103141, 3.092353, 3.123527, 
    3.108189, 3.138274, 3.151157, 3.163321, 3.177577, 3.056792, 3.052612, 
    3.0601, 3.070482, 3.080138, 3.09301, 3.09433, 3.096746, 3.103012, 
    3.108288, 3.09751, 3.109611, 3.06437, 3.088019, 3.051032, 3.062135, 
    3.069869, 3.066475, 3.084133, 3.088306, 3.105304, 3.096509, 3.147973, 
    3.125329, 3.188466, 3.170727, 3.051152, 3.056778, 3.076416, 3.067061, 
    3.093871, 3.100497, 3.105891, 3.11275, 3.113473, 3.117444, 3.110927, 
    3.117187, 3.093038, 3.103896, 3.074167, 3.081383, 3.078062, 3.074422, 
    3.085667, 3.09768, 3.097937, 3.101796, 3.112646, 3.09398, 3.150903, 
    3.115988, 3.062921, 3.073793, 3.075349, 3.071133, 3.099832, 3.089411, 
    3.117347, 3.109918, 3.122069, 3.116048, 3.115163, 3.107321, 3.10237, 
    3.089888, 3.079759, 3.071744, 3.073606, 3.082415, 3.098416, 3.113538, 
    3.110276, 3.121148, 3.091922, 3.104282, 3.0995, 3.111961, 3.084683, 
    3.107916, 3.078765, 3.081313, 3.089204, 3.105122, 3.108652, 3.11239, 
    3.110096, 3.098823, 3.096979, 3.089012, 3.086815, 3.080758, 3.07575, 
    3.080325, 3.085135, 3.098828, 3.111204, 3.124326, 3.127543, 3.142931, 
    3.130399, 3.151098, 3.133491, 3.164017, 3.109267, 3.132976, 3.089564, 
    3.094293, 3.10286, 3.122229, 3.111904, 3.123982, 3.096907, 3.082719, 
    3.079057, 3.072231, 3.079213, 3.078644, 3.085335, 3.083184, 3.099283, 
    3.090628, 3.115141, 3.123887, 3.148688, 3.163962, 3.179569, 3.186477, 
    3.188581, 3.189461,
  2.893865, 2.909182, 2.906199, 2.91859, 2.911711, 2.919832, 2.896965, 
    2.909792, 2.901598, 2.895241, 2.942753, 2.919143, 2.967429, 2.952258, 
    2.990482, 2.965065, 2.995516, 2.989745, 3.006982, 3.002058, 3.024093, 
    3.009256, 3.035564, 3.020544, 3.02289, 3.008768, 2.923882, 2.939806, 
    2.92294, 2.925207, 2.924189, 2.911853, 2.905653, 2.892696, 2.895045, 
    2.904562, 2.926226, 2.918857, 2.937453, 2.937032, 2.957841, 2.948445, 
    2.98359, 2.973568, 3.002263, 2.995177, 3.00193, 2.999881, 3.001957, 
    2.99155, 2.996017, 2.986714, 2.950203, 2.960898, 2.92909, 2.910094, 
    2.897527, 2.888635, 2.889891, 2.892286, 2.904618, 2.916248, 2.925136, 
    2.931093, 2.936972, 2.954825, 2.964305, 2.98562, 2.981763, 2.988298, 
    2.994473, 3.004655, 3.002977, 3.00747, 2.988125, 3.001014, 2.979569, 
    2.985502, 2.938576, 2.920844, 2.913335, 2.906772, 2.890857, 2.901841, 
    2.897507, 2.907825, 2.914396, 2.911144, 2.931256, 2.923425, 2.964868, 
    2.946962, 2.993767, 2.982555, 2.996385, 2.989389, 3.00132, 2.990611, 
    3.009143, 3.01318, 3.010421, 3.021029, 2.990002, 3.001931, 2.911053, 
    2.911584, 2.914054, 2.903207, 2.902544, 2.892632, 2.90145, 2.905212, 
    2.914777, 2.920447, 2.925844, 2.937739, 2.951067, 2.969783, 2.983284, 
    2.992354, 2.986792, 2.991708, 2.986213, 2.98364, 3.011667, 2.996058, 
    3.019502, 3.018201, 3.007577, 3.018347, 2.911956, 2.908906, 2.898337, 
    2.906605, 2.891554, 2.899972, 2.904821, 2.923589, 2.927724, 2.931564, 
    2.939157, 2.948925, 2.966122, 2.981147, 2.994825, 2.993847, 2.994191, 
    2.997174, 2.989711, 2.998388, 2.999833, 2.996056, 3.018027, 3.011737, 
    3.018173, 3.014076, 2.909897, 2.915031, 2.912256, 2.917477, 2.913798, 
    2.930184, 2.93511, 2.958246, 2.948733, 2.963883, 2.950269, 2.952678, 
    2.964381, 2.951003, 2.980318, 2.960421, 2.99729, 2.977504, 2.998504, 
    2.994767, 3.000956, 3.006508, 3.013503, 3.026446, 3.023445, 3.034294, 
    2.922698, 2.929383, 2.928793, 2.935799, 2.940989, 2.952261, 2.97041, 
    2.963575, 2.976132, 2.978658, 2.959584, 2.971285, 2.933862, 2.939884, 
    2.936297, 2.923226, 2.96515, 2.943577, 2.983508, 2.97175, 3.005716, 
    2.989012, 3.021794, 3.035853, 3.049129, 3.064706, 2.933035, 2.928488, 
    2.936633, 2.947932, 2.958445, 2.972466, 2.973903, 2.976537, 2.983366, 
    2.989118, 2.977371, 2.990561, 2.941284, 2.967028, 2.92677, 2.938849, 
    2.947265, 2.94357, 2.962794, 2.96734, 2.985866, 2.976277, 3.032379, 
    3.007683, 3.076607, 3.057221, 2.9269, 2.933019, 2.954392, 2.944207, 
    2.973403, 2.980624, 2.986504, 2.993974, 2.994761, 2.999087, 2.991996, 
    2.998807, 2.972496, 2.984329, 2.951942, 2.9598, 2.956183, 2.952219, 
    2.964465, 2.977556, 2.977834, 2.982042, 2.993868, 2.973522, 3.035581, 
    2.997508, 2.939702, 2.951538, 2.95323, 2.948639, 2.9799, 2.968544, 
    2.998981, 2.990896, 3.004127, 2.997566, 2.996603, 2.988064, 2.982667, 
    2.969064, 2.958031, 2.949304, 2.951332, 2.960924, 2.978357, 2.994833, 
    2.991287, 3.003123, 2.971279, 2.984752, 2.979539, 2.993114, 2.963394, 
    2.988719, 2.956948, 2.959723, 2.968319, 2.985668, 2.989515, 2.993583, 
    2.99109, 2.978801, 2.97679, 2.968109, 2.965716, 2.959118, 2.953665, 
    2.958647, 2.963887, 2.978805, 2.992295, 3.006587, 3.010092, 3.026879, 
    3.01321, 3.035794, 3.016587, 3.049895, 2.990189, 3.016021, 2.96871, 
    2.973863, 2.983203, 3.004304, 2.993052, 3.006214, 2.976712, 2.961256, 
    2.957266, 2.949835, 2.957436, 2.956817, 2.964103, 2.96176, 2.979302, 
    2.969869, 2.996578, 3.00611, 3.033156, 3.049832, 3.06688, 3.074431, 
    3.076732, 3.077694,
  2.944312, 2.960424, 2.957285, 2.970329, 2.963086, 2.971638, 2.947571, 
    2.961066, 2.952444, 2.945758, 2.995805, 2.970912, 3.021869, 3.005837, 
    3.046266, 3.01937, 3.051717, 3.045485, 3.064276, 3.058881, 3.082962, 
    3.066768, 3.095155, 3.079147, 3.081684, 3.066233, 2.975904, 2.992695, 
    2.974913, 2.977301, 2.976228, 2.963236, 2.95671, 2.943083, 2.945552, 
    2.955562, 2.978375, 2.970611, 2.990212, 2.989768, 3.011735, 3.001812, 
    3.038967, 3.028361, 3.059106, 3.051346, 3.058741, 3.056497, 3.05877, 
    3.047397, 3.052265, 3.042275, 3.003668, 3.014965, 2.981394, 2.961385, 
    2.948162, 2.938815, 2.940135, 2.942652, 2.955621, 2.967863, 2.977226, 
    2.983505, 2.989704, 3.008549, 3.018567, 3.041116, 3.037033, 3.043952, 
    3.050575, 3.061726, 3.059888, 3.064811, 3.043768, 3.057738, 3.03471, 
    3.040992, 2.991397, 2.972703, 2.964797, 2.957888, 2.94115, 2.952699, 
    2.948141, 2.958995, 2.965913, 2.962489, 2.983677, 2.975423, 3.019161, 
    3.000246, 3.049801, 3.037871, 3.052668, 3.045108, 3.058072, 3.046402, 
    3.066645, 3.07107, 3.068045, 3.079679, 3.045757, 3.058742, 2.962394, 
    2.962952, 2.965553, 2.954137, 2.953439, 2.943016, 2.952289, 2.956246, 
    2.966314, 2.972286, 2.977973, 2.990513, 3.00458, 3.024358, 3.038643, 
    3.048256, 3.042357, 3.047564, 3.041744, 3.03902, 3.069412, 3.05231, 
    3.078004, 3.076576, 3.064928, 3.076737, 2.963344, 2.960133, 2.949014, 
    2.957712, 2.941883, 2.950734, 2.955835, 2.975596, 2.979954, 2.984001, 
    2.99201, 3.002319, 3.020487, 3.036381, 3.05096, 3.049889, 3.050266, 
    3.053532, 3.045449, 3.054861, 3.056444, 3.052308, 3.076385, 3.069487, 
    3.076546, 3.072053, 2.961176, 2.966582, 2.96366, 2.969157, 2.965284, 
    2.982547, 2.987741, 3.012164, 3.002116, 3.018121, 3.003737, 3.006282, 
    3.018646, 3.004513, 3.035503, 3.014461, 3.053659, 3.032526, 3.054989, 
    3.050897, 3.057674, 3.063756, 3.071424, 3.085462, 3.082273, 3.093804, 
    2.974658, 2.981702, 2.98108, 2.988467, 2.993942, 3.005841, 3.025021, 
    3.017794, 3.031074, 3.033747, 3.013577, 3.025946, 2.986425, 2.992777, 
    2.988993, 2.975213, 3.01946, 2.996674, 3.03888, 3.026438, 3.062889, 
    3.044709, 3.080518, 3.095463, 3.109589, 3.126186, 2.985552, 2.980758, 
    2.989347, 3.001271, 3.012373, 3.027195, 3.028715, 3.031502, 3.03873, 
    3.044821, 3.032384, 3.046349, 2.994254, 3.021445, 2.978949, 2.991685, 
    3.000566, 2.996666, 3.016969, 3.021774, 3.041377, 3.031227, 3.091769, 
    3.065044, 3.13888, 3.118208, 2.979085, 2.985535, 3.008091, 2.997339, 
    3.028187, 3.035828, 3.042052, 3.050029, 3.05089, 3.055627, 3.047869, 
    3.05532, 3.027227, 3.03975, 3.005504, 3.013805, 3.009983, 3.005797, 
    3.018735, 3.03258, 3.032875, 3.037328, 3.049915, 3.028312, 3.095174, 
    3.053899, 2.992584, 3.005078, 3.006864, 3.002016, 3.035061, 3.023047, 
    3.055511, 3.046704, 3.061147, 3.053962, 3.052906, 3.043704, 3.037989, 
    3.023597, 3.011936, 3.002719, 3.004859, 3.014992, 3.033429, 3.050969, 
    3.047119, 3.060047, 3.02594, 3.040197, 3.03468, 3.049087, 3.017603, 
    3.044399, 3.010791, 3.013723, 3.022809, 3.041168, 3.045242, 3.0496, 
    3.04691, 3.033898, 3.03177, 3.022588, 3.020058, 3.013084, 3.007323, 
    3.012587, 3.018125, 3.033902, 3.048191, 3.063843, 3.067685, 3.085922, 
    3.071104, 3.095401, 3.074809, 3.110406, 3.045956, 3.074187, 3.023223, 
    3.028673, 3.038557, 3.061342, 3.049019, 3.063435, 3.031687, 3.015344, 
    3.011127, 3.003278, 3.011307, 3.010653, 3.018353, 3.015876, 3.034428, 
    3.024449, 3.05288, 3.06332, 3.092594, 3.110337, 3.128503, 3.136558, 
    3.139013, 3.14004,
  2.969938, 2.988338, 2.98475, 2.999671, 2.991382, 3.001169, 2.973656, 
    2.989072, 2.979219, 2.971587, 3.028894, 3.000339, 3.058904, 3.040431, 
    3.087099, 3.056021, 3.093413, 3.086195, 3.107979, 3.101719, 3.129798, 
    3.110874, 3.144477, 3.125264, 3.128261, 3.110252, 3.006057, 3.025321, 
    3.004921, 3.007657, 3.006428, 2.991554, 2.984093, 2.968536, 2.971352, 
    2.982781, 3.008888, 2.999994, 3.022469, 3.021959, 3.047222, 3.0358, 
    3.078652, 3.066396, 3.101979, 3.092983, 3.101557, 3.098953, 3.10159, 
    3.088408, 3.094048, 3.082479, 3.037935, 3.050943, 3.01235, 2.989436, 
    2.97433, 2.963669, 2.965173, 2.968044, 2.982849, 2.996848, 3.007572, 
    3.014772, 3.021886, 3.043553, 3.055095, 3.081139, 3.076417, 3.084421, 
    3.092089, 3.10502, 3.102887, 3.108601, 3.084208, 3.100393, 3.073731, 
    3.080995, 3.02383, 3.00239, 2.993339, 2.985439, 2.966331, 2.979511, 
    2.974307, 2.986705, 2.994616, 2.9907, 3.014969, 3.005505, 3.055781, 
    3.033999, 3.091193, 3.077385, 3.094515, 3.085759, 3.100781, 3.087257, 
    3.11073, 3.115872, 3.112357, 3.125884, 3.086509, 3.101557, 2.99059, 
    2.991229, 2.994204, 2.981153, 2.980356, 2.968459, 2.979042, 2.983563, 
    2.995075, 3.001911, 3.008427, 3.022815, 3.038985, 3.061775, 3.078278, 
    3.089403, 3.082575, 3.088602, 3.081866, 3.078714, 3.113945, 3.094101, 
    3.123934, 3.122273, 3.108737, 3.12246, 2.991677, 2.988005, 2.975303, 
    2.985238, 2.967167, 2.977267, 2.983094, 3.005704, 3.010698, 3.015341, 
    3.024534, 3.036383, 3.057309, 3.075662, 3.092536, 3.091295, 3.091732, 
    3.095517, 3.086153, 3.097057, 3.098893, 3.094098, 3.122051, 3.114033, 
    3.122238, 3.117013, 2.989198, 2.995382, 2.992038, 2.998329, 2.993896, 
    3.013672, 3.019633, 3.047715, 3.03615, 3.054581, 3.038015, 3.040942, 
    3.055187, 3.038907, 3.074648, 3.050363, 3.095664, 3.071208, 3.097205, 
    3.092463, 3.100318, 3.107377, 3.116283, 3.132805, 3.128969, 3.142848, 
    3.004629, 3.012703, 3.01199, 3.020466, 3.026753, 3.040435, 3.062541, 
    3.054204, 3.069529, 3.072618, 3.049343, 3.063609, 3.018121, 3.025415, 
    3.021069, 3.005265, 3.056125, 3.029892, 3.078552, 3.064176, 3.106369, 
    3.085297, 3.12686, 3.144848, 3.161419, 3.180853, 3.01712, 3.011621, 
    3.021475, 3.035177, 3.047956, 3.065051, 3.066806, 3.070024, 3.078379, 
    3.085426, 3.071044, 3.087195, 3.027112, 3.058414, 3.009546, 3.024161, 
    3.034367, 3.029883, 3.053253, 3.058794, 3.08144, 3.069707, 3.140397, 
    3.108872, 3.195752, 3.171504, 3.009703, 3.017101, 3.043026, 3.030656, 
    3.066195, 3.075023, 3.082222, 3.091457, 3.092455, 3.097945, 3.088955, 
    3.097589, 3.065087, 3.079558, 3.040047, 3.049606, 3.045204, 3.040385, 
    3.055289, 3.07127, 3.07161, 3.076758, 3.091325, 3.06634, 3.1445, 
    3.095942, 3.025194, 3.039557, 3.041613, 3.036035, 3.074137, 3.060263, 
    3.097811, 3.087606, 3.104348, 3.096015, 3.094791, 3.084134, 3.077523, 
    3.060898, 3.047453, 3.036843, 3.039306, 3.050975, 3.07225, 3.092546, 
    3.088086, 3.103072, 3.063601, 3.080076, 3.073696, 3.090366, 3.053984, 
    3.084938, 3.046135, 3.049512, 3.059988, 3.081199, 3.085913, 3.090961, 
    3.087844, 3.072792, 3.070334, 3.059733, 3.056815, 3.048776, 3.042142, 
    3.048203, 3.054585, 3.072798, 3.089328, 3.107477, 3.111938, 3.133359, 
    3.115911, 3.144773, 3.120218, 3.162375, 3.08674, 3.119495, 3.060465, 
    3.066756, 3.078179, 3.104575, 3.090287, 3.107004, 3.070238, 3.05138, 
    3.046521, 3.037487, 3.046728, 3.045975, 3.054848, 3.051993, 3.073405, 
    3.06188, 3.094761, 3.106871, 3.141391, 3.162294, 3.18357, 3.193024, 
    3.195909, 3.197116,
  3.254741, 3.278218, 3.27363, 3.292737, 3.282113, 3.29466, 3.259476, 
    3.279157, 3.266568, 3.256841, 3.329907, 3.293594, 3.367681, 3.34439, 
    3.403476, 3.364038, 3.411533, 3.402324, 3.430179, 3.422155, 3.458265, 
    3.433895, 3.477267, 3.452414, 3.45628, 3.433097, 3.300939, 3.325432, 
    3.299479, 3.302996, 3.301417, 3.282333, 3.272791, 3.252957, 3.256542, 
    3.271116, 3.30458, 3.293151, 3.321862, 3.321224, 3.352938, 3.33857, 
    3.392721, 3.377164, 3.422489, 3.410983, 3.421947, 3.418616, 3.421991, 
    3.405146, 3.412344, 3.397591, 3.341253, 3.357629, 3.309036, 3.279623, 
    3.260335, 3.24677, 3.248682, 3.252332, 3.271201, 3.289116, 3.302887, 
    3.312155, 3.321133, 3.348318, 3.362868, 3.395885, 3.389879, 3.400063, 
    3.409842, 3.426385, 3.423651, 3.430977, 3.399792, 3.420458, 3.386468, 
    3.395701, 3.323565, 3.296227, 3.284619, 3.274511, 3.250153, 3.266941, 
    3.260305, 3.276129, 3.286255, 3.28124, 3.31241, 3.30023, 3.363734, 
    3.336309, 3.408699, 3.39111, 3.41294, 3.401767, 3.420955, 3.403677, 
    3.43371, 3.440318, 3.4358, 3.453213, 3.402724, 3.421948, 3.2811, 
    3.281917, 3.285727, 3.269036, 3.268019, 3.25286, 3.266342, 3.272114, 
    3.286843, 3.295613, 3.303987, 3.322295, 3.342572, 3.371312, 3.392245, 
    3.406414, 3.397712, 3.405393, 3.396809, 3.3928, 3.43784, 3.412412, 
    3.450698, 3.448558, 3.431152, 3.448799, 3.28249, 3.277792, 3.261575, 
    3.274255, 3.251216, 3.264078, 3.271514, 3.300485, 3.306909, 3.312889, 
    3.324445, 3.339303, 3.365666, 3.388921, 3.410413, 3.408829, 3.409386, 
    3.414221, 3.40227, 3.416191, 3.418538, 3.412408, 3.448272, 3.437953, 
    3.448513, 3.441786, 3.279318, 3.287236, 3.282954, 3.291016, 3.285333, 
    3.310739, 3.318315, 3.353559, 3.339009, 3.362219, 3.341353, 3.345033, 
    3.362985, 3.342474, 3.387632, 3.356896, 3.414409, 3.383265, 3.416379, 
    3.410319, 3.420363, 3.429406, 3.440847, 3.462151, 3.457195, 3.475155, 
    3.299103, 3.309491, 3.308573, 3.319357, 3.327225, 3.344395, 3.372282, 
    3.361744, 3.381135, 3.385054, 3.355611, 3.373633, 3.316427, 3.325549, 
    3.320111, 3.299921, 3.364169, 3.331158, 3.392593, 3.374351, 3.428114, 
    3.401179, 3.454473, 3.477749, 3.499924, 3.526197, 3.315176, 3.308097, 
    3.320619, 3.337789, 3.353863, 3.375459, 3.377682, 3.381763, 3.392373, 
    3.401343, 3.383056, 3.403599, 3.327674, 3.367062, 3.305427, 3.323979, 
    3.336771, 3.331147, 3.360543, 3.367542, 3.396268, 3.381361, 3.471978, 
    3.431325, 3.546064, 3.513538, 3.305628, 3.315152, 3.347654, 3.332116, 
    3.376909, 3.388108, 3.397263, 3.409035, 3.41031, 3.417326, 3.405843, 
    3.41687, 3.375505, 3.393873, 3.343907, 3.355943, 3.350395, 3.344331, 
    3.363113, 3.383343, 3.383775, 3.390312, 3.408867, 3.377093, 3.477297, 
    3.414765, 3.325272, 3.343291, 3.345876, 3.338865, 3.386982, 3.3694, 
    3.417154, 3.404122, 3.425524, 3.414857, 3.413294, 3.399697, 3.391284, 
    3.370203, 3.353229, 3.33988, 3.342975, 3.357669, 3.384588, 3.410426, 
    3.404735, 3.423888, 3.373624, 3.394532, 3.386423, 3.407643, 3.361465, 
    3.400721, 3.351568, 3.355824, 3.369052, 3.395961, 3.401964, 3.408402, 
    3.404426, 3.385276, 3.382156, 3.368729, 3.365041, 3.354896, 3.346541, 
    3.354174, 3.362225, 3.385283, 3.406319, 3.429536, 3.435262, 3.462867, 
    3.440368, 3.477652, 3.44591, 3.501212, 3.403018, 3.44498, 3.369656, 
    3.37762, 3.392119, 3.425814, 3.407542, 3.428928, 3.382034, 3.358179, 
    3.352055, 3.340689, 3.352316, 3.351367, 3.362557, 3.358953, 3.386053, 
    3.371446, 3.413255, 3.428757, 3.473265, 3.501104, 3.529883, 3.542462, 
    3.546271, 3.547866,
  3.812393, 3.852924, 3.844952, 3.878324, 3.859713, 3.881707, 3.820515, 
    3.854559, 3.83273, 3.815992, 3.945428, 3.879831, 4.016907, 3.972589, 
    4.084889, 4.009923, 4.100391, 4.082681, 4.136661, 4.120984, 4.192374, 
    4.143956, 4.230835, 4.180657, 4.188393, 4.142387, 3.892786, 3.937096, 
    3.890205, 3.896428, 3.893631, 3.860096, 3.843497, 3.80934, 3.815479, 
    3.840594, 3.899235, 3.879052, 3.93047, 3.929288, 3.988761, 3.961638, 
    4.064354, 4.034963, 4.121634, 4.099329, 4.12058, 4.114101, 4.120664, 
    4.088093, 4.101956, 4.073629, 3.96668, 3.997681, 3.907147, 3.855371, 
    3.821992, 3.798779, 3.802038, 3.808271, 3.840742, 3.871965, 3.896233, 
    3.912702, 3.929118, 3.980006, 4.007683, 4.070376, 4.058958, 4.078353, 
    4.097129, 4.129234, 4.123899, 4.138225, 4.077835, 4.117682, 4.052496, 
    4.070027, 3.93363, 3.884468, 3.86409, 3.846481, 3.804549, 3.833373, 
    3.82194, 3.849291, 3.866952, 3.858189, 3.913155, 3.891532, 4.00934, 
    3.957397, 4.094926, 4.061294, 4.103108, 4.081614, 4.118647, 4.085275, 
    4.143593, 4.15662, 4.147705, 4.182254, 4.083448, 4.120581, 3.857945, 
    3.85937, 3.866028, 3.836994, 3.835237, 3.809173, 3.832339, 3.842323, 
    3.867982, 3.883384, 3.898182, 3.931272, 3.969163, 4.023889, 4.06345, 
    4.09053, 4.073862, 4.088568, 4.072139, 4.064504, 4.151726, 4.102087, 
    4.177233, 4.172968, 4.138568, 4.173448, 3.860372, 3.852184, 3.824124, 
    3.846036, 3.806363, 3.828434, 3.841284, 3.891984, 3.903368, 3.91401, 
    3.935263, 3.963014, 4.01304, 4.05714, 4.098228, 4.095177, 4.096251, 
    4.105585, 4.082578, 4.109398, 4.113951, 4.102079, 4.172398, 4.151948, 
    4.172878, 4.159524, 3.85484, 3.86867, 3.86118, 3.875299, 3.865339, 
    3.910178, 3.923903, 3.989941, 3.962463, 4.006441, 3.966868, 3.973802, 
    4.007906, 3.968978, 4.0547, 3.996286, 4.105948, 4.046445, 4.109763, 
    4.098048, 4.117496, 4.135146, 4.157666, 4.200188, 4.190227, 4.226529, 
    3.889542, 3.907957, 3.906323, 3.92583, 3.940431, 3.972598, 4.025756, 
    4.005533, 4.042431, 4.049824, 3.99384, 4.028343, 3.920414, 3.937314, 
    3.927225, 3.890987, 4.010172, 3.947763, 4.064112, 4.029688, 4.132617, 
    4.080488, 4.184773, 4.231818, 4.277538, 4.332246, 3.918106, 3.905478, 
    3.928167, 3.960172, 3.990517, 4.031764, 4.035937, 4.043613, 4.063693, 
    4.080802, 4.046052, 4.085124, 3.941268, 4.015719, 3.900735, 3.934397, 
    3.958264, 3.947742, 4.003239, 4.01664, 4.071107, 4.042855, 4.220065, 
    4.138907, 4.374605, 4.306057, 3.901093, 3.918061, 3.978752, 3.949552, 
    4.034485, 4.055602, 4.073004, 4.095573, 4.09803, 4.111598, 4.089432, 
    4.110715, 4.031851, 4.066545, 3.971679, 3.994471, 3.98394, 3.972478, 
    4.008152, 4.046594, 4.047409, 4.05978, 4.09525, 4.03483, 4.230896, 
    4.106637, 3.936798, 3.970517, 3.975394, 3.962193, 4.053471, 4.020208, 
    4.111266, 4.086128, 4.127552, 4.106816, 4.103791, 4.077653, 4.061625, 
    4.021753, 3.989313, 3.964099, 3.969922, 3.997757, 4.048943, 4.098255, 
    4.087304, 4.124361, 4.028325, 4.0678, 4.052412, 4.092893, 4.005001, 
    4.079612, 3.986161, 3.994245, 4.019541, 4.070521, 4.081992, 4.094354, 
    4.086712, 4.050242, 4.044355, 4.018919, 4.011842, 3.992481, 3.976649, 
    3.991108, 4.006452, 4.050256, 4.090347, 4.1354, 4.146646, 4.201631, 
    4.156718, 4.231621, 4.167703, 4.280221, 4.084012, 4.165855, 4.020701, 
    4.03582, 4.06321, 4.128119, 4.0927, 4.134209, 4.044125, 3.99873, 
    3.987085, 3.965621, 3.98758, 3.985781, 4.007088, 4.000206, 4.051713, 
    4.024146, 4.103716, 4.133875, 4.222682, 4.279996, 4.339895, 4.366773, 
    4.375056, 4.378533,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24813.87, 24834.3, 24830.29, 24847.02, 24837.71, 24848.71, 24817.97, 
    24835.12, 24824.14, 24815.69, 24880.24, 24847.78, 24915.03, 24893.52, 
    24948.02, 24911.65, 24955.49, 24946.95, 24972.88, 24965.38, 24999.34, 
    24976.36, 25017.42, 24993.8, 24997.46, 24975.61, 24854.24, 24876.15, 
    24852.95, 24856.05, 24854.66, 24837.9, 24829.56, 24812.32, 24815.43, 
    24828.1, 24857.45, 24847.39, 24872.9, 24872.32, 24901.39, 24888.17, 
    24938.08, 24923.79, 24965.69, 24954.98, 24965.18, 24962.08, 24965.22, 
    24949.57, 24956.24, 24942.57, 24890.63, 24905.72, 24861.38, 24835.53, 
    24818.72, 24806.96, 24808.62, 24811.78, 24828.18, 24843.84, 24855.96, 
    24864.14, 24872.24, 24897.13, 24910.57, 24941, 24935.46, 24944.86, 
    24953.92, 24969.32, 24966.77, 24973.62, 24944.61, 24963.79, 24932.32, 
    24940.83, 24874.45, 24850.09, 24839.9, 24831.06, 24809.89, 24824.46, 
    24818.69, 24832.48, 24841.33, 24836.94, 24864.36, 24853.61, 24911.37, 
    24886.1, 24952.86, 24936.6, 24956.8, 24946.44, 24964.26, 24948.21, 
    24976.18, 24982.39, 24978.14, 24994.56, 24947.32, 24965.18, 24836.82, 
    24837.54, 24840.87, 24826.29, 24825.4, 24812.24, 24823.94, 24828.97, 
    24841.85, 24849.55, 24856.92, 24873.29, 24891.85, 24918.4, 24937.64, 
    24950.74, 24942.69, 24949.8, 24941.85, 24938.15, 24980.06, 24956.31, 
    24992.18, 24990.16, 24973.79, 24990.38, 24838.04, 24833.93, 24819.8, 
    24830.84, 24810.81, 24821.97, 24828.45, 24853.84, 24859.5, 24864.79, 
    24875.26, 24888.84, 24913.16, 24934.58, 24954.45, 24952.98, 24953.5, 
    24957.99, 24946.9, 24959.82, 24962, 24956.3, 24989.88, 24980.17, 
    24990.11, 24983.77, 24835.26, 24842.2, 24838.44, 24845.51, 24840.53, 
    24862.89, 24869.67, 24901.96, 24888.58, 24909.96, 24890.73, 24894.11, 
    24910.67, 24891.76, 24933.39, 24905.04, 24958.16, 24929.38, 24959.99, 
    24954.36, 24963.7, 24972.15, 24982.89, 25003.02, 24998.32, 25015.4, 
    24852.62, 24861.78, 24860.97, 24870.62, 24877.79, 24893.52, 24919.3, 
    24909.53, 24927.43, 24931.02, 24903.85, 24920.55, 24867.96, 24876.26, 
    24871.31, 24853.34, 24911.77, 24881.38, 24937.96, 24921.21, 24970.94, 
    24945.89, 24995.75, 25017.88, 25039.16, 25064.5, 24866.82, 24860.55, 
    24871.77, 24887.46, 24902.24, 24922.22, 24924.26, 24928, 24937.76, 
    24946.04, 24929.19, 24948.13, 24878.2, 24914.45, 24858.2, 24874.83, 
    24886.52, 24881.38, 24908.41, 24914.9, 24941.35, 24927.63, 25012.37, 
    24973.95, 25084.01, 25052.34, 24858.37, 24866.79, 24896.52, 24882.26, 
    24923.55, 24933.83, 24942.27, 24953.17, 24954.35, 24960.88, 24950.21, 
    24960.45, 24922.27, 24939.14, 24893.07, 24904.16, 24899.04, 24893.46, 
    24910.79, 24929.45, 24929.85, 24935.86, 24953.02, 24923.72, 25017.45, 
    24958.49, 24876.01, 24892.51, 24894.88, 24888.44, 24932.8, 24916.62, 
    24960.71, 24948.62, 24968.52, 24958.58, 24957.12, 24944.52, 24936.76, 
    24917.37, 24901.66, 24889.38, 24892.22, 24905.76, 24930.6, 24954.46, 
    24949.19, 24966.99, 24920.54, 24939.75, 24932.28, 24951.88, 24909.27, 
    24945.47, 24900.12, 24904.05, 24916.3, 24941.07, 24946.62, 24952.58, 
    24948.9, 24931.23, 24928.36, 24916, 24912.58, 24903.19, 24895.49, 
    24902.53, 24909.97, 24931.23, 24950.65, 24972.27, 24977.64, 25003.7, 
    24982.44, 25017.79, 24987.66, 25040.41, 24947.6, 24986.78, 24916.86, 
    24924.2, 24937.53, 24968.79, 24951.79, 24971.7, 24928.25, 24906.23, 
    24900.57, 24890.12, 24900.81, 24899.94, 24910.28, 24906.94, 24931.94, 
    24918.53, 24957.09, 24971.54, 25013.6, 25040.3, 25068.05, 25080.42, 
    25084.22, 25085.81 ;

 HCSOI =
  24813.87, 24834.3, 24830.29, 24847.02, 24837.71, 24848.71, 24817.97, 
    24835.12, 24824.14, 24815.69, 24880.24, 24847.78, 24915.03, 24893.52, 
    24948.02, 24911.65, 24955.49, 24946.95, 24972.88, 24965.38, 24999.34, 
    24976.36, 25017.42, 24993.8, 24997.46, 24975.61, 24854.24, 24876.15, 
    24852.95, 24856.05, 24854.66, 24837.9, 24829.56, 24812.32, 24815.43, 
    24828.1, 24857.45, 24847.39, 24872.9, 24872.32, 24901.39, 24888.17, 
    24938.08, 24923.79, 24965.69, 24954.98, 24965.18, 24962.08, 24965.22, 
    24949.57, 24956.24, 24942.57, 24890.63, 24905.72, 24861.38, 24835.53, 
    24818.72, 24806.96, 24808.62, 24811.78, 24828.18, 24843.84, 24855.96, 
    24864.14, 24872.24, 24897.13, 24910.57, 24941, 24935.46, 24944.86, 
    24953.92, 24969.32, 24966.77, 24973.62, 24944.61, 24963.79, 24932.32, 
    24940.83, 24874.45, 24850.09, 24839.9, 24831.06, 24809.89, 24824.46, 
    24818.69, 24832.48, 24841.33, 24836.94, 24864.36, 24853.61, 24911.37, 
    24886.1, 24952.86, 24936.6, 24956.8, 24946.44, 24964.26, 24948.21, 
    24976.18, 24982.39, 24978.14, 24994.56, 24947.32, 24965.18, 24836.82, 
    24837.54, 24840.87, 24826.29, 24825.4, 24812.24, 24823.94, 24828.97, 
    24841.85, 24849.55, 24856.92, 24873.29, 24891.85, 24918.4, 24937.64, 
    24950.74, 24942.69, 24949.8, 24941.85, 24938.15, 24980.06, 24956.31, 
    24992.18, 24990.16, 24973.79, 24990.38, 24838.04, 24833.93, 24819.8, 
    24830.84, 24810.81, 24821.97, 24828.45, 24853.84, 24859.5, 24864.79, 
    24875.26, 24888.84, 24913.16, 24934.58, 24954.45, 24952.98, 24953.5, 
    24957.99, 24946.9, 24959.82, 24962, 24956.3, 24989.88, 24980.17, 
    24990.11, 24983.77, 24835.26, 24842.2, 24838.44, 24845.51, 24840.53, 
    24862.89, 24869.67, 24901.96, 24888.58, 24909.96, 24890.73, 24894.11, 
    24910.67, 24891.76, 24933.39, 24905.04, 24958.16, 24929.38, 24959.99, 
    24954.36, 24963.7, 24972.15, 24982.89, 25003.02, 24998.32, 25015.4, 
    24852.62, 24861.78, 24860.97, 24870.62, 24877.79, 24893.52, 24919.3, 
    24909.53, 24927.43, 24931.02, 24903.85, 24920.55, 24867.96, 24876.26, 
    24871.31, 24853.34, 24911.77, 24881.38, 24937.96, 24921.21, 24970.94, 
    24945.89, 24995.75, 25017.88, 25039.16, 25064.5, 24866.82, 24860.55, 
    24871.77, 24887.46, 24902.24, 24922.22, 24924.26, 24928, 24937.76, 
    24946.04, 24929.19, 24948.13, 24878.2, 24914.45, 24858.2, 24874.83, 
    24886.52, 24881.38, 24908.41, 24914.9, 24941.35, 24927.63, 25012.37, 
    24973.95, 25084.01, 25052.34, 24858.37, 24866.79, 24896.52, 24882.26, 
    24923.55, 24933.83, 24942.27, 24953.17, 24954.35, 24960.88, 24950.21, 
    24960.45, 24922.27, 24939.14, 24893.07, 24904.16, 24899.04, 24893.46, 
    24910.79, 24929.45, 24929.85, 24935.86, 24953.02, 24923.72, 25017.45, 
    24958.49, 24876.01, 24892.51, 24894.88, 24888.44, 24932.8, 24916.62, 
    24960.71, 24948.62, 24968.52, 24958.58, 24957.12, 24944.52, 24936.76, 
    24917.37, 24901.66, 24889.38, 24892.22, 24905.76, 24930.6, 24954.46, 
    24949.19, 24966.99, 24920.54, 24939.75, 24932.28, 24951.88, 24909.27, 
    24945.47, 24900.12, 24904.05, 24916.3, 24941.07, 24946.62, 24952.58, 
    24948.9, 24931.23, 24928.36, 24916, 24912.58, 24903.19, 24895.49, 
    24902.53, 24909.97, 24931.23, 24950.65, 24972.27, 24977.64, 25003.7, 
    24982.44, 25017.79, 24987.66, 25040.41, 24947.6, 24986.78, 24916.86, 
    24924.2, 24937.53, 24968.79, 24951.79, 24971.7, 24928.25, 24906.23, 
    24900.57, 24890.12, 24900.81, 24899.94, 24910.28, 24906.94, 24931.94, 
    24918.53, 24957.09, 24971.54, 25013.6, 25040.3, 25068.05, 25080.42, 
    25084.22, 25085.81 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371698e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441075e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379093e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377207e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523353e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.56315e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529406e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.532169e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547246e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.46224e-08, 6.465288e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532766e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472856e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 HR_vr =
  2.669659e-07, 2.676731e-07, 2.675357e-07, 2.681056e-07, 2.677895e-07, 
    2.681626e-07, 2.671093e-07, 2.677012e-07, 2.673234e-07, 2.670296e-07, 
    2.692103e-07, 2.68131e-07, 2.703289e-07, 2.696422e-07, 2.713656e-07, 
    2.702221e-07, 2.715959e-07, 2.713326e-07, 2.721245e-07, 2.718978e-07, 
    2.729097e-07, 2.722292e-07, 2.734334e-07, 2.727472e-07, 2.728546e-07, 
    2.722067e-07, 2.683483e-07, 2.69076e-07, 2.683052e-07, 2.68409e-07, 
    2.683624e-07, 2.677961e-07, 2.675105e-07, 2.669118e-07, 2.670205e-07, 
    2.674602e-07, 2.684557e-07, 2.681179e-07, 2.689687e-07, 2.689495e-07, 
    2.698954e-07, 2.694691e-07, 2.710565e-07, 2.706058e-07, 2.719072e-07, 
    2.715802e-07, 2.718919e-07, 2.717974e-07, 2.718931e-07, 2.714134e-07, 
    2.71619e-07, 2.711967e-07, 2.69549e-07, 2.700337e-07, 2.685868e-07, 
    2.677151e-07, 2.671353e-07, 2.667236e-07, 2.667818e-07, 2.668928e-07, 
    2.674628e-07, 2.679981e-07, 2.684058e-07, 2.686783e-07, 2.689468e-07, 
    2.697587e-07, 2.701878e-07, 2.711476e-07, 2.709744e-07, 2.712677e-07, 
    2.715476e-07, 2.720174e-07, 2.719401e-07, 2.72147e-07, 2.712599e-07, 
    2.718496e-07, 2.708759e-07, 2.711423e-07, 2.690199e-07, 2.68209e-07, 
    2.678642e-07, 2.675621e-07, 2.668266e-07, 2.673346e-07, 2.671344e-07, 
    2.676106e-07, 2.67913e-07, 2.677634e-07, 2.686858e-07, 2.683274e-07, 
    2.702132e-07, 2.694017e-07, 2.71515e-07, 2.7101e-07, 2.71636e-07, 
    2.713166e-07, 2.718637e-07, 2.713713e-07, 2.72224e-07, 2.724095e-07, 
    2.722827e-07, 2.727694e-07, 2.71344e-07, 2.718919e-07, 2.677592e-07, 
    2.677836e-07, 2.678973e-07, 2.673977e-07, 2.673671e-07, 2.669088e-07, 
    2.673166e-07, 2.674902e-07, 2.679305e-07, 2.681908e-07, 2.684382e-07, 
    2.689818e-07, 2.695882e-07, 2.704351e-07, 2.710427e-07, 2.714497e-07, 
    2.712002e-07, 2.714205e-07, 2.711742e-07, 2.710587e-07, 2.7234e-07, 
    2.716209e-07, 2.726995e-07, 2.726398e-07, 2.721519e-07, 2.726465e-07, 
    2.678008e-07, 2.676604e-07, 2.671728e-07, 2.675544e-07, 2.668589e-07, 
    2.672483e-07, 2.674722e-07, 2.683349e-07, 2.685242e-07, 2.686998e-07, 
    2.690464e-07, 2.694909e-07, 2.702699e-07, 2.709467e-07, 2.715639e-07, 
    2.715187e-07, 2.715346e-07, 2.716724e-07, 2.71331e-07, 2.717285e-07, 
    2.717952e-07, 2.716208e-07, 2.726318e-07, 2.723432e-07, 2.726385e-07, 
    2.724506e-07, 2.67706e-07, 2.679422e-07, 2.678146e-07, 2.680545e-07, 
    2.678855e-07, 2.686368e-07, 2.688618e-07, 2.699137e-07, 2.694822e-07, 
    2.701688e-07, 2.695519e-07, 2.696613e-07, 2.701912e-07, 2.695853e-07, 
    2.709095e-07, 2.700121e-07, 2.716778e-07, 2.70783e-07, 2.717338e-07, 
    2.715612e-07, 2.718469e-07, 2.721027e-07, 2.724243e-07, 2.730173e-07, 
    2.7288e-07, 2.733755e-07, 2.682941e-07, 2.686001e-07, 2.685732e-07, 
    2.688932e-07, 2.691299e-07, 2.696424e-07, 2.704634e-07, 2.701548e-07, 
    2.707212e-07, 2.708349e-07, 2.699743e-07, 2.705029e-07, 2.688049e-07, 
    2.690795e-07, 2.68916e-07, 2.683183e-07, 2.70226e-07, 2.692477e-07, 
    2.710528e-07, 2.705238e-07, 2.720663e-07, 2.712997e-07, 2.728044e-07, 
    2.734466e-07, 2.740501e-07, 2.747547e-07, 2.687671e-07, 2.685592e-07, 
    2.689313e-07, 2.694458e-07, 2.699227e-07, 2.705561e-07, 2.706209e-07, 
    2.707395e-07, 2.710464e-07, 2.713044e-07, 2.70777e-07, 2.713691e-07, 
    2.691433e-07, 2.703108e-07, 2.684806e-07, 2.690324e-07, 2.694155e-07, 
    2.692474e-07, 2.701195e-07, 2.703249e-07, 2.711586e-07, 2.707278e-07, 
    2.732882e-07, 2.721568e-07, 2.752905e-07, 2.744165e-07, 2.684866e-07, 
    2.687663e-07, 2.69739e-07, 2.692764e-07, 2.705983e-07, 2.709232e-07, 
    2.711872e-07, 2.715246e-07, 2.71561e-07, 2.717607e-07, 2.714334e-07, 
    2.717478e-07, 2.705575e-07, 2.710896e-07, 2.696279e-07, 2.69984e-07, 
    2.698202e-07, 2.696405e-07, 2.70195e-07, 2.707853e-07, 2.707978e-07, 
    2.709869e-07, 2.715198e-07, 2.706037e-07, 2.734342e-07, 2.716879e-07, 
    2.690713e-07, 2.696096e-07, 2.696863e-07, 2.694779e-07, 2.708908e-07, 
    2.703792e-07, 2.717559e-07, 2.713841e-07, 2.719931e-07, 2.716906e-07, 
    2.71646e-07, 2.712572e-07, 2.71015e-07, 2.704027e-07, 2.699039e-07, 
    2.695081e-07, 2.696002e-07, 2.700349e-07, 2.708214e-07, 2.715643e-07, 
    2.714016e-07, 2.719468e-07, 2.705026e-07, 2.711086e-07, 2.708745e-07, 
    2.714848e-07, 2.701466e-07, 2.712866e-07, 2.698549e-07, 2.699805e-07, 
    2.70369e-07, 2.711498e-07, 2.713223e-07, 2.715065e-07, 2.713928e-07, 
    2.708413e-07, 2.707509e-07, 2.703596e-07, 2.702515e-07, 2.699532e-07, 
    2.69706e-07, 2.699319e-07, 2.701689e-07, 2.708415e-07, 2.71447e-07, 
    2.721064e-07, 2.722676e-07, 2.73037e-07, 2.724109e-07, 2.734439e-07, 
    2.725658e-07, 2.740848e-07, 2.713524e-07, 2.725399e-07, 2.703867e-07, 
    2.706191e-07, 2.710391e-07, 2.720013e-07, 2.71482e-07, 2.720892e-07, 
    2.707473e-07, 2.700499e-07, 2.698693e-07, 2.695322e-07, 2.69877e-07, 
    2.69849e-07, 2.701787e-07, 2.700727e-07, 2.708638e-07, 2.70439e-07, 
    2.716449e-07, 2.720844e-07, 2.733236e-07, 2.740819e-07, 2.748527e-07, 
    2.751926e-07, 2.752961e-07, 2.753393e-07,
  2.414858e-07, 2.423968e-07, 2.422197e-07, 2.42954e-07, 2.425468e-07, 
    2.430274e-07, 2.416706e-07, 2.424329e-07, 2.419463e-07, 2.415678e-07, 
    2.443772e-07, 2.429867e-07, 2.458195e-07, 2.449343e-07, 2.471562e-07, 
    2.456817e-07, 2.474533e-07, 2.471138e-07, 2.481353e-07, 2.478427e-07, 
    2.491479e-07, 2.482702e-07, 2.498238e-07, 2.489384e-07, 2.49077e-07, 
    2.482413e-07, 2.432668e-07, 2.442042e-07, 2.432112e-07, 2.433449e-07, 
    2.432849e-07, 2.425552e-07, 2.421872e-07, 2.414161e-07, 2.415562e-07, 
    2.421225e-07, 2.434051e-07, 2.429699e-07, 2.440663e-07, 2.440416e-07, 
    2.452606e-07, 2.447112e-07, 2.467577e-07, 2.461765e-07, 2.47855e-07, 
    2.474331e-07, 2.478351e-07, 2.477133e-07, 2.478367e-07, 2.47218e-07, 
    2.474831e-07, 2.469385e-07, 2.448141e-07, 2.45439e-07, 2.43574e-07, 
    2.424507e-07, 2.41704e-07, 2.411737e-07, 2.412487e-07, 2.413916e-07, 
    2.421258e-07, 2.428156e-07, 2.433408e-07, 2.436921e-07, 2.44038e-07, 
    2.450842e-07, 2.456375e-07, 2.468751e-07, 2.46652e-07, 2.4703e-07, 
    2.473912e-07, 2.479971e-07, 2.478974e-07, 2.481642e-07, 2.470201e-07, 
    2.477806e-07, 2.465248e-07, 2.468684e-07, 2.441319e-07, 2.430873e-07, 
    2.426429e-07, 2.422538e-07, 2.413063e-07, 2.419607e-07, 2.417028e-07, 
    2.423163e-07, 2.427059e-07, 2.425132e-07, 2.437017e-07, 2.432398e-07, 
    2.456703e-07, 2.446242e-07, 2.47349e-07, 2.466978e-07, 2.475051e-07, 
    2.470932e-07, 2.477988e-07, 2.471638e-07, 2.482635e-07, 2.485028e-07, 
    2.483393e-07, 2.489672e-07, 2.471286e-07, 2.478351e-07, 2.425078e-07, 
    2.425392e-07, 2.426856e-07, 2.420419e-07, 2.420026e-07, 2.414123e-07, 
    2.419375e-07, 2.421611e-07, 2.427284e-07, 2.430639e-07, 2.433826e-07, 
    2.44083e-07, 2.448646e-07, 2.459564e-07, 2.4674e-07, 2.472649e-07, 
    2.469431e-07, 2.472272e-07, 2.469096e-07, 2.467607e-07, 2.484131e-07, 
    2.474856e-07, 2.488769e-07, 2.488e-07, 2.481706e-07, 2.488086e-07, 
    2.425613e-07, 2.423805e-07, 2.417523e-07, 2.422439e-07, 2.41348e-07, 
    2.418496e-07, 2.421378e-07, 2.432494e-07, 2.434935e-07, 2.437197e-07, 
    2.441664e-07, 2.447393e-07, 2.457434e-07, 2.466162e-07, 2.474122e-07, 
    2.473539e-07, 2.473744e-07, 2.475521e-07, 2.471118e-07, 2.476244e-07, 
    2.477104e-07, 2.474855e-07, 2.487897e-07, 2.484173e-07, 2.487983e-07, 
    2.485559e-07, 2.424393e-07, 2.427435e-07, 2.425791e-07, 2.428882e-07, 
    2.426704e-07, 2.436384e-07, 2.439284e-07, 2.452842e-07, 2.44728e-07, 
    2.45613e-07, 2.44818e-07, 2.449589e-07, 2.456418e-07, 2.44861e-07, 
    2.46568e-07, 2.45411e-07, 2.47559e-07, 2.464049e-07, 2.476313e-07, 
    2.474087e-07, 2.477772e-07, 2.481071e-07, 2.48522e-07, 2.492869e-07, 
    2.491098e-07, 2.497491e-07, 2.431969e-07, 2.435912e-07, 2.435565e-07, 
    2.43969e-07, 2.442739e-07, 2.449345e-07, 2.45993e-07, 2.455951e-07, 
    2.463254e-07, 2.46472e-07, 2.453624e-07, 2.460438e-07, 2.43855e-07, 
    2.44209e-07, 2.439983e-07, 2.43228e-07, 2.456868e-07, 2.444258e-07, 
    2.467529e-07, 2.460709e-07, 2.480601e-07, 2.470713e-07, 2.490123e-07, 
    2.498407e-07, 2.506197e-07, 2.51529e-07, 2.438064e-07, 2.435385e-07, 
    2.440181e-07, 2.44681e-07, 2.452958e-07, 2.461125e-07, 2.46196e-07, 
    2.463489e-07, 2.467448e-07, 2.470775e-07, 2.463972e-07, 2.471609e-07, 
    2.44291e-07, 2.457962e-07, 2.434372e-07, 2.441482e-07, 2.44642e-07, 
    2.444254e-07, 2.455496e-07, 2.458144e-07, 2.468894e-07, 2.463339e-07, 
    2.496363e-07, 2.481767e-07, 2.522208e-07, 2.510926e-07, 2.434449e-07, 
    2.438055e-07, 2.450591e-07, 2.444628e-07, 2.46167e-07, 2.465859e-07, 
    2.469264e-07, 2.473614e-07, 2.474084e-07, 2.47666e-07, 2.472438e-07, 
    2.476493e-07, 2.461142e-07, 2.468005e-07, 2.449159e-07, 2.453749e-07, 
    2.451638e-07, 2.449321e-07, 2.45647e-07, 2.464079e-07, 2.464242e-07, 
    2.46668e-07, 2.473548e-07, 2.461739e-07, 2.498244e-07, 2.475716e-07, 
    2.441984e-07, 2.448921e-07, 2.449912e-07, 2.447225e-07, 2.46544e-07, 
    2.458844e-07, 2.476597e-07, 2.471803e-07, 2.479657e-07, 2.475755e-07, 
    2.475181e-07, 2.470166e-07, 2.467042e-07, 2.459147e-07, 2.452717e-07, 
    2.447615e-07, 2.448802e-07, 2.454405e-07, 2.464544e-07, 2.474126e-07, 
    2.472028e-07, 2.47906e-07, 2.460435e-07, 2.46825e-07, 2.46523e-07, 
    2.473101e-07, 2.455845e-07, 2.470541e-07, 2.452085e-07, 2.453705e-07, 
    2.458713e-07, 2.468779e-07, 2.471005e-07, 2.473381e-07, 2.471915e-07, 
    2.464802e-07, 2.463636e-07, 2.458592e-07, 2.457198e-07, 2.453352e-07, 
    2.450167e-07, 2.453077e-07, 2.456133e-07, 2.464805e-07, 2.472613e-07, 
    2.481118e-07, 2.483198e-07, 2.493122e-07, 2.485044e-07, 2.49837e-07, 
    2.487041e-07, 2.506642e-07, 2.471392e-07, 2.486708e-07, 2.458941e-07, 
    2.461937e-07, 2.467352e-07, 2.479761e-07, 2.473064e-07, 2.480896e-07, 
    2.46359e-07, 2.454598e-07, 2.45227e-07, 2.447925e-07, 2.45237e-07, 
    2.452008e-07, 2.456259e-07, 2.454893e-07, 2.465093e-07, 2.459616e-07, 
    2.475166e-07, 2.480834e-07, 2.496821e-07, 2.506607e-07, 2.516557e-07, 
    2.520946e-07, 2.522281e-07, 2.522839e-07,
  2.259477e-07, 2.26945e-07, 2.267512e-07, 2.275552e-07, 2.271093e-07, 
    2.276357e-07, 2.2615e-07, 2.269846e-07, 2.264519e-07, 2.260375e-07, 
    2.291142e-07, 2.275911e-07, 2.306949e-07, 2.297247e-07, 2.321607e-07, 
    2.305439e-07, 2.324865e-07, 2.321141e-07, 2.332346e-07, 2.329137e-07, 
    2.343459e-07, 2.333827e-07, 2.350877e-07, 2.341159e-07, 2.34268e-07, 
    2.333509e-07, 2.278978e-07, 2.289247e-07, 2.278369e-07, 2.279834e-07, 
    2.279177e-07, 2.271185e-07, 2.267156e-07, 2.258715e-07, 2.260248e-07, 
    2.266447e-07, 2.280493e-07, 2.275727e-07, 2.287736e-07, 2.287465e-07, 
    2.300823e-07, 2.294802e-07, 2.317236e-07, 2.310863e-07, 2.329271e-07, 
    2.324644e-07, 2.329054e-07, 2.327717e-07, 2.329071e-07, 2.322284e-07, 
    2.325192e-07, 2.319219e-07, 2.29593e-07, 2.302778e-07, 2.282343e-07, 
    2.270041e-07, 2.261866e-07, 2.256062e-07, 2.256882e-07, 2.258447e-07, 
    2.266484e-07, 2.274036e-07, 2.279789e-07, 2.283636e-07, 2.287426e-07, 
    2.29889e-07, 2.304954e-07, 2.318524e-07, 2.316076e-07, 2.320223e-07, 
    2.324183e-07, 2.33083e-07, 2.329736e-07, 2.332664e-07, 2.320114e-07, 
    2.328456e-07, 2.314682e-07, 2.31845e-07, 2.288455e-07, 2.277012e-07, 
    2.272145e-07, 2.267885e-07, 2.257513e-07, 2.264676e-07, 2.261853e-07, 
    2.268569e-07, 2.272835e-07, 2.270725e-07, 2.283741e-07, 2.278683e-07, 
    2.305314e-07, 2.293849e-07, 2.323722e-07, 2.316579e-07, 2.325433e-07, 
    2.320916e-07, 2.328655e-07, 2.32169e-07, 2.333753e-07, 2.336378e-07, 
    2.334585e-07, 2.341475e-07, 2.321304e-07, 2.329054e-07, 2.270666e-07, 
    2.27101e-07, 2.272614e-07, 2.265566e-07, 2.265134e-07, 2.258673e-07, 
    2.264423e-07, 2.26687e-07, 2.273082e-07, 2.276756e-07, 2.280247e-07, 
    2.287919e-07, 2.296483e-07, 2.30845e-07, 2.317042e-07, 2.322798e-07, 
    2.319269e-07, 2.322385e-07, 2.318902e-07, 2.317269e-07, 2.335395e-07, 
    2.325219e-07, 2.340484e-07, 2.33964e-07, 2.332733e-07, 2.339735e-07, 
    2.271252e-07, 2.269272e-07, 2.262394e-07, 2.267777e-07, 2.257969e-07, 
    2.26346e-07, 2.266616e-07, 2.278788e-07, 2.281461e-07, 2.283939e-07, 
    2.288833e-07, 2.29511e-07, 2.306115e-07, 2.315684e-07, 2.324414e-07, 
    2.323774e-07, 2.324e-07, 2.325949e-07, 2.32112e-07, 2.326742e-07, 
    2.327685e-07, 2.325218e-07, 2.339527e-07, 2.335441e-07, 2.339622e-07, 
    2.336962e-07, 2.269916e-07, 2.273247e-07, 2.271447e-07, 2.274832e-07, 
    2.272447e-07, 2.283048e-07, 2.286225e-07, 2.301081e-07, 2.294986e-07, 
    2.304686e-07, 2.295972e-07, 2.297516e-07, 2.305001e-07, 2.296443e-07, 
    2.315156e-07, 2.302472e-07, 2.326025e-07, 2.313367e-07, 2.326818e-07, 
    2.324376e-07, 2.328418e-07, 2.332037e-07, 2.336589e-07, 2.344984e-07, 
    2.34304e-07, 2.350058e-07, 2.278213e-07, 2.282532e-07, 2.282152e-07, 
    2.28667e-07, 2.290011e-07, 2.297249e-07, 2.308851e-07, 2.30449e-07, 
    2.312496e-07, 2.314103e-07, 2.301939e-07, 2.309408e-07, 2.285421e-07, 
    2.289299e-07, 2.286991e-07, 2.278554e-07, 2.305494e-07, 2.291674e-07, 
    2.317184e-07, 2.309705e-07, 2.331521e-07, 2.320675e-07, 2.34197e-07, 
    2.351063e-07, 2.359616e-07, 2.369604e-07, 2.284888e-07, 2.281954e-07, 
    2.287208e-07, 2.294472e-07, 2.301209e-07, 2.310161e-07, 2.311077e-07, 
    2.312753e-07, 2.317094e-07, 2.320744e-07, 2.313283e-07, 2.321658e-07, 
    2.290198e-07, 2.306694e-07, 2.280845e-07, 2.288633e-07, 2.294044e-07, 
    2.291671e-07, 2.303991e-07, 2.306893e-07, 2.31868e-07, 2.312589e-07, 
    2.348819e-07, 2.332801e-07, 2.377204e-07, 2.36481e-07, 2.280929e-07, 
    2.284878e-07, 2.298614e-07, 2.29208e-07, 2.310759e-07, 2.315353e-07, 
    2.319086e-07, 2.323857e-07, 2.324372e-07, 2.327198e-07, 2.322567e-07, 
    2.327015e-07, 2.31018e-07, 2.317706e-07, 2.297045e-07, 2.302076e-07, 
    2.299762e-07, 2.297223e-07, 2.305058e-07, 2.313401e-07, 2.313579e-07, 
    2.316253e-07, 2.323784e-07, 2.310834e-07, 2.350885e-07, 2.326163e-07, 
    2.289184e-07, 2.296784e-07, 2.29787e-07, 2.294926e-07, 2.314892e-07, 
    2.307661e-07, 2.327129e-07, 2.32187e-07, 2.330486e-07, 2.326205e-07, 
    2.325575e-07, 2.320075e-07, 2.31665e-07, 2.307993e-07, 2.300945e-07, 
    2.295353e-07, 2.296654e-07, 2.302795e-07, 2.313911e-07, 2.324419e-07, 
    2.322117e-07, 2.329831e-07, 2.309405e-07, 2.317974e-07, 2.314662e-07, 
    2.323295e-07, 2.304374e-07, 2.320487e-07, 2.300252e-07, 2.302027e-07, 
    2.307517e-07, 2.318554e-07, 2.320996e-07, 2.323601e-07, 2.321994e-07, 
    2.314193e-07, 2.312915e-07, 2.307384e-07, 2.305857e-07, 2.301641e-07, 
    2.298149e-07, 2.301339e-07, 2.304688e-07, 2.314196e-07, 2.322759e-07, 
    2.332089e-07, 2.334371e-07, 2.345262e-07, 2.336396e-07, 2.351022e-07, 
    2.338588e-07, 2.360105e-07, 2.32142e-07, 2.338223e-07, 2.307767e-07, 
    2.311052e-07, 2.316989e-07, 2.3306e-07, 2.323254e-07, 2.331845e-07, 
    2.312864e-07, 2.303006e-07, 2.300455e-07, 2.295693e-07, 2.300564e-07, 
    2.300168e-07, 2.304827e-07, 2.30333e-07, 2.314512e-07, 2.308507e-07, 
    2.325559e-07, 2.331777e-07, 2.349322e-07, 2.360066e-07, 2.370995e-07, 
    2.375817e-07, 2.377284e-07, 2.377897e-07,
  2.166374e-07, 2.176639e-07, 2.174644e-07, 2.182922e-07, 2.17833e-07, 
    2.18375e-07, 2.168455e-07, 2.177047e-07, 2.171562e-07, 2.167298e-07, 
    2.198984e-07, 2.183291e-07, 2.21528e-07, 2.205275e-07, 2.230404e-07, 
    2.213723e-07, 2.233767e-07, 2.229923e-07, 2.241491e-07, 2.238177e-07, 
    2.252972e-07, 2.243021e-07, 2.260639e-07, 2.250596e-07, 2.252167e-07, 
    2.242692e-07, 2.18645e-07, 2.197031e-07, 2.185823e-07, 2.187332e-07, 
    2.186655e-07, 2.178425e-07, 2.174277e-07, 2.165589e-07, 2.167167e-07, 
    2.173548e-07, 2.18801e-07, 2.183101e-07, 2.195472e-07, 2.195193e-07, 
    2.208962e-07, 2.202755e-07, 2.225893e-07, 2.219317e-07, 2.238316e-07, 
    2.233539e-07, 2.238091e-07, 2.236711e-07, 2.238109e-07, 2.231103e-07, 
    2.234105e-07, 2.227939e-07, 2.203917e-07, 2.210978e-07, 2.189916e-07, 
    2.177248e-07, 2.168832e-07, 2.162859e-07, 2.163704e-07, 2.165313e-07, 
    2.173585e-07, 2.181361e-07, 2.187285e-07, 2.191248e-07, 2.195153e-07, 
    2.20697e-07, 2.213223e-07, 2.227222e-07, 2.224696e-07, 2.228975e-07, 
    2.233063e-07, 2.239926e-07, 2.238796e-07, 2.241819e-07, 2.228862e-07, 
    2.237474e-07, 2.223257e-07, 2.227146e-07, 2.196215e-07, 2.184426e-07, 
    2.179414e-07, 2.175027e-07, 2.164353e-07, 2.171725e-07, 2.168819e-07, 
    2.175732e-07, 2.180124e-07, 2.177951e-07, 2.191357e-07, 2.186145e-07, 
    2.213594e-07, 2.201773e-07, 2.232586e-07, 2.225214e-07, 2.234353e-07, 
    2.22969e-07, 2.23768e-07, 2.230489e-07, 2.242945e-07, 2.245656e-07, 
    2.243803e-07, 2.250921e-07, 2.230091e-07, 2.238091e-07, 2.177891e-07, 
    2.178245e-07, 2.179895e-07, 2.17264e-07, 2.172196e-07, 2.165546e-07, 
    2.171463e-07, 2.173983e-07, 2.180378e-07, 2.184161e-07, 2.187757e-07, 
    2.195661e-07, 2.204488e-07, 2.216829e-07, 2.225692e-07, 2.231633e-07, 
    2.22799e-07, 2.231207e-07, 2.227611e-07, 2.225926e-07, 2.24464e-07, 
    2.234133e-07, 2.249898e-07, 2.249025e-07, 2.241891e-07, 2.249124e-07, 
    2.178494e-07, 2.176455e-07, 2.169376e-07, 2.174916e-07, 2.164822e-07, 
    2.170472e-07, 2.173721e-07, 2.186254e-07, 2.189008e-07, 2.191561e-07, 
    2.196603e-07, 2.203072e-07, 2.21442e-07, 2.224291e-07, 2.233301e-07, 
    2.232641e-07, 2.232873e-07, 2.234886e-07, 2.229901e-07, 2.235704e-07, 
    2.236678e-07, 2.234132e-07, 2.248909e-07, 2.244687e-07, 2.249007e-07, 
    2.246258e-07, 2.177118e-07, 2.180548e-07, 2.178694e-07, 2.18218e-07, 
    2.179725e-07, 2.190643e-07, 2.193916e-07, 2.209229e-07, 2.202945e-07, 
    2.212946e-07, 2.203961e-07, 2.205553e-07, 2.213272e-07, 2.204446e-07, 
    2.223747e-07, 2.210663e-07, 2.234964e-07, 2.221901e-07, 2.235783e-07, 
    2.233262e-07, 2.237435e-07, 2.241172e-07, 2.245874e-07, 2.254547e-07, 
    2.252539e-07, 2.259791e-07, 2.185662e-07, 2.190111e-07, 2.189719e-07, 
    2.194374e-07, 2.197817e-07, 2.205278e-07, 2.217242e-07, 2.212743e-07, 
    2.221002e-07, 2.222659e-07, 2.210112e-07, 2.217816e-07, 2.193088e-07, 
    2.197084e-07, 2.194705e-07, 2.186013e-07, 2.21378e-07, 2.199532e-07, 
    2.225839e-07, 2.218122e-07, 2.24064e-07, 2.229443e-07, 2.251433e-07, 
    2.260831e-07, 2.269675e-07, 2.280007e-07, 2.192538e-07, 2.189516e-07, 
    2.194928e-07, 2.202415e-07, 2.20936e-07, 2.218593e-07, 2.219538e-07, 
    2.221267e-07, 2.225746e-07, 2.229512e-07, 2.221814e-07, 2.230456e-07, 
    2.198011e-07, 2.215016e-07, 2.188373e-07, 2.196397e-07, 2.201973e-07, 
    2.199527e-07, 2.212229e-07, 2.215222e-07, 2.227383e-07, 2.221097e-07, 
    2.258512e-07, 2.241962e-07, 2.287873e-07, 2.275047e-07, 2.18846e-07, 
    2.192528e-07, 2.206685e-07, 2.199949e-07, 2.219209e-07, 2.223949e-07, 
    2.227802e-07, 2.232726e-07, 2.233258e-07, 2.236175e-07, 2.231394e-07, 
    2.235987e-07, 2.218613e-07, 2.226377e-07, 2.205067e-07, 2.210254e-07, 
    2.207868e-07, 2.20525e-07, 2.213329e-07, 2.221935e-07, 2.222119e-07, 
    2.224878e-07, 2.232653e-07, 2.219287e-07, 2.260648e-07, 2.235109e-07, 
    2.196964e-07, 2.204799e-07, 2.205918e-07, 2.202883e-07, 2.223474e-07, 
    2.216014e-07, 2.236104e-07, 2.230675e-07, 2.23957e-07, 2.23515e-07, 
    2.2345e-07, 2.228823e-07, 2.225288e-07, 2.216356e-07, 2.209087e-07, 
    2.203323e-07, 2.204663e-07, 2.210995e-07, 2.222461e-07, 2.233306e-07, 
    2.230931e-07, 2.238894e-07, 2.217813e-07, 2.226654e-07, 2.223237e-07, 
    2.232146e-07, 2.212623e-07, 2.229249e-07, 2.208373e-07, 2.210204e-07, 
    2.215866e-07, 2.227254e-07, 2.229772e-07, 2.232462e-07, 2.230802e-07, 
    2.222752e-07, 2.221433e-07, 2.215728e-07, 2.214153e-07, 2.209805e-07, 
    2.206205e-07, 2.209494e-07, 2.212948e-07, 2.222756e-07, 2.231593e-07, 
    2.241226e-07, 2.243583e-07, 2.254835e-07, 2.245676e-07, 2.26079e-07, 
    2.247941e-07, 2.270182e-07, 2.230212e-07, 2.247562e-07, 2.216123e-07, 
    2.219511e-07, 2.225639e-07, 2.239689e-07, 2.232104e-07, 2.240974e-07, 
    2.221382e-07, 2.211214e-07, 2.208583e-07, 2.203674e-07, 2.208695e-07, 
    2.208287e-07, 2.213091e-07, 2.211547e-07, 2.223081e-07, 2.216886e-07, 
    2.234484e-07, 2.240904e-07, 2.259032e-07, 2.270141e-07, 2.281447e-07, 
    2.286437e-07, 2.287956e-07, 2.288591e-07,
  2.081373e-07, 2.091061e-07, 2.089177e-07, 2.096995e-07, 2.092658e-07, 
    2.097778e-07, 2.083337e-07, 2.091446e-07, 2.086269e-07, 2.082245e-07, 
    2.11218e-07, 2.097344e-07, 2.127605e-07, 2.118131e-07, 2.141941e-07, 
    2.126131e-07, 2.145131e-07, 2.141484e-07, 2.152462e-07, 2.149316e-07, 
    2.163369e-07, 2.153914e-07, 2.170658e-07, 2.16111e-07, 2.162603e-07, 
    2.153602e-07, 2.100328e-07, 2.110333e-07, 2.099735e-07, 2.101162e-07, 
    2.100521e-07, 2.092748e-07, 2.088832e-07, 2.080633e-07, 2.082121e-07, 
    2.088143e-07, 2.101803e-07, 2.097164e-07, 2.108857e-07, 2.108593e-07, 
    2.121621e-07, 2.115746e-07, 2.137662e-07, 2.131429e-07, 2.149447e-07, 
    2.144914e-07, 2.149234e-07, 2.147924e-07, 2.149252e-07, 2.142603e-07, 
    2.145451e-07, 2.139602e-07, 2.116846e-07, 2.12353e-07, 2.103604e-07, 
    2.091637e-07, 2.083692e-07, 2.078058e-07, 2.078854e-07, 2.080373e-07, 
    2.088178e-07, 2.09552e-07, 2.101117e-07, 2.104863e-07, 2.108555e-07, 
    2.119736e-07, 2.125657e-07, 2.138923e-07, 2.136527e-07, 2.140586e-07, 
    2.144463e-07, 2.150976e-07, 2.149904e-07, 2.152774e-07, 2.140478e-07, 
    2.148649e-07, 2.135163e-07, 2.13885e-07, 2.109561e-07, 2.098415e-07, 
    2.093683e-07, 2.089539e-07, 2.079467e-07, 2.086422e-07, 2.08368e-07, 
    2.090204e-07, 2.094352e-07, 2.0923e-07, 2.104966e-07, 2.10004e-07, 
    2.126008e-07, 2.114817e-07, 2.144011e-07, 2.137019e-07, 2.145687e-07, 
    2.141263e-07, 2.148844e-07, 2.142021e-07, 2.153842e-07, 2.156418e-07, 
    2.154658e-07, 2.161419e-07, 2.141643e-07, 2.149235e-07, 2.092243e-07, 
    2.092577e-07, 2.094136e-07, 2.087286e-07, 2.086867e-07, 2.080592e-07, 
    2.086175e-07, 2.088554e-07, 2.094592e-07, 2.098165e-07, 2.101563e-07, 
    2.109036e-07, 2.117387e-07, 2.129072e-07, 2.137472e-07, 2.143106e-07, 
    2.139651e-07, 2.142701e-07, 2.139292e-07, 2.137694e-07, 2.155453e-07, 
    2.145478e-07, 2.160447e-07, 2.159618e-07, 2.152842e-07, 2.159711e-07, 
    2.092812e-07, 2.090887e-07, 2.084205e-07, 2.089434e-07, 2.079909e-07, 
    2.08524e-07, 2.088307e-07, 2.100144e-07, 2.102745e-07, 2.105159e-07, 
    2.109926e-07, 2.116046e-07, 2.12679e-07, 2.136144e-07, 2.144688e-07, 
    2.144062e-07, 2.144283e-07, 2.146192e-07, 2.141463e-07, 2.146969e-07, 
    2.147894e-07, 2.145477e-07, 2.159507e-07, 2.155497e-07, 2.1596e-07, 
    2.156989e-07, 2.091513e-07, 2.094752e-07, 2.093002e-07, 2.096294e-07, 
    2.093975e-07, 2.104291e-07, 2.107386e-07, 2.121874e-07, 2.115926e-07, 
    2.125394e-07, 2.116887e-07, 2.118394e-07, 2.125704e-07, 2.117347e-07, 
    2.135629e-07, 2.123232e-07, 2.146267e-07, 2.133879e-07, 2.147043e-07, 
    2.144651e-07, 2.148611e-07, 2.152159e-07, 2.156624e-07, 2.164866e-07, 
    2.162957e-07, 2.169852e-07, 2.099583e-07, 2.103788e-07, 2.103417e-07, 
    2.107818e-07, 2.111074e-07, 2.118133e-07, 2.129463e-07, 2.125201e-07, 
    2.133025e-07, 2.134597e-07, 2.12271e-07, 2.130008e-07, 2.106602e-07, 
    2.110382e-07, 2.108131e-07, 2.099915e-07, 2.126184e-07, 2.112697e-07, 
    2.137611e-07, 2.130297e-07, 2.151654e-07, 2.141029e-07, 2.161906e-07, 
    2.170842e-07, 2.179255e-07, 2.189097e-07, 2.106083e-07, 2.103225e-07, 
    2.108342e-07, 2.115425e-07, 2.121998e-07, 2.130743e-07, 2.131638e-07, 
    2.133277e-07, 2.137523e-07, 2.141094e-07, 2.133796e-07, 2.14199e-07, 
    2.111259e-07, 2.127355e-07, 2.102146e-07, 2.109732e-07, 2.115007e-07, 
    2.112692e-07, 2.124714e-07, 2.127549e-07, 2.139076e-07, 2.133116e-07, 
    2.168636e-07, 2.15291e-07, 2.196594e-07, 2.184372e-07, 2.102227e-07, 
    2.106073e-07, 2.119466e-07, 2.113092e-07, 2.131327e-07, 2.135819e-07, 
    2.139472e-07, 2.144143e-07, 2.144648e-07, 2.147416e-07, 2.14288e-07, 
    2.147237e-07, 2.130762e-07, 2.138122e-07, 2.117934e-07, 2.122845e-07, 
    2.120585e-07, 2.118107e-07, 2.125756e-07, 2.133911e-07, 2.134084e-07, 
    2.1367e-07, 2.144076e-07, 2.131401e-07, 2.170669e-07, 2.146406e-07, 
    2.110267e-07, 2.117681e-07, 2.118739e-07, 2.115867e-07, 2.135369e-07, 
    2.1283e-07, 2.147349e-07, 2.142198e-07, 2.150638e-07, 2.146443e-07, 
    2.145826e-07, 2.140441e-07, 2.137089e-07, 2.128624e-07, 2.12174e-07, 
    2.116283e-07, 2.117552e-07, 2.123547e-07, 2.13441e-07, 2.144694e-07, 
    2.14244e-07, 2.149997e-07, 2.130004e-07, 2.138384e-07, 2.135145e-07, 
    2.143593e-07, 2.125088e-07, 2.140846e-07, 2.121063e-07, 2.122797e-07, 
    2.128159e-07, 2.138953e-07, 2.141341e-07, 2.143893e-07, 2.142318e-07, 
    2.134685e-07, 2.133435e-07, 2.128029e-07, 2.126537e-07, 2.122419e-07, 
    2.119011e-07, 2.122125e-07, 2.125396e-07, 2.134688e-07, 2.143068e-07, 
    2.15221e-07, 2.154448e-07, 2.165141e-07, 2.156437e-07, 2.170804e-07, 
    2.15859e-07, 2.17974e-07, 2.141759e-07, 2.158229e-07, 2.128403e-07, 
    2.131613e-07, 2.137422e-07, 2.150752e-07, 2.143553e-07, 2.151972e-07, 
    2.133386e-07, 2.123754e-07, 2.121262e-07, 2.116615e-07, 2.121368e-07, 
    2.120981e-07, 2.125531e-07, 2.124069e-07, 2.134997e-07, 2.129126e-07, 
    2.145811e-07, 2.151905e-07, 2.169129e-07, 2.1797e-07, 2.190467e-07, 
    2.195224e-07, 2.196672e-07, 2.197278e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371698e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441075e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379093e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377207e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523353e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.56315e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529406e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.532169e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547246e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.46224e-08, 6.465288e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532766e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472856e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  8.591897e-13, 8.615078e-13, 8.610575e-13, 8.629254e-13, 8.618897e-13, 
    8.631123e-13, 8.596602e-13, 8.615995e-13, 8.603619e-13, 8.593989e-13, 
    8.66545e-13, 8.630088e-13, 8.702151e-13, 8.679639e-13, 8.736153e-13, 
    8.698645e-13, 8.743711e-13, 8.735079e-13, 8.761065e-13, 8.753624e-13, 
    8.78681e-13, 8.764498e-13, 8.804005e-13, 8.781488e-13, 8.785009e-13, 
    8.76376e-13, 8.637216e-13, 8.661048e-13, 8.635801e-13, 8.639202e-13, 
    8.637678e-13, 8.619109e-13, 8.60974e-13, 8.590129e-13, 8.593692e-13, 
    8.608098e-13, 8.640731e-13, 8.629664e-13, 8.65756e-13, 8.656931e-13, 
    8.687941e-13, 8.673965e-13, 8.726022e-13, 8.711244e-13, 8.753935e-13, 
    8.743204e-13, 8.75343e-13, 8.750331e-13, 8.75347e-13, 8.737731e-13, 
    8.744475e-13, 8.730623e-13, 8.676582e-13, 8.692477e-13, 8.645031e-13, 
    8.616442e-13, 8.597451e-13, 8.58396e-13, 8.585868e-13, 8.589503e-13, 
    8.608182e-13, 8.625737e-13, 8.639103e-13, 8.648039e-13, 8.65684e-13, 
    8.683441e-13, 8.697523e-13, 8.729006e-13, 8.723333e-13, 8.732947e-13, 
    8.742137e-13, 8.757548e-13, 8.755013e-13, 8.761798e-13, 8.732698e-13, 
    8.75204e-13, 8.720105e-13, 8.72884e-13, 8.659207e-13, 8.632651e-13, 
    8.621332e-13, 8.611439e-13, 8.587334e-13, 8.603982e-13, 8.59742e-13, 
    8.613034e-13, 8.622946e-13, 8.618045e-13, 8.648283e-13, 8.636531e-13, 
    8.698358e-13, 8.671749e-13, 8.741065e-13, 8.724498e-13, 8.745035e-13, 
    8.734559e-13, 8.752503e-13, 8.736355e-13, 8.764325e-13, 8.770408e-13, 
    8.766251e-13, 8.782224e-13, 8.735458e-13, 8.753427e-13, 8.617907e-13, 
    8.618706e-13, 8.622432e-13, 8.606048e-13, 8.605048e-13, 8.59003e-13, 
    8.603395e-13, 8.609082e-13, 8.623522e-13, 8.632054e-13, 8.640164e-13, 
    8.657984e-13, 8.677864e-13, 8.70564e-13, 8.725572e-13, 8.738925e-13, 
    8.73074e-13, 8.737966e-13, 8.729887e-13, 8.7261e-13, 8.768127e-13, 
    8.744536e-13, 8.779927e-13, 8.777971e-13, 8.761959e-13, 8.778192e-13, 
    8.619267e-13, 8.614667e-13, 8.598681e-13, 8.611192e-13, 8.588395e-13, 
    8.601155e-13, 8.608488e-13, 8.636771e-13, 8.642987e-13, 8.648741e-13, 
    8.660106e-13, 8.67468e-13, 8.700222e-13, 8.72242e-13, 8.742672e-13, 
    8.74119e-13, 8.741711e-13, 8.746231e-13, 8.735031e-13, 8.748069e-13, 
    8.750254e-13, 8.744537e-13, 8.777709e-13, 8.768238e-13, 8.77793e-13, 
    8.771764e-13, 8.616163e-13, 8.623903e-13, 8.619721e-13, 8.627584e-13, 
    8.622042e-13, 8.646666e-13, 8.654043e-13, 8.688535e-13, 8.674392e-13, 
    8.696903e-13, 8.676682e-13, 8.680265e-13, 8.697626e-13, 8.677777e-13, 
    8.721191e-13, 8.691759e-13, 8.746406e-13, 8.717039e-13, 8.748245e-13, 
    8.742585e-13, 8.751958e-13, 8.760347e-13, 8.7709e-13, 8.79035e-13, 
    8.785849e-13, 8.802109e-13, 8.63544e-13, 8.645469e-13, 8.644591e-13, 
    8.655085e-13, 8.66284e-13, 8.679648e-13, 8.706572e-13, 8.696453e-13, 
    8.715032e-13, 8.718759e-13, 8.690534e-13, 8.707863e-13, 8.652181e-13, 
    8.661182e-13, 8.655827e-13, 8.636229e-13, 8.698778e-13, 8.666697e-13, 
    8.725901e-13, 8.708555e-13, 8.75915e-13, 8.733995e-13, 8.783369e-13, 
    8.804428e-13, 8.824252e-13, 8.847366e-13, 8.650945e-13, 8.644133e-13, 
    8.656333e-13, 8.673193e-13, 8.688838e-13, 8.709612e-13, 8.71174e-13, 
    8.715628e-13, 8.725696e-13, 8.73416e-13, 8.716852e-13, 8.736282e-13, 
    8.663259e-13, 8.701563e-13, 8.641552e-13, 8.659634e-13, 8.672201e-13, 
    8.666694e-13, 8.695298e-13, 8.702032e-13, 8.729369e-13, 8.715247e-13, 
    8.799228e-13, 8.762111e-13, 8.864965e-13, 8.83627e-13, 8.641751e-13, 
    8.650924e-13, 8.682811e-13, 8.667646e-13, 8.711001e-13, 8.721653e-13, 
    8.730316e-13, 8.741377e-13, 8.742575e-13, 8.749126e-13, 8.738389e-13, 
    8.748704e-13, 8.709657e-13, 8.727113e-13, 8.679175e-13, 8.690851e-13, 
    8.685482e-13, 8.679588e-13, 8.697773e-13, 8.717123e-13, 8.717544e-13, 
    8.723739e-13, 8.741185e-13, 8.711177e-13, 8.803999e-13, 8.746705e-13, 
    8.660921e-13, 8.67856e-13, 8.681088e-13, 8.674256e-13, 8.720589e-13, 
    8.703811e-13, 8.748967e-13, 8.736773e-13, 8.756752e-13, 8.746825e-13, 
    8.745364e-13, 8.73261e-13, 8.724663e-13, 8.704579e-13, 8.688223e-13, 
    8.675248e-13, 8.678266e-13, 8.692517e-13, 8.718308e-13, 8.742679e-13, 
    8.737341e-13, 8.755234e-13, 8.70786e-13, 8.727731e-13, 8.720053e-13, 
    8.740076e-13, 8.696182e-13, 8.733541e-13, 8.686619e-13, 8.690739e-13, 
    8.703478e-13, 8.729073e-13, 8.734744e-13, 8.740784e-13, 8.737059e-13, 
    8.718964e-13, 8.716e-13, 8.703171e-13, 8.699623e-13, 8.689842e-13, 
    8.681738e-13, 8.689141e-13, 8.696911e-13, 8.718975e-13, 8.73883e-13, 
    8.760465e-13, 8.765759e-13, 8.790982e-13, 8.77044e-13, 8.804316e-13, 
    8.775502e-13, 8.825364e-13, 8.735716e-13, 8.77467e-13, 8.70406e-13, 
    8.711681e-13, 8.725444e-13, 8.757007e-13, 8.739981e-13, 8.759895e-13, 
    8.715886e-13, 8.693005e-13, 8.68709e-13, 8.676036e-13, 8.687343e-13, 
    8.686424e-13, 8.697238e-13, 8.693764e-13, 8.719707e-13, 8.705776e-13, 
    8.745325e-13, 8.75974e-13, 8.800403e-13, 8.825286e-13, 8.850598e-13, 
    8.861758e-13, 8.865154e-13, 8.866573e-13 ;

 LITR1C =
  3.066802e-05, 3.066791e-05, 3.066793e-05, 3.066783e-05, 3.066788e-05, 
    3.066782e-05, 3.0668e-05, 3.06679e-05, 3.066796e-05, 3.066801e-05, 
    3.066765e-05, 3.066783e-05, 3.066747e-05, 3.066758e-05, 3.06673e-05, 
    3.066748e-05, 3.066726e-05, 3.06673e-05, 3.066717e-05, 3.066721e-05, 
    3.066704e-05, 3.066715e-05, 3.066696e-05, 3.066707e-05, 3.066705e-05, 
    3.066716e-05, 3.066779e-05, 3.066767e-05, 3.06678e-05, 3.066778e-05, 
    3.066779e-05, 3.066788e-05, 3.066793e-05, 3.066803e-05, 3.066801e-05, 
    3.066794e-05, 3.066778e-05, 3.066783e-05, 3.066769e-05, 3.06677e-05, 
    3.066754e-05, 3.066761e-05, 3.066735e-05, 3.066742e-05, 3.066721e-05, 
    3.066726e-05, 3.066721e-05, 3.066723e-05, 3.066721e-05, 3.066729e-05, 
    3.066726e-05, 3.066732e-05, 3.06676e-05, 3.066752e-05, 3.066775e-05, 
    3.06679e-05, 3.066799e-05, 3.066806e-05, 3.066805e-05, 3.066803e-05, 
    3.066794e-05, 3.066785e-05, 3.066778e-05, 3.066774e-05, 3.06677e-05, 
    3.066756e-05, 3.066749e-05, 3.066733e-05, 3.066736e-05, 3.066731e-05, 
    3.066727e-05, 3.066719e-05, 3.06672e-05, 3.066717e-05, 3.066731e-05, 
    3.066722e-05, 3.066738e-05, 3.066733e-05, 3.066768e-05, 3.066782e-05, 
    3.066787e-05, 3.066792e-05, 3.066804e-05, 3.066796e-05, 3.066799e-05, 
    3.066791e-05, 3.066787e-05, 3.066789e-05, 3.066774e-05, 3.06678e-05, 
    3.066749e-05, 3.066762e-05, 3.066727e-05, 3.066735e-05, 3.066725e-05, 
    3.066731e-05, 3.066722e-05, 3.06673e-05, 3.066715e-05, 3.066712e-05, 
    3.066715e-05, 3.066707e-05, 3.06673e-05, 3.066721e-05, 3.066789e-05, 
    3.066789e-05, 3.066787e-05, 3.066795e-05, 3.066795e-05, 3.066803e-05, 
    3.066796e-05, 3.066794e-05, 3.066786e-05, 3.066782e-05, 3.066778e-05, 
    3.066769e-05, 3.066759e-05, 3.066745e-05, 3.066735e-05, 3.066728e-05, 
    3.066732e-05, 3.066729e-05, 3.066733e-05, 3.066735e-05, 3.066714e-05, 
    3.066726e-05, 3.066708e-05, 3.066709e-05, 3.066717e-05, 3.066708e-05, 
    3.066788e-05, 3.066791e-05, 3.066799e-05, 3.066792e-05, 3.066804e-05, 
    3.066798e-05, 3.066794e-05, 3.06678e-05, 3.066776e-05, 3.066774e-05, 
    3.066768e-05, 3.06676e-05, 3.066748e-05, 3.066736e-05, 3.066726e-05, 
    3.066727e-05, 3.066727e-05, 3.066724e-05, 3.06673e-05, 3.066724e-05, 
    3.066723e-05, 3.066726e-05, 3.066709e-05, 3.066714e-05, 3.066709e-05, 
    3.066712e-05, 3.06679e-05, 3.066786e-05, 3.066788e-05, 3.066784e-05, 
    3.066787e-05, 3.066775e-05, 3.066771e-05, 3.066754e-05, 3.066761e-05, 
    3.06675e-05, 3.066759e-05, 3.066758e-05, 3.066749e-05, 3.066759e-05, 
    3.066737e-05, 3.066752e-05, 3.066724e-05, 3.066739e-05, 3.066724e-05, 
    3.066726e-05, 3.066722e-05, 3.066718e-05, 3.066712e-05, 3.066702e-05, 
    3.066705e-05, 3.066696e-05, 3.06678e-05, 3.066775e-05, 3.066776e-05, 
    3.06677e-05, 3.066767e-05, 3.066758e-05, 3.066744e-05, 3.06675e-05, 
    3.06674e-05, 3.066738e-05, 3.066752e-05, 3.066744e-05, 3.066772e-05, 
    3.066767e-05, 3.06677e-05, 3.06678e-05, 3.066748e-05, 3.066764e-05, 
    3.066735e-05, 3.066743e-05, 3.066718e-05, 3.066731e-05, 3.066706e-05, 
    3.066695e-05, 3.066686e-05, 3.066674e-05, 3.066772e-05, 3.066776e-05, 
    3.06677e-05, 3.066761e-05, 3.066754e-05, 3.066743e-05, 3.066742e-05, 
    3.06674e-05, 3.066735e-05, 3.066731e-05, 3.066739e-05, 3.06673e-05, 
    3.066766e-05, 3.066747e-05, 3.066777e-05, 3.066768e-05, 3.066762e-05, 
    3.066764e-05, 3.06675e-05, 3.066747e-05, 3.066733e-05, 3.06674e-05, 
    3.066698e-05, 3.066716e-05, 3.066665e-05, 3.066679e-05, 3.066777e-05, 
    3.066772e-05, 3.066756e-05, 3.066764e-05, 3.066742e-05, 3.066737e-05, 
    3.066732e-05, 3.066727e-05, 3.066726e-05, 3.066723e-05, 3.066728e-05, 
    3.066723e-05, 3.066743e-05, 3.066734e-05, 3.066758e-05, 3.066752e-05, 
    3.066755e-05, 3.066758e-05, 3.066749e-05, 3.066739e-05, 3.066739e-05, 
    3.066736e-05, 3.066727e-05, 3.066742e-05, 3.066696e-05, 3.066724e-05, 
    3.066767e-05, 3.066759e-05, 3.066757e-05, 3.066761e-05, 3.066738e-05, 
    3.066746e-05, 3.066723e-05, 3.066729e-05, 3.066719e-05, 3.066724e-05, 
    3.066725e-05, 3.066731e-05, 3.066735e-05, 3.066746e-05, 3.066754e-05, 
    3.06676e-05, 3.066759e-05, 3.066752e-05, 3.066739e-05, 3.066726e-05, 
    3.066729e-05, 3.06672e-05, 3.066744e-05, 3.066734e-05, 3.066738e-05, 
    3.066728e-05, 3.06675e-05, 3.066731e-05, 3.066755e-05, 3.066752e-05, 
    3.066746e-05, 3.066733e-05, 3.06673e-05, 3.066727e-05, 3.066729e-05, 
    3.066738e-05, 3.06674e-05, 3.066746e-05, 3.066748e-05, 3.066753e-05, 
    3.066757e-05, 3.066753e-05, 3.06675e-05, 3.066738e-05, 3.066728e-05, 
    3.066718e-05, 3.066715e-05, 3.066702e-05, 3.066712e-05, 3.066695e-05, 
    3.06671e-05, 3.066685e-05, 3.06673e-05, 3.06671e-05, 3.066746e-05, 
    3.066742e-05, 3.066735e-05, 3.066719e-05, 3.066728e-05, 3.066718e-05, 
    3.06674e-05, 3.066751e-05, 3.066754e-05, 3.06676e-05, 3.066754e-05, 
    3.066755e-05, 3.066749e-05, 3.066751e-05, 3.066738e-05, 3.066745e-05, 
    3.066725e-05, 3.066718e-05, 3.066698e-05, 3.066685e-05, 3.066672e-05, 
    3.066667e-05, 3.066665e-05, 3.066664e-05 ;

 LITR1C_TO_SOIL1C =
  5.722613e-13, 5.738049e-13, 5.735051e-13, 5.74749e-13, 5.740592e-13, 
    5.748734e-13, 5.725745e-13, 5.73866e-13, 5.730418e-13, 5.724006e-13, 
    5.771593e-13, 5.748045e-13, 5.796034e-13, 5.781042e-13, 5.818676e-13, 
    5.793699e-13, 5.823709e-13, 5.817962e-13, 5.835266e-13, 5.830311e-13, 
    5.85241e-13, 5.837552e-13, 5.86386e-13, 5.848866e-13, 5.851211e-13, 
    5.837061e-13, 5.752792e-13, 5.768662e-13, 5.75185e-13, 5.754114e-13, 
    5.753099e-13, 5.740733e-13, 5.734495e-13, 5.721435e-13, 5.723808e-13, 
    5.733401e-13, 5.755133e-13, 5.747763e-13, 5.76634e-13, 5.765921e-13, 
    5.786571e-13, 5.777264e-13, 5.81193e-13, 5.802089e-13, 5.830518e-13, 
    5.823372e-13, 5.830181e-13, 5.828117e-13, 5.830208e-13, 5.819727e-13, 
    5.824219e-13, 5.814994e-13, 5.779006e-13, 5.789591e-13, 5.757996e-13, 
    5.738957e-13, 5.726311e-13, 5.717327e-13, 5.718598e-13, 5.721018e-13, 
    5.733457e-13, 5.745147e-13, 5.754048e-13, 5.759999e-13, 5.76586e-13, 
    5.783574e-13, 5.792952e-13, 5.813917e-13, 5.81014e-13, 5.816541e-13, 
    5.822661e-13, 5.832924e-13, 5.831236e-13, 5.835754e-13, 5.816376e-13, 
    5.829256e-13, 5.80799e-13, 5.813806e-13, 5.767436e-13, 5.749752e-13, 
    5.742214e-13, 5.735626e-13, 5.719574e-13, 5.730661e-13, 5.726291e-13, 
    5.736688e-13, 5.743289e-13, 5.740025e-13, 5.760162e-13, 5.752335e-13, 
    5.793508e-13, 5.775788e-13, 5.821948e-13, 5.810915e-13, 5.824591e-13, 
    5.817615e-13, 5.829565e-13, 5.818811e-13, 5.837437e-13, 5.841487e-13, 
    5.838719e-13, 5.849356e-13, 5.818214e-13, 5.83018e-13, 5.739933e-13, 
    5.740465e-13, 5.742946e-13, 5.732036e-13, 5.73137e-13, 5.72137e-13, 
    5.73027e-13, 5.734057e-13, 5.743673e-13, 5.749354e-13, 5.754755e-13, 
    5.766621e-13, 5.77986e-13, 5.798357e-13, 5.81163e-13, 5.820523e-13, 
    5.815072e-13, 5.819884e-13, 5.814504e-13, 5.811982e-13, 5.839969e-13, 
    5.824259e-13, 5.847827e-13, 5.846524e-13, 5.835861e-13, 5.846671e-13, 
    5.740839e-13, 5.737776e-13, 5.72713e-13, 5.735462e-13, 5.72028e-13, 
    5.728778e-13, 5.733661e-13, 5.752495e-13, 5.756635e-13, 5.760466e-13, 
    5.768035e-13, 5.77774e-13, 5.794749e-13, 5.809531e-13, 5.823018e-13, 
    5.822031e-13, 5.822378e-13, 5.825387e-13, 5.817929e-13, 5.826611e-13, 
    5.828066e-13, 5.824259e-13, 5.84635e-13, 5.840043e-13, 5.846497e-13, 
    5.84239e-13, 5.738772e-13, 5.743927e-13, 5.741141e-13, 5.746378e-13, 
    5.742688e-13, 5.759085e-13, 5.763997e-13, 5.786967e-13, 5.777548e-13, 
    5.792539e-13, 5.779073e-13, 5.781459e-13, 5.79302e-13, 5.779802e-13, 
    5.808713e-13, 5.789113e-13, 5.825504e-13, 5.805948e-13, 5.826729e-13, 
    5.822959e-13, 5.829202e-13, 5.834787e-13, 5.841815e-13, 5.854768e-13, 
    5.85177e-13, 5.862598e-13, 5.751609e-13, 5.758287e-13, 5.757703e-13, 
    5.764691e-13, 5.769856e-13, 5.781048e-13, 5.798978e-13, 5.79224e-13, 
    5.804612e-13, 5.807093e-13, 5.788297e-13, 5.799838e-13, 5.762757e-13, 
    5.768751e-13, 5.765185e-13, 5.752134e-13, 5.793788e-13, 5.772424e-13, 
    5.811849e-13, 5.800298e-13, 5.833991e-13, 5.81724e-13, 5.850119e-13, 
    5.864142e-13, 5.877343e-13, 5.892736e-13, 5.761934e-13, 5.757398e-13, 
    5.765523e-13, 5.77675e-13, 5.787168e-13, 5.801003e-13, 5.802419e-13, 
    5.805008e-13, 5.811713e-13, 5.817349e-13, 5.805823e-13, 5.818762e-13, 
    5.770135e-13, 5.795642e-13, 5.755679e-13, 5.76772e-13, 5.776089e-13, 
    5.772422e-13, 5.79147e-13, 5.795955e-13, 5.814159e-13, 5.804754e-13, 
    5.86068e-13, 5.835962e-13, 5.904455e-13, 5.885346e-13, 5.755811e-13, 
    5.76192e-13, 5.783155e-13, 5.773056e-13, 5.801927e-13, 5.80902e-13, 
    5.814789e-13, 5.822155e-13, 5.822953e-13, 5.827316e-13, 5.820165e-13, 
    5.827034e-13, 5.801032e-13, 5.812657e-13, 5.780733e-13, 5.788508e-13, 
    5.784933e-13, 5.781008e-13, 5.793118e-13, 5.806004e-13, 5.806284e-13, 
    5.81041e-13, 5.822027e-13, 5.802044e-13, 5.863856e-13, 5.825703e-13, 
    5.768578e-13, 5.780324e-13, 5.782007e-13, 5.777458e-13, 5.808312e-13, 
    5.797139e-13, 5.82721e-13, 5.819089e-13, 5.832393e-13, 5.825784e-13, 
    5.824811e-13, 5.816317e-13, 5.811025e-13, 5.797651e-13, 5.786759e-13, 
    5.778118e-13, 5.780128e-13, 5.789618e-13, 5.806793e-13, 5.823023e-13, 
    5.819468e-13, 5.831383e-13, 5.799835e-13, 5.813068e-13, 5.807955e-13, 
    5.821289e-13, 5.792059e-13, 5.816937e-13, 5.78569e-13, 5.788434e-13, 
    5.796917e-13, 5.813962e-13, 5.817738e-13, 5.82176e-13, 5.81928e-13, 
    5.80723e-13, 5.805256e-13, 5.796712e-13, 5.79435e-13, 5.787837e-13, 
    5.78244e-13, 5.78737e-13, 5.792544e-13, 5.807237e-13, 5.820459e-13, 
    5.834866e-13, 5.838391e-13, 5.855188e-13, 5.841509e-13, 5.864068e-13, 
    5.84488e-13, 5.878084e-13, 5.818385e-13, 5.844326e-13, 5.797305e-13, 
    5.80238e-13, 5.811545e-13, 5.832564e-13, 5.821226e-13, 5.834487e-13, 
    5.805179e-13, 5.789943e-13, 5.786004e-13, 5.778643e-13, 5.786172e-13, 
    5.78556e-13, 5.792762e-13, 5.790448e-13, 5.807725e-13, 5.798448e-13, 
    5.824785e-13, 5.834384e-13, 5.861462e-13, 5.878032e-13, 5.894888e-13, 
    5.90232e-13, 5.904581e-13, 5.905526e-13 ;

 LITR1C_vr =
  0.001751176, 0.001751169, 0.00175117, 0.001751165, 0.001751168, 
    0.001751164, 0.001751174, 0.001751169, 0.001751172, 0.001751175, 
    0.001751155, 0.001751165, 0.001751144, 0.001751151, 0.001751134, 
    0.001751145, 0.001751132, 0.001751135, 0.001751127, 0.001751129, 
    0.00175112, 0.001751126, 0.001751115, 0.001751121, 0.00175112, 
    0.001751126, 0.001751163, 0.001751156, 0.001751163, 0.001751162, 
    0.001751163, 0.001751168, 0.001751171, 0.001751176, 0.001751175, 
    0.001751171, 0.001751162, 0.001751165, 0.001751157, 0.001751157, 
    0.001751148, 0.001751152, 0.001751137, 0.001751142, 0.001751129, 
    0.001751132, 0.001751129, 0.00175113, 0.001751129, 0.001751134, 
    0.001751132, 0.001751136, 0.001751151, 0.001751147, 0.00175116, 
    0.001751169, 0.001751174, 0.001751178, 0.001751177, 0.001751176, 
    0.001751171, 0.001751166, 0.001751162, 0.00175116, 0.001751157, 
    0.001751149, 0.001751145, 0.001751136, 0.001751138, 0.001751135, 
    0.001751133, 0.001751128, 0.001751129, 0.001751127, 0.001751135, 
    0.00175113, 0.001751139, 0.001751136, 0.001751156, 0.001751164, 
    0.001751167, 0.00175117, 0.001751177, 0.001751172, 0.001751174, 
    0.00175117, 0.001751167, 0.001751168, 0.00175116, 0.001751163, 
    0.001751145, 0.001751153, 0.001751133, 0.001751138, 0.001751132, 
    0.001751135, 0.00175113, 0.001751134, 0.001751126, 0.001751125, 
    0.001751126, 0.001751121, 0.001751135, 0.001751129, 0.001751168, 
    0.001751168, 0.001751167, 0.001751172, 0.001751172, 0.001751176, 
    0.001751172, 0.001751171, 0.001751167, 0.001751164, 0.001751162, 
    0.001751157, 0.001751151, 0.001751143, 0.001751137, 0.001751134, 
    0.001751136, 0.001751134, 0.001751136, 0.001751137, 0.001751125, 
    0.001751132, 0.001751122, 0.001751122, 0.001751127, 0.001751122, 
    0.001751168, 0.001751169, 0.001751174, 0.00175117, 0.001751177, 
    0.001751173, 0.001751171, 0.001751163, 0.001751161, 0.001751159, 
    0.001751156, 0.001751152, 0.001751145, 0.001751138, 0.001751132, 
    0.001751133, 0.001751133, 0.001751131, 0.001751135, 0.001751131, 
    0.00175113, 0.001751132, 0.001751122, 0.001751125, 0.001751122, 
    0.001751124, 0.001751169, 0.001751167, 0.001751168, 0.001751165, 
    0.001751167, 0.00175116, 0.001751158, 0.001751148, 0.001751152, 
    0.001751146, 0.001751151, 0.00175115, 0.001751145, 0.001751151, 
    0.001751139, 0.001751147, 0.001751131, 0.00175114, 0.001751131, 
    0.001751133, 0.00175113, 0.001751127, 0.001751124, 0.001751119, 
    0.00175112, 0.001751115, 0.001751163, 0.00175116, 0.001751161, 
    0.001751158, 0.001751155, 0.001751151, 0.001751143, 0.001751146, 
    0.00175114, 0.001751139, 0.001751147, 0.001751142, 0.001751158, 
    0.001751156, 0.001751157, 0.001751163, 0.001751145, 0.001751154, 
    0.001751137, 0.001751142, 0.001751128, 0.001751135, 0.001751121, 
    0.001751115, 0.001751109, 0.001751102, 0.001751159, 0.001751161, 
    0.001751157, 0.001751152, 0.001751148, 0.001751142, 0.001751141, 
    0.00175114, 0.001751137, 0.001751135, 0.00175114, 0.001751134, 
    0.001751155, 0.001751144, 0.001751162, 0.001751156, 0.001751153, 
    0.001751154, 0.001751146, 0.001751144, 0.001751136, 0.00175114, 
    0.001751116, 0.001751127, 0.001751097, 0.001751106, 0.001751161, 
    0.001751159, 0.00175115, 0.001751154, 0.001751142, 0.001751138, 
    0.001751136, 0.001751133, 0.001751133, 0.001751131, 0.001751134, 
    0.001751131, 0.001751142, 0.001751137, 0.001751151, 0.001751147, 
    0.001751149, 0.001751151, 0.001751145, 0.00175114, 0.00175114, 
    0.001751138, 0.001751133, 0.001751142, 0.001751115, 0.001751131, 
    0.001751156, 0.001751151, 0.00175115, 0.001751152, 0.001751139, 
    0.001751144, 0.001751131, 0.001751134, 0.001751128, 0.001751131, 
    0.001751132, 0.001751135, 0.001751138, 0.001751143, 0.001751148, 
    0.001751152, 0.001751151, 0.001751147, 0.001751139, 0.001751132, 
    0.001751134, 0.001751129, 0.001751142, 0.001751137, 0.001751139, 
    0.001751133, 0.001751146, 0.001751135, 0.001751148, 0.001751147, 
    0.001751144, 0.001751136, 0.001751135, 0.001751133, 0.001751134, 
    0.001751139, 0.00175114, 0.001751144, 0.001751145, 0.001751148, 
    0.00175115, 0.001751148, 0.001751146, 0.001751139, 0.001751134, 
    0.001751127, 0.001751126, 0.001751119, 0.001751125, 0.001751115, 
    0.001751123, 0.001751109, 0.001751134, 0.001751123, 0.001751143, 
    0.001751141, 0.001751137, 0.001751128, 0.001751133, 0.001751128, 
    0.00175114, 0.001751147, 0.001751148, 0.001751152, 0.001751148, 
    0.001751149, 0.001751145, 0.001751147, 0.001751139, 0.001751143, 
    0.001751132, 0.001751128, 0.001751116, 0.001751109, 0.001751101, 
    0.001751098, 0.001751097, 0.001751097,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.73289e-07, 9.732854e-07, 9.732861e-07, 9.732831e-07, 9.732847e-07, 
    9.732828e-07, 9.732884e-07, 9.732853e-07, 9.732872e-07, 9.732887e-07, 
    9.732773e-07, 9.73283e-07, 9.732715e-07, 9.732751e-07, 9.732661e-07, 
    9.732721e-07, 9.732648e-07, 9.732663e-07, 9.732621e-07, 9.732632e-07, 
    9.73258e-07, 9.732615e-07, 9.732553e-07, 9.732588e-07, 9.732582e-07, 
    9.732616e-07, 9.732819e-07, 9.73278e-07, 9.732821e-07, 9.732815e-07, 
    9.732818e-07, 9.732847e-07, 9.732862e-07, 9.732894e-07, 9.732888e-07, 
    9.732865e-07, 9.732813e-07, 9.73283e-07, 9.732786e-07, 9.732787e-07, 
    9.732738e-07, 9.73276e-07, 9.732677e-07, 9.732701e-07, 9.732632e-07, 
    9.732649e-07, 9.732634e-07, 9.732638e-07, 9.732634e-07, 9.732659e-07, 
    9.732647e-07, 9.73267e-07, 9.732756e-07, 9.73273e-07, 9.732806e-07, 
    9.732852e-07, 9.732883e-07, 9.732904e-07, 9.732901e-07, 9.732895e-07, 
    9.732865e-07, 9.732837e-07, 9.732815e-07, 9.732802e-07, 9.732787e-07, 
    9.732745e-07, 9.732722e-07, 9.732672e-07, 9.732681e-07, 9.732665e-07, 
    9.732652e-07, 9.732627e-07, 9.732631e-07, 9.73262e-07, 9.732667e-07, 
    9.732636e-07, 9.732687e-07, 9.732672e-07, 9.732784e-07, 9.732826e-07, 
    9.732844e-07, 9.73286e-07, 9.732898e-07, 9.732871e-07, 9.732883e-07, 
    9.732858e-07, 9.732842e-07, 9.73285e-07, 9.732801e-07, 9.73282e-07, 
    9.732721e-07, 9.732763e-07, 9.732653e-07, 9.732679e-07, 9.732647e-07, 
    9.732663e-07, 9.732635e-07, 9.732661e-07, 9.732615e-07, 9.732606e-07, 
    9.732613e-07, 9.732587e-07, 9.732662e-07, 9.732634e-07, 9.73285e-07, 
    9.732848e-07, 9.732843e-07, 9.732869e-07, 9.73287e-07, 9.732894e-07, 
    9.732872e-07, 9.732863e-07, 9.73284e-07, 9.732827e-07, 9.732814e-07, 
    9.732786e-07, 9.732754e-07, 9.73271e-07, 9.732678e-07, 9.732656e-07, 
    9.73267e-07, 9.732657e-07, 9.732671e-07, 9.732677e-07, 9.73261e-07, 
    9.732647e-07, 9.732591e-07, 9.732594e-07, 9.73262e-07, 9.732594e-07, 
    9.732847e-07, 9.732854e-07, 9.73288e-07, 9.73286e-07, 9.732896e-07, 
    9.732876e-07, 9.732864e-07, 9.732819e-07, 9.73281e-07, 9.732801e-07, 
    9.732782e-07, 9.732759e-07, 9.732718e-07, 9.732682e-07, 9.732651e-07, 
    9.732653e-07, 9.732652e-07, 9.732645e-07, 9.732663e-07, 9.732642e-07, 
    9.732638e-07, 9.732647e-07, 9.732595e-07, 9.73261e-07, 9.732594e-07, 
    9.732604e-07, 9.732852e-07, 9.732839e-07, 9.732846e-07, 9.732834e-07, 
    9.732843e-07, 9.732804e-07, 9.732792e-07, 9.732737e-07, 9.73276e-07, 
    9.732723e-07, 9.732755e-07, 9.73275e-07, 9.732722e-07, 9.732754e-07, 
    9.732685e-07, 9.732731e-07, 9.732645e-07, 9.732692e-07, 9.732642e-07, 
    9.732651e-07, 9.732636e-07, 9.732622e-07, 9.732605e-07, 9.732574e-07, 
    9.732581e-07, 9.732556e-07, 9.732821e-07, 9.732805e-07, 9.732806e-07, 
    9.73279e-07, 9.732778e-07, 9.732751e-07, 9.732707e-07, 9.732724e-07, 
    9.732695e-07, 9.732688e-07, 9.732734e-07, 9.732706e-07, 9.732795e-07, 
    9.73278e-07, 9.732789e-07, 9.73282e-07, 9.73272e-07, 9.732771e-07, 
    9.732677e-07, 9.732705e-07, 9.732624e-07, 9.732664e-07, 9.732586e-07, 
    9.732552e-07, 9.73252e-07, 9.732483e-07, 9.732797e-07, 9.732807e-07, 
    9.732788e-07, 9.732761e-07, 9.732736e-07, 9.732703e-07, 9.732699e-07, 
    9.732694e-07, 9.732678e-07, 9.732664e-07, 9.732692e-07, 9.732661e-07, 
    9.732777e-07, 9.732717e-07, 9.732812e-07, 9.732782e-07, 9.732763e-07, 
    9.732771e-07, 9.732726e-07, 9.732715e-07, 9.732672e-07, 9.732694e-07, 
    9.732561e-07, 9.73262e-07, 9.732455e-07, 9.732502e-07, 9.732811e-07, 
    9.732797e-07, 9.732746e-07, 9.73277e-07, 9.732701e-07, 9.732684e-07, 
    9.73267e-07, 9.732653e-07, 9.732651e-07, 9.73264e-07, 9.732657e-07, 
    9.73264e-07, 9.732703e-07, 9.732676e-07, 9.732752e-07, 9.732734e-07, 
    9.732742e-07, 9.732751e-07, 9.732722e-07, 9.732692e-07, 9.73269e-07, 
    9.73268e-07, 9.732653e-07, 9.732701e-07, 9.732553e-07, 9.732644e-07, 
    9.732781e-07, 9.732753e-07, 9.732748e-07, 9.73276e-07, 9.732686e-07, 
    9.732712e-07, 9.73264e-07, 9.73266e-07, 9.732628e-07, 9.732644e-07, 
    9.732646e-07, 9.732667e-07, 9.732679e-07, 9.732711e-07, 9.732737e-07, 
    9.732757e-07, 9.732753e-07, 9.73273e-07, 9.732689e-07, 9.732651e-07, 
    9.732659e-07, 9.73263e-07, 9.732706e-07, 9.732674e-07, 9.732687e-07, 
    9.732654e-07, 9.732724e-07, 9.732665e-07, 9.732739e-07, 9.732734e-07, 
    9.732713e-07, 9.732672e-07, 9.732663e-07, 9.732653e-07, 9.73266e-07, 
    9.732688e-07, 9.732693e-07, 9.732713e-07, 9.732719e-07, 9.732735e-07, 
    9.732747e-07, 9.732736e-07, 9.732723e-07, 9.732688e-07, 9.732656e-07, 
    9.732622e-07, 9.732613e-07, 9.732573e-07, 9.732606e-07, 9.732552e-07, 
    9.732598e-07, 9.732519e-07, 9.732662e-07, 9.732599e-07, 9.732712e-07, 
    9.732699e-07, 9.732678e-07, 9.732628e-07, 9.732655e-07, 9.732623e-07, 
    9.732693e-07, 9.73273e-07, 9.732739e-07, 9.732756e-07, 9.732738e-07, 
    9.73274e-07, 9.732723e-07, 9.732728e-07, 9.732687e-07, 9.73271e-07, 
    9.732646e-07, 9.732623e-07, 9.732559e-07, 9.732519e-07, 9.732479e-07, 
    9.732461e-07, 9.732455e-07, 9.732453e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  -2.646978e-25, 2.205815e-25, 1.078398e-25, -1.666616e-25, -4.264576e-25, 
    -3.921449e-25, -4.509666e-25, -6.862535e-26, -7.842898e-26, 
    -2.843051e-25, 4.41163e-25, 6.568427e-25, -7.107626e-25, 3.921449e-26, 
    -7.744861e-25, -3.431268e-26, -5.784137e-25, 3.529304e-25, 7.25468e-25, 
    -1.862688e-25, 4.705739e-25, 5.293956e-25, -2.058761e-25, -3.725376e-25, 
    3.039123e-25, 4.509666e-25, 2.254833e-25, 4.901811e-26, -1.519561e-25, 
    -2.254833e-25, 2.156797e-25, 5.882173e-25, -1.421525e-25, 5.391992e-25, 
    -5.882173e-26, 1.539169e-24, -3.578322e-25, -1.220551e-24, -6.274318e-25, 
    -4.705739e-25, -5.588064e-25, 2.745014e-25, 2.745014e-25, -1.372507e-25, 
    3.137159e-25, 6.323336e-25, 6.862535e-26, -2.745014e-25, -2.941087e-26, 
    -1.470543e-26, 1.372507e-25, -1.176435e-24, -7.842898e-26, 2.450905e-26, 
    1.053889e-24, 3.529304e-25, -2.59796e-25, 2.646978e-25, -2.745014e-25, 
    2.156797e-25, 8.578169e-25, 3.431268e-25, -1.372507e-25, -4.41163e-25, 
    2.941087e-26, 3.725376e-25, 1.960724e-25, 2.843051e-25, 3.039123e-25, 
    1.56858e-25, 4.509666e-25, -3.921449e-25, 7.842898e-26, 1.127417e-25, 
    -2.058761e-25, 9.803622e-25, -7.940934e-25, 1.666616e-25, 2.058761e-25, 
    -2.254833e-25, 1.764652e-25, -8.82326e-26, 1.313685e-24, 2.646978e-25, 
    1.960724e-25, 4.607703e-25, -5.588064e-25, -7.548789e-25, 4.41163e-25, 
    -8.725224e-25, -9.509513e-25, 4.901811e-26, -3.774394e-25, 4.803775e-25, 
    -7.744861e-25, -7.646825e-25, 2.59796e-25, -3.676358e-25, 2.205815e-25, 
    3.676358e-25, -4.117521e-25, -4.901811e-27, 0, 5.735119e-25, 
    -3.921449e-26, -2.941087e-26, -4.41163e-25, 3.088141e-25, -8.333079e-25, 
    3.431268e-25, 8.333079e-26, 6.127264e-25, 1.372507e-25, 7.352717e-26, 
    -8.82326e-26, 3.725376e-25, 2.499924e-25, 1.323489e-25, 2.745014e-25, 
    -1.911706e-25, 6.47039e-25, -9.803622e-27, 1.666616e-25, 4.999847e-25, 
    -2.058761e-25, -3.431268e-25, 3.921449e-25, -2.009742e-25, 9.215405e-25, 
    1.127417e-24, 4.803775e-25, 7.352717e-25, 1.372507e-25, 9.85264e-25, 
    -8.82326e-26, 2.058761e-25, -4.607703e-25, 6.47039e-25, 8.03897e-25, 
    -8.382097e-25, 2.352869e-25, -2.205815e-25, 9.901658e-25, 9.803622e-27, 
    1.56858e-25, -3.725376e-25, 4.019485e-25, 3.431268e-25, 8.82326e-26, 
    -1.176435e-25, -2.450905e-26, 3.62734e-25, 2.156797e-25, -8.235043e-25, 
    3.186177e-25, -5.44101e-25, 4.607703e-25, 1.196042e-24, 3.62734e-25, 
    3.921449e-26, -6.666463e-25, -2.254833e-25, -1.176435e-25, 1.078398e-25, 
    -9.803622e-27, -6.862535e-26, 3.039123e-25, 1.862688e-25, 6.862535e-25, 
    3.039123e-25, 3.529304e-25, 3.62734e-25, -1.176435e-25, -5.882173e-26, 
    6.078246e-25, -9.803622e-27, 6.960572e-25, 3.480286e-25, 1.470543e-25, 
    -1.274471e-25, 1.166631e-24, -4.901811e-27, 8.03897e-25, 6.862535e-26, 
    -3.431268e-25, -2.254833e-25, -1.421525e-25, -9.901658e-25, 3.676358e-25, 
    -2.205815e-25, -3.38225e-25, 2.745014e-25, 2.941087e-25, 1.078398e-25, 
    3.62734e-25, 3.137159e-25, 1.127417e-25, -4.999847e-25, 3.823413e-25, 
    4.901811e-26, 1.078398e-25, -6.862535e-26, 2.941087e-25, -5.882173e-26, 
    -1.56858e-25, 1.02938e-25, 2.695996e-25, 1.519561e-25, -3.921449e-26, 
    -1.176435e-25, -1.764652e-25, 1.764652e-25, -3.186177e-25, 9.803622e-26, 
    -1.274471e-25, -3.431268e-26, 1.127417e-24, -3.823413e-25, 2.450906e-25, 
    -2.548942e-25, 2.941087e-25, 8.03897e-25, 1.225453e-25, 1.666616e-25, 
    3.62734e-25, -3.823413e-25, 1.960724e-25, 6.617445e-25, 4.313593e-25, 
    -5.931191e-25, 7.352717e-26, 5.097883e-25, 4.215557e-25, 4.019485e-25, 
    -5.588064e-25, -2.941087e-25, 1.078398e-25, 2.107779e-25, 1.862688e-25, 
    -1.470543e-26, 1.323489e-24, -2.450906e-25, 3.872431e-25, -5.097883e-25, 
    4.313593e-25, -1.470543e-26, -6.47039e-25, -1.470543e-25, 2.941087e-26, 
    2.745014e-25, 1.176435e-25, 4.215557e-25, 3.970467e-25, -8.82326e-26, 
    3.823413e-25, -3.921449e-25, -3.38225e-25, -1.519561e-25, 5.244938e-25, 
    3.725376e-25, -6.274318e-25, 2.450906e-25, 6.568427e-25, -1.764652e-25, 
    0, -9.803622e-26, -3.921449e-26, 4.999847e-25, -3.039123e-25, 
    -4.117521e-25, 4.313593e-25, 5.98021e-25, -4.509666e-25, -5.588064e-25, 
    2.745014e-25, 2.941087e-25, 1.078398e-25, 1.764652e-25, 4.705739e-25, 
    -2.548942e-25, -6.862535e-26, -3.431268e-25, 6.372354e-25, 1.068595e-24, 
    -8.333079e-26, 2.254833e-25, -3.62734e-25, -2.401887e-25, -1.176435e-25, 
    0, 4.215557e-25, 9.313441e-25, -2.352869e-25, 1.323489e-25, 1.470543e-25, 
    6.960572e-25, 5.882173e-26, 4.215557e-25, -2.990105e-25, 4.901811e-27, 
    5.686101e-25, -2.941087e-26, 6.862535e-25, 1.470543e-25, 3.480286e-25, 
    1.088202e-24, -2.59796e-25, -8.82326e-26, -3.62734e-25, 1.323489e-25, 
    1.176435e-25, -1.81367e-25, -2.941087e-26, -4.803775e-25, -5.882173e-26, 
    -1.264667e-24, 6.862535e-26, -1.764652e-25, -2.156797e-25, 2.646978e-25, 
    -3.529304e-25, 3.823413e-25, 4.117521e-25, 1.068595e-24, 1.470543e-26, 
    2.843051e-25, 5.98021e-25, -1.176435e-25, 3.137159e-25, 3.333231e-25, 
    9.901658e-25, 4.901811e-25, 2.941087e-25, -1.323489e-25, -3.62734e-25, 
    2.646978e-25, 4.264576e-25, 1.372507e-25,
  9.436731e-32, 9.436693e-32, 9.436701e-32, 9.436671e-32, 9.436688e-32, 
    9.436668e-32, 9.436723e-32, 9.436692e-32, 9.436712e-32, 9.436728e-32, 
    9.436613e-32, 9.436669e-32, 9.436554e-32, 9.43659e-32, 9.4365e-32, 
    9.436559e-32, 9.436487e-32, 9.436501e-32, 9.43646e-32, 9.436471e-32, 
    9.436418e-32, 9.436454e-32, 9.436391e-32, 9.436427e-32, 9.436421e-32, 
    9.436455e-32, 9.436658e-32, 9.43662e-32, 9.436661e-32, 9.436655e-32, 
    9.436658e-32, 9.436687e-32, 9.436702e-32, 9.436733e-32, 9.436728e-32, 
    9.436705e-32, 9.436652e-32, 9.43667e-32, 9.436625e-32, 9.436626e-32, 
    9.436577e-32, 9.436599e-32, 9.436516e-32, 9.43654e-32, 9.436471e-32, 
    9.436488e-32, 9.436472e-32, 9.436477e-32, 9.436472e-32, 9.436497e-32, 
    9.436486e-32, 9.436508e-32, 9.436595e-32, 9.436569e-32, 9.436645e-32, 
    9.436691e-32, 9.436722e-32, 9.436743e-32, 9.436741e-32, 9.436735e-32, 
    9.436705e-32, 9.436676e-32, 9.436655e-32, 9.436641e-32, 9.436626e-32, 
    9.436584e-32, 9.436561e-32, 9.436511e-32, 9.43652e-32, 9.436505e-32, 
    9.43649e-32, 9.436465e-32, 9.43647e-32, 9.436458e-32, 9.436505e-32, 
    9.436474e-32, 9.436525e-32, 9.436511e-32, 9.436623e-32, 9.436665e-32, 
    9.436684e-32, 9.436699e-32, 9.436738e-32, 9.436711e-32, 9.436722e-32, 
    9.436697e-32, 9.436681e-32, 9.436689e-32, 9.436641e-32, 9.436659e-32, 
    9.43656e-32, 9.436603e-32, 9.436492e-32, 9.436518e-32, 9.436485e-32, 
    9.436502e-32, 9.436473e-32, 9.4365e-32, 9.436454e-32, 9.436445e-32, 
    9.436451e-32, 9.436426e-32, 9.436501e-32, 9.436472e-32, 9.436689e-32, 
    9.436688e-32, 9.436682e-32, 9.436708e-32, 9.436709e-32, 9.436733e-32, 
    9.436712e-32, 9.436703e-32, 9.43668e-32, 9.436666e-32, 9.436654e-32, 
    9.436625e-32, 9.436593e-32, 9.436548e-32, 9.436517e-32, 9.436495e-32, 
    9.436508e-32, 9.436497e-32, 9.43651e-32, 9.436515e-32, 9.436448e-32, 
    9.436486e-32, 9.43643e-32, 9.436433e-32, 9.436458e-32, 9.436433e-32, 
    9.436687e-32, 9.436694e-32, 9.43672e-32, 9.4367e-32, 9.436736e-32, 
    9.436716e-32, 9.436704e-32, 9.436659e-32, 9.436649e-32, 9.436639e-32, 
    9.436621e-32, 9.436598e-32, 9.436557e-32, 9.436521e-32, 9.436489e-32, 
    9.436491e-32, 9.436491e-32, 9.436484e-32, 9.436501e-32, 9.436481e-32, 
    9.436477e-32, 9.436486e-32, 9.436433e-32, 9.436448e-32, 9.436433e-32, 
    9.436443e-32, 9.436692e-32, 9.436679e-32, 9.436686e-32, 9.436674e-32, 
    9.436682e-32, 9.436643e-32, 9.436631e-32, 9.436576e-32, 9.436598e-32, 
    9.436562e-32, 9.436595e-32, 9.436589e-32, 9.436561e-32, 9.436593e-32, 
    9.436524e-32, 9.436571e-32, 9.436483e-32, 9.43653e-32, 9.43648e-32, 
    9.43649e-32, 9.436474e-32, 9.436461e-32, 9.436444e-32, 9.436413e-32, 
    9.43642e-32, 9.436394e-32, 9.436661e-32, 9.436645e-32, 9.436646e-32, 
    9.436629e-32, 9.436617e-32, 9.43659e-32, 9.436547e-32, 9.436563e-32, 
    9.436534e-32, 9.436527e-32, 9.436572e-32, 9.436545e-32, 9.436634e-32, 
    9.436619e-32, 9.436628e-32, 9.436659e-32, 9.436559e-32, 9.436611e-32, 
    9.436516e-32, 9.436544e-32, 9.436463e-32, 9.436503e-32, 9.436424e-32, 
    9.43639e-32, 9.436358e-32, 9.436321e-32, 9.436636e-32, 9.436647e-32, 
    9.436628e-32, 9.436601e-32, 9.436575e-32, 9.436542e-32, 9.436539e-32, 
    9.436532e-32, 9.436517e-32, 9.436502e-32, 9.436531e-32, 9.4365e-32, 
    9.436617e-32, 9.436555e-32, 9.436651e-32, 9.436622e-32, 9.436602e-32, 
    9.436611e-32, 9.436565e-32, 9.436554e-32, 9.436511e-32, 9.436533e-32, 
    9.436398e-32, 9.436458e-32, 9.436293e-32, 9.436339e-32, 9.436651e-32, 
    9.436636e-32, 9.436585e-32, 9.436609e-32, 9.43654e-32, 9.436523e-32, 
    9.436509e-32, 9.436491e-32, 9.43649e-32, 9.436479e-32, 9.436496e-32, 
    9.43648e-32, 9.436542e-32, 9.436514e-32, 9.436591e-32, 9.436572e-32, 
    9.436581e-32, 9.43659e-32, 9.436561e-32, 9.43653e-32, 9.43653e-32, 
    9.43652e-32, 9.436491e-32, 9.43654e-32, 9.436391e-32, 9.436482e-32, 
    9.43662e-32, 9.436592e-32, 9.436588e-32, 9.436599e-32, 9.436524e-32, 
    9.436551e-32, 9.436479e-32, 9.436498e-32, 9.436467e-32, 9.436482e-32, 
    9.436485e-32, 9.436505e-32, 9.436518e-32, 9.43655e-32, 9.436577e-32, 
    9.436597e-32, 9.436592e-32, 9.436569e-32, 9.436528e-32, 9.436489e-32, 
    9.436498e-32, 9.436469e-32, 9.436545e-32, 9.436513e-32, 9.436525e-32, 
    9.436493e-32, 9.436564e-32, 9.436504e-32, 9.436579e-32, 9.436572e-32, 
    9.436552e-32, 9.436511e-32, 9.436502e-32, 9.436492e-32, 9.436498e-32, 
    9.436527e-32, 9.436532e-32, 9.436552e-32, 9.436558e-32, 9.436574e-32, 
    9.436587e-32, 9.436575e-32, 9.436562e-32, 9.436527e-32, 9.436495e-32, 
    9.436461e-32, 9.436452e-32, 9.436412e-32, 9.436445e-32, 9.43639e-32, 
    9.436437e-32, 9.436357e-32, 9.4365e-32, 9.436438e-32, 9.436551e-32, 
    9.436539e-32, 9.436517e-32, 9.436466e-32, 9.436494e-32, 9.436461e-32, 
    9.436532e-32, 9.436569e-32, 9.436578e-32, 9.436596e-32, 9.436578e-32, 
    9.436579e-32, 9.436562e-32, 9.436568e-32, 9.436526e-32, 9.436548e-32, 
    9.436485e-32, 9.436462e-32, 9.436397e-32, 9.436357e-32, 9.436316e-32, 
    9.436299e-32, 9.436293e-32, 9.436291e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.035863e-14, 4.04675e-14, 4.044635e-14, 4.053407e-14, 4.048543e-14, 
    4.054285e-14, 4.038072e-14, 4.04718e-14, 4.041368e-14, 4.036846e-14, 
    4.070406e-14, 4.053799e-14, 4.087643e-14, 4.07707e-14, 4.103612e-14, 
    4.085996e-14, 4.107161e-14, 4.103108e-14, 4.115311e-14, 4.111817e-14, 
    4.127402e-14, 4.116924e-14, 4.135478e-14, 4.124903e-14, 4.126556e-14, 
    4.116577e-14, 4.057147e-14, 4.068339e-14, 4.056482e-14, 4.05808e-14, 
    4.057364e-14, 4.048643e-14, 4.044243e-14, 4.035033e-14, 4.036706e-14, 
    4.043472e-14, 4.058798e-14, 4.0536e-14, 4.066701e-14, 4.066406e-14, 
    4.08097e-14, 4.074406e-14, 4.098854e-14, 4.091914e-14, 4.111963e-14, 
    4.106923e-14, 4.111726e-14, 4.11027e-14, 4.111745e-14, 4.104353e-14, 
    4.10752e-14, 4.101014e-14, 4.075635e-14, 4.0831e-14, 4.060817e-14, 
    4.04739e-14, 4.038471e-14, 4.032135e-14, 4.033032e-14, 4.034738e-14, 
    4.043511e-14, 4.051755e-14, 4.058033e-14, 4.062229e-14, 4.066363e-14, 
    4.078856e-14, 4.08547e-14, 4.100255e-14, 4.097591e-14, 4.102106e-14, 
    4.106422e-14, 4.11366e-14, 4.112469e-14, 4.115656e-14, 4.101989e-14, 
    4.111073e-14, 4.096075e-14, 4.100177e-14, 4.067475e-14, 4.055003e-14, 
    4.049687e-14, 4.045041e-14, 4.03372e-14, 4.041539e-14, 4.038457e-14, 
    4.04579e-14, 4.050445e-14, 4.048143e-14, 4.062344e-14, 4.056825e-14, 
    4.085862e-14, 4.073365e-14, 4.105919e-14, 4.098138e-14, 4.107783e-14, 
    4.102863e-14, 4.111291e-14, 4.103707e-14, 4.116843e-14, 4.119699e-14, 
    4.117747e-14, 4.125249e-14, 4.103285e-14, 4.111725e-14, 4.048078e-14, 
    4.048454e-14, 4.050203e-14, 4.042509e-14, 4.042039e-14, 4.034986e-14, 
    4.041263e-14, 4.043934e-14, 4.050716e-14, 4.054723e-14, 4.058531e-14, 
    4.0669e-14, 4.076237e-14, 4.089282e-14, 4.098643e-14, 4.104914e-14, 
    4.10107e-14, 4.104463e-14, 4.100669e-14, 4.098891e-14, 4.118628e-14, 
    4.107549e-14, 4.12417e-14, 4.123251e-14, 4.115731e-14, 4.123355e-14, 
    4.048717e-14, 4.046557e-14, 4.039049e-14, 4.044925e-14, 4.034218e-14, 
    4.040211e-14, 4.043655e-14, 4.056938e-14, 4.059857e-14, 4.062559e-14, 
    4.067897e-14, 4.074741e-14, 4.086737e-14, 4.097162e-14, 4.106674e-14, 
    4.105977e-14, 4.106222e-14, 4.108345e-14, 4.103085e-14, 4.109208e-14, 
    4.110234e-14, 4.107549e-14, 4.123128e-14, 4.11868e-14, 4.123232e-14, 
    4.120336e-14, 4.047259e-14, 4.050895e-14, 4.04893e-14, 4.052623e-14, 
    4.050021e-14, 4.061585e-14, 4.065049e-14, 4.081248e-14, 4.074606e-14, 
    4.085178e-14, 4.075682e-14, 4.077364e-14, 4.085518e-14, 4.076196e-14, 
    4.096585e-14, 4.082762e-14, 4.108427e-14, 4.094635e-14, 4.109291e-14, 
    4.106633e-14, 4.111034e-14, 4.114974e-14, 4.11993e-14, 4.129065e-14, 
    4.126951e-14, 4.134588e-14, 4.056313e-14, 4.061023e-14, 4.06061e-14, 
    4.065539e-14, 4.069181e-14, 4.077075e-14, 4.089719e-14, 4.084967e-14, 
    4.093693e-14, 4.095443e-14, 4.082187e-14, 4.090325e-14, 4.064175e-14, 
    4.068402e-14, 4.065887e-14, 4.056683e-14, 4.086059e-14, 4.070992e-14, 
    4.098797e-14, 4.09065e-14, 4.114412e-14, 4.102598e-14, 4.125786e-14, 
    4.135677e-14, 4.144987e-14, 4.155842e-14, 4.063594e-14, 4.060395e-14, 
    4.066125e-14, 4.074043e-14, 4.081391e-14, 4.091147e-14, 4.092146e-14, 
    4.093972e-14, 4.098701e-14, 4.102676e-14, 4.094547e-14, 4.103672e-14, 
    4.069378e-14, 4.087367e-14, 4.059183e-14, 4.067675e-14, 4.073577e-14, 
    4.070991e-14, 4.084424e-14, 4.087587e-14, 4.100426e-14, 4.093794e-14, 
    4.133234e-14, 4.115803e-14, 4.164107e-14, 4.150631e-14, 4.059276e-14, 
    4.063585e-14, 4.07856e-14, 4.071438e-14, 4.091799e-14, 4.096802e-14, 
    4.10087e-14, 4.106065e-14, 4.106628e-14, 4.109705e-14, 4.104662e-14, 
    4.109506e-14, 4.091168e-14, 4.099366e-14, 4.076852e-14, 4.082336e-14, 
    4.079814e-14, 4.077046e-14, 4.085587e-14, 4.094674e-14, 4.094872e-14, 
    4.097782e-14, 4.105975e-14, 4.091882e-14, 4.135475e-14, 4.108568e-14, 
    4.06828e-14, 4.076564e-14, 4.077751e-14, 4.074542e-14, 4.096302e-14, 
    4.088423e-14, 4.10963e-14, 4.103903e-14, 4.113286e-14, 4.108624e-14, 
    4.107938e-14, 4.101948e-14, 4.098216e-14, 4.088784e-14, 4.081102e-14, 
    4.075008e-14, 4.076426e-14, 4.083118e-14, 4.095231e-14, 4.106677e-14, 
    4.10417e-14, 4.112573e-14, 4.090324e-14, 4.099656e-14, 4.096051e-14, 
    4.105454e-14, 4.08484e-14, 4.102385e-14, 4.080348e-14, 4.082283e-14, 
    4.088266e-14, 4.100287e-14, 4.10295e-14, 4.105787e-14, 4.104037e-14, 
    4.095539e-14, 4.094147e-14, 4.088122e-14, 4.086456e-14, 4.081863e-14, 
    4.078056e-14, 4.081533e-14, 4.085182e-14, 4.095544e-14, 4.104869e-14, 
    4.115029e-14, 4.117516e-14, 4.129362e-14, 4.119714e-14, 4.135624e-14, 
    4.122092e-14, 4.145509e-14, 4.103406e-14, 4.121701e-14, 4.08854e-14, 
    4.092119e-14, 4.098583e-14, 4.113405e-14, 4.10541e-14, 4.114762e-14, 
    4.094093e-14, 4.083347e-14, 4.08057e-14, 4.075378e-14, 4.080689e-14, 
    4.080257e-14, 4.085336e-14, 4.083704e-14, 4.095888e-14, 4.089345e-14, 
    4.10792e-14, 4.114689e-14, 4.133786e-14, 4.145472e-14, 4.15736e-14, 
    4.162601e-14, 4.164196e-14, 4.164863e-14 ;

 LITR1N_vr =
  5.557581e-05, 5.55756e-05, 5.557564e-05, 5.557547e-05, 5.557557e-05, 
    5.557546e-05, 5.557577e-05, 5.557559e-05, 5.557571e-05, 5.557579e-05, 
    5.557514e-05, 5.557546e-05, 5.557481e-05, 5.557501e-05, 5.55745e-05, 
    5.557484e-05, 5.557443e-05, 5.557451e-05, 5.557427e-05, 5.557434e-05, 
    5.557404e-05, 5.557424e-05, 5.557388e-05, 5.557409e-05, 5.557406e-05, 
    5.557425e-05, 5.55754e-05, 5.557518e-05, 5.557541e-05, 5.557538e-05, 
    5.557539e-05, 5.557557e-05, 5.557565e-05, 5.557583e-05, 5.55758e-05, 
    5.557567e-05, 5.557537e-05, 5.557547e-05, 5.557522e-05, 5.557522e-05, 
    5.557494e-05, 5.557507e-05, 5.557459e-05, 5.557472e-05, 5.557434e-05, 
    5.557443e-05, 5.557434e-05, 5.557437e-05, 5.557434e-05, 5.557448e-05, 
    5.557442e-05, 5.557455e-05, 5.557504e-05, 5.55749e-05, 5.557533e-05, 
    5.557559e-05, 5.557576e-05, 5.557589e-05, 5.557587e-05, 5.557583e-05, 
    5.557566e-05, 5.55755e-05, 5.557538e-05, 5.55753e-05, 5.557522e-05, 
    5.557498e-05, 5.557485e-05, 5.557456e-05, 5.557462e-05, 5.557453e-05, 
    5.557444e-05, 5.55743e-05, 5.557433e-05, 5.557427e-05, 5.557453e-05, 
    5.557435e-05, 5.557464e-05, 5.557456e-05, 5.55752e-05, 5.557544e-05, 
    5.557554e-05, 5.557563e-05, 5.557586e-05, 5.55757e-05, 5.557576e-05, 
    5.557562e-05, 5.557553e-05, 5.557558e-05, 5.55753e-05, 5.55754e-05, 
    5.557484e-05, 5.557508e-05, 5.557446e-05, 5.55746e-05, 5.557442e-05, 
    5.557451e-05, 5.557435e-05, 5.55745e-05, 5.557424e-05, 5.557419e-05, 
    5.557423e-05, 5.557408e-05, 5.557451e-05, 5.557434e-05, 5.557558e-05, 
    5.557557e-05, 5.557554e-05, 5.557569e-05, 5.557569e-05, 5.557583e-05, 
    5.557571e-05, 5.557566e-05, 5.557553e-05, 5.557545e-05, 5.557537e-05, 
    5.557521e-05, 5.557503e-05, 5.557478e-05, 5.557459e-05, 5.557447e-05, 
    5.557455e-05, 5.557448e-05, 5.557456e-05, 5.557459e-05, 5.557421e-05, 
    5.557442e-05, 5.55741e-05, 5.557412e-05, 5.557426e-05, 5.557412e-05, 
    5.557557e-05, 5.557561e-05, 5.557575e-05, 5.557564e-05, 5.557585e-05, 
    5.557573e-05, 5.557566e-05, 5.55754e-05, 5.557535e-05, 5.55753e-05, 
    5.557519e-05, 5.557506e-05, 5.557483e-05, 5.557462e-05, 5.557444e-05, 
    5.557445e-05, 5.557445e-05, 5.557441e-05, 5.557451e-05, 5.557439e-05, 
    5.557437e-05, 5.557442e-05, 5.557412e-05, 5.557421e-05, 5.557412e-05, 
    5.557418e-05, 5.557559e-05, 5.557552e-05, 5.557556e-05, 5.557549e-05, 
    5.557554e-05, 5.557531e-05, 5.557524e-05, 5.557493e-05, 5.557506e-05, 
    5.557486e-05, 5.557504e-05, 5.557501e-05, 5.557485e-05, 5.557503e-05, 
    5.557463e-05, 5.55749e-05, 5.55744e-05, 5.557467e-05, 5.557439e-05, 
    5.557444e-05, 5.557435e-05, 5.557428e-05, 5.557418e-05, 5.5574e-05, 
    5.557405e-05, 5.55739e-05, 5.557542e-05, 5.557532e-05, 5.557533e-05, 
    5.557524e-05, 5.557516e-05, 5.557501e-05, 5.557477e-05, 5.557486e-05, 
    5.557469e-05, 5.557466e-05, 5.557491e-05, 5.557476e-05, 5.557526e-05, 
    5.557518e-05, 5.557523e-05, 5.557541e-05, 5.557484e-05, 5.557513e-05, 
    5.557459e-05, 5.557475e-05, 5.557429e-05, 5.557452e-05, 5.557407e-05, 
    5.557388e-05, 5.55737e-05, 5.557349e-05, 5.557527e-05, 5.557534e-05, 
    5.557523e-05, 5.557507e-05, 5.557493e-05, 5.557474e-05, 5.557472e-05, 
    5.557468e-05, 5.557459e-05, 5.557452e-05, 5.557467e-05, 5.55745e-05, 
    5.557516e-05, 5.557482e-05, 5.557536e-05, 5.557519e-05, 5.557508e-05, 
    5.557513e-05, 5.557487e-05, 5.557481e-05, 5.557456e-05, 5.557469e-05, 
    5.557392e-05, 5.557426e-05, 5.557333e-05, 5.557359e-05, 5.557536e-05, 
    5.557527e-05, 5.557498e-05, 5.557512e-05, 5.557473e-05, 5.557463e-05, 
    5.557455e-05, 5.557445e-05, 5.557444e-05, 5.557438e-05, 5.557448e-05, 
    5.557439e-05, 5.557474e-05, 5.557458e-05, 5.557502e-05, 5.557491e-05, 
    5.557496e-05, 5.557502e-05, 5.557485e-05, 5.557467e-05, 5.557467e-05, 
    5.557461e-05, 5.557445e-05, 5.557473e-05, 5.557388e-05, 5.55744e-05, 
    5.557518e-05, 5.557502e-05, 5.5575e-05, 5.557506e-05, 5.557464e-05, 
    5.557479e-05, 5.557438e-05, 5.557449e-05, 5.557431e-05, 5.55744e-05, 
    5.557442e-05, 5.557453e-05, 5.55746e-05, 5.557479e-05, 5.557494e-05, 
    5.557505e-05, 5.557503e-05, 5.55749e-05, 5.557466e-05, 5.557444e-05, 
    5.557449e-05, 5.557432e-05, 5.557476e-05, 5.557458e-05, 5.557464e-05, 
    5.557446e-05, 5.557486e-05, 5.557452e-05, 5.557495e-05, 5.557491e-05, 
    5.55748e-05, 5.557456e-05, 5.557451e-05, 5.557446e-05, 5.557449e-05, 
    5.557466e-05, 5.557468e-05, 5.55748e-05, 5.557483e-05, 5.557492e-05, 
    5.557499e-05, 5.557493e-05, 5.557486e-05, 5.557466e-05, 5.557447e-05, 
    5.557428e-05, 5.557423e-05, 5.5574e-05, 5.557419e-05, 5.557388e-05, 
    5.557414e-05, 5.557369e-05, 5.55745e-05, 5.557415e-05, 5.557479e-05, 
    5.557472e-05, 5.55746e-05, 5.557431e-05, 5.557446e-05, 5.557428e-05, 
    5.557468e-05, 5.557489e-05, 5.557495e-05, 5.557504e-05, 5.557494e-05, 
    5.557495e-05, 5.557485e-05, 5.557488e-05, 5.557465e-05, 5.557478e-05, 
    5.557442e-05, 5.557428e-05, 5.557391e-05, 5.557369e-05, 5.557346e-05, 
    5.557336e-05, 5.557332e-05, 5.557331e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  6.994304e-13, 7.013172e-13, 7.009506e-13, 7.02471e-13, 7.01628e-13, 
    7.026231e-13, 6.998134e-13, 7.013917e-13, 7.003845e-13, 6.996007e-13, 
    7.05417e-13, 7.025388e-13, 7.084041e-13, 7.065718e-13, 7.111716e-13, 
    7.081188e-13, 7.117866e-13, 7.110842e-13, 7.131991e-13, 7.125936e-13, 
    7.152945e-13, 7.134786e-13, 7.166941e-13, 7.148614e-13, 7.15148e-13, 
    7.134185e-13, 7.03119e-13, 7.050587e-13, 7.030038e-13, 7.032806e-13, 
    7.031566e-13, 7.016452e-13, 7.008827e-13, 6.992865e-13, 6.995765e-13, 
    7.00749e-13, 7.034051e-13, 7.025043e-13, 7.047748e-13, 7.047236e-13, 
    7.072476e-13, 7.0611e-13, 7.10347e-13, 7.091442e-13, 7.126189e-13, 
    7.117455e-13, 7.125777e-13, 7.123255e-13, 7.12581e-13, 7.112999e-13, 
    7.118489e-13, 7.107214e-13, 7.06323e-13, 7.076167e-13, 7.037551e-13, 
    7.014282e-13, 6.998825e-13, 6.987845e-13, 6.989397e-13, 6.992355e-13, 
    7.007559e-13, 7.021847e-13, 7.032726e-13, 7.039998e-13, 7.047162e-13, 
    7.068813e-13, 7.080275e-13, 7.105898e-13, 7.101281e-13, 7.109106e-13, 
    7.116586e-13, 7.129129e-13, 7.127066e-13, 7.132588e-13, 7.108904e-13, 
    7.124646e-13, 7.098654e-13, 7.105763e-13, 7.049088e-13, 7.027475e-13, 
    7.018262e-13, 7.01021e-13, 6.99059e-13, 7.004141e-13, 6.9988e-13, 
    7.011508e-13, 7.019575e-13, 7.015587e-13, 7.040197e-13, 7.030633e-13, 
    7.080954e-13, 7.059297e-13, 7.115714e-13, 7.10223e-13, 7.118945e-13, 
    7.110418e-13, 7.125024e-13, 7.11188e-13, 7.134645e-13, 7.139596e-13, 
    7.136212e-13, 7.149213e-13, 7.11115e-13, 7.125775e-13, 7.015474e-13, 
    7.016124e-13, 7.019157e-13, 7.005822e-13, 7.005007e-13, 6.992785e-13, 
    7.003663e-13, 7.008292e-13, 7.020044e-13, 7.026989e-13, 7.033589e-13, 
    7.048093e-13, 7.064273e-13, 7.08688e-13, 7.103104e-13, 7.113972e-13, 
    7.10731e-13, 7.113191e-13, 7.106616e-13, 7.103534e-13, 7.13774e-13, 
    7.118539e-13, 7.147344e-13, 7.145752e-13, 7.132719e-13, 7.145932e-13, 
    7.016581e-13, 7.012837e-13, 6.999826e-13, 7.010009e-13, 6.991454e-13, 
    7.00184e-13, 7.007807e-13, 7.030828e-13, 7.035887e-13, 7.04057e-13, 
    7.049821e-13, 7.061683e-13, 7.082471e-13, 7.100538e-13, 7.117022e-13, 
    7.115815e-13, 7.11624e-13, 7.119918e-13, 7.110802e-13, 7.121414e-13, 
    7.123193e-13, 7.118539e-13, 7.145539e-13, 7.13783e-13, 7.145718e-13, 
    7.1407e-13, 7.014055e-13, 7.020355e-13, 7.01695e-13, 7.023351e-13, 
    7.01884e-13, 7.038881e-13, 7.044885e-13, 7.072959e-13, 7.061448e-13, 
    7.07977e-13, 7.063312e-13, 7.066227e-13, 7.080358e-13, 7.064203e-13, 
    7.099538e-13, 7.075583e-13, 7.120061e-13, 7.096158e-13, 7.121558e-13, 
    7.11695e-13, 7.124579e-13, 7.131407e-13, 7.139996e-13, 7.155827e-13, 
    7.152164e-13, 7.165398e-13, 7.029745e-13, 7.037907e-13, 7.037192e-13, 
    7.045733e-13, 7.052046e-13, 7.065726e-13, 7.08764e-13, 7.079404e-13, 
    7.094526e-13, 7.097558e-13, 7.074586e-13, 7.08869e-13, 7.04337e-13, 
    7.050696e-13, 7.046338e-13, 7.030386e-13, 7.081296e-13, 7.055185e-13, 
    7.103371e-13, 7.089253e-13, 7.130433e-13, 7.109959e-13, 7.150145e-13, 
    7.167285e-13, 7.183419e-13, 7.202233e-13, 7.042364e-13, 7.03682e-13, 
    7.04675e-13, 7.060472e-13, 7.073205e-13, 7.090114e-13, 7.091846e-13, 
    7.09501e-13, 7.103205e-13, 7.110093e-13, 7.096006e-13, 7.11182e-13, 
    7.052387e-13, 7.083563e-13, 7.034719e-13, 7.049436e-13, 7.059665e-13, 
    7.055183e-13, 7.078463e-13, 7.083944e-13, 7.106194e-13, 7.0947e-13, 
    7.163053e-13, 7.132842e-13, 7.216556e-13, 7.193201e-13, 7.034881e-13, 
    7.042347e-13, 7.0683e-13, 7.055957e-13, 7.091244e-13, 7.099914e-13, 
    7.106965e-13, 7.115967e-13, 7.116942e-13, 7.122274e-13, 7.113536e-13, 
    7.121931e-13, 7.09015e-13, 7.104358e-13, 7.065341e-13, 7.074844e-13, 
    7.070474e-13, 7.065677e-13, 7.080478e-13, 7.096227e-13, 7.09657e-13, 
    7.101612e-13, 7.115811e-13, 7.091387e-13, 7.166936e-13, 7.120304e-13, 
    7.050484e-13, 7.06484e-13, 7.066898e-13, 7.061337e-13, 7.099048e-13, 
    7.085392e-13, 7.122145e-13, 7.11222e-13, 7.128481e-13, 7.120402e-13, 
    7.119213e-13, 7.108832e-13, 7.102364e-13, 7.086017e-13, 7.072705e-13, 
    7.062144e-13, 7.064601e-13, 7.0762e-13, 7.097192e-13, 7.117028e-13, 
    7.112683e-13, 7.127246e-13, 7.088688e-13, 7.104861e-13, 7.098612e-13, 
    7.114908e-13, 7.079183e-13, 7.10959e-13, 7.071399e-13, 7.074753e-13, 
    7.085121e-13, 7.105953e-13, 7.110569e-13, 7.115484e-13, 7.112453e-13, 
    7.097725e-13, 7.095313e-13, 7.084871e-13, 7.081984e-13, 7.074023e-13, 
    7.067427e-13, 7.073452e-13, 7.079776e-13, 7.097734e-13, 7.113894e-13, 
    7.131503e-13, 7.135812e-13, 7.156341e-13, 7.139622e-13, 7.167194e-13, 
    7.143742e-13, 7.184325e-13, 7.11136e-13, 7.143065e-13, 7.085595e-13, 
    7.091798e-13, 7.103e-13, 7.128689e-13, 7.114832e-13, 7.131039e-13, 
    7.09522e-13, 7.076597e-13, 7.071783e-13, 7.062786e-13, 7.071989e-13, 
    7.071241e-13, 7.080042e-13, 7.077215e-13, 7.09833e-13, 7.086992e-13, 
    7.119182e-13, 7.130913e-13, 7.164009e-13, 7.184261e-13, 7.204863e-13, 
    7.213946e-13, 7.21671e-13, 7.217866e-13 ;

 LITR2C =
  1.9396e-05, 1.939598e-05, 1.939598e-05, 1.939597e-05, 1.939597e-05, 
    1.939596e-05, 1.939599e-05, 1.939598e-05, 1.939599e-05, 1.939599e-05, 
    1.939593e-05, 1.939597e-05, 1.939591e-05, 1.939592e-05, 1.939588e-05, 
    1.939591e-05, 1.939587e-05, 1.939588e-05, 1.939585e-05, 1.939586e-05, 
    1.939583e-05, 1.939585e-05, 1.939582e-05, 1.939584e-05, 1.939583e-05, 
    1.939585e-05, 1.939596e-05, 1.939594e-05, 1.939596e-05, 1.939596e-05, 
    1.939596e-05, 1.939597e-05, 1.939598e-05, 1.9396e-05, 1.9396e-05, 
    1.939598e-05, 1.939596e-05, 1.939597e-05, 1.939594e-05, 1.939594e-05, 
    1.939592e-05, 1.939593e-05, 1.939588e-05, 1.93959e-05, 1.939586e-05, 
    1.939587e-05, 1.939586e-05, 1.939586e-05, 1.939586e-05, 1.939587e-05, 
    1.939587e-05, 1.939588e-05, 1.939593e-05, 1.939591e-05, 1.939595e-05, 
    1.939598e-05, 1.939599e-05, 1.9396e-05, 1.9396e-05, 1.9396e-05, 
    1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939595e-05, 1.939594e-05, 
    1.939592e-05, 1.939591e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939587e-05, 1.939586e-05, 1.939586e-05, 1.939585e-05, 1.939588e-05, 
    1.939586e-05, 1.939589e-05, 1.939588e-05, 1.939594e-05, 1.939596e-05, 
    1.939597e-05, 1.939598e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.939598e-05, 1.939597e-05, 1.939597e-05, 1.939595e-05, 1.939596e-05, 
    1.939591e-05, 1.939593e-05, 1.939587e-05, 1.939589e-05, 1.939587e-05, 
    1.939588e-05, 1.939586e-05, 1.939588e-05, 1.939585e-05, 1.939585e-05, 
    1.939585e-05, 1.939584e-05, 1.939588e-05, 1.939586e-05, 1.939597e-05, 
    1.939597e-05, 1.939597e-05, 1.939599e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939596e-05, 
    1.939594e-05, 1.939593e-05, 1.93959e-05, 1.939589e-05, 1.939587e-05, 
    1.939588e-05, 1.939587e-05, 1.939588e-05, 1.939588e-05, 1.939585e-05, 
    1.939587e-05, 1.939584e-05, 1.939584e-05, 1.939585e-05, 1.939584e-05, 
    1.939597e-05, 1.939598e-05, 1.939599e-05, 1.939598e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939596e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939587e-05, 1.939587e-05, 1.939588e-05, 1.939587e-05, 
    1.939586e-05, 1.939587e-05, 1.939584e-05, 1.939585e-05, 1.939584e-05, 
    1.939585e-05, 1.939598e-05, 1.939597e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939595e-05, 1.939595e-05, 1.939592e-05, 1.939593e-05, 
    1.939591e-05, 1.939593e-05, 1.939592e-05, 1.939591e-05, 1.939593e-05, 
    1.939589e-05, 1.939591e-05, 1.939587e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939586e-05, 1.939586e-05, 1.939585e-05, 1.939583e-05, 
    1.939583e-05, 1.939582e-05, 1.939596e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939594e-05, 1.939592e-05, 1.93959e-05, 1.939591e-05, 
    1.939589e-05, 1.939589e-05, 1.939591e-05, 1.93959e-05, 1.939595e-05, 
    1.939594e-05, 1.939594e-05, 1.939596e-05, 1.939591e-05, 1.939593e-05, 
    1.939589e-05, 1.93959e-05, 1.939586e-05, 1.939588e-05, 1.939584e-05, 
    1.939582e-05, 1.93958e-05, 1.939578e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 1.93959e-05, 
    1.939589e-05, 1.939589e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939594e-05, 1.939591e-05, 1.939596e-05, 1.939594e-05, 1.939593e-05, 
    1.939593e-05, 1.939591e-05, 1.939591e-05, 1.939588e-05, 1.939589e-05, 
    1.939582e-05, 1.939585e-05, 1.939577e-05, 1.939579e-05, 1.939595e-05, 
    1.939595e-05, 1.939592e-05, 1.939593e-05, 1.93959e-05, 1.939589e-05, 
    1.939588e-05, 1.939587e-05, 1.939587e-05, 1.939587e-05, 1.939587e-05, 
    1.939587e-05, 1.93959e-05, 1.939588e-05, 1.939592e-05, 1.939591e-05, 
    1.939592e-05, 1.939592e-05, 1.939591e-05, 1.939589e-05, 1.939589e-05, 
    1.939589e-05, 1.939587e-05, 1.93959e-05, 1.939582e-05, 1.939587e-05, 
    1.939594e-05, 1.939592e-05, 1.939592e-05, 1.939593e-05, 1.939589e-05, 
    1.93959e-05, 1.939587e-05, 1.939588e-05, 1.939586e-05, 1.939587e-05, 
    1.939587e-05, 1.939588e-05, 1.939589e-05, 1.93959e-05, 1.939592e-05, 
    1.939593e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939586e-05, 1.93959e-05, 1.939588e-05, 1.939589e-05, 
    1.939587e-05, 1.939591e-05, 1.939588e-05, 1.939592e-05, 1.939591e-05, 
    1.93959e-05, 1.939588e-05, 1.939588e-05, 1.939587e-05, 1.939587e-05, 
    1.939589e-05, 1.939589e-05, 1.93959e-05, 1.939591e-05, 1.939591e-05, 
    1.939592e-05, 1.939592e-05, 1.939591e-05, 1.939589e-05, 1.939587e-05, 
    1.939586e-05, 1.939585e-05, 1.939583e-05, 1.939585e-05, 1.939582e-05, 
    1.939584e-05, 1.93958e-05, 1.939588e-05, 1.939584e-05, 1.93959e-05, 
    1.93959e-05, 1.939589e-05, 1.939586e-05, 1.939587e-05, 1.939586e-05, 
    1.939589e-05, 1.939591e-05, 1.939592e-05, 1.939593e-05, 1.939592e-05, 
    1.939592e-05, 1.939591e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939587e-05, 1.939586e-05, 1.939582e-05, 1.93958e-05, 1.939578e-05, 
    1.939577e-05, 1.939577e-05, 1.939577e-05 ;

 LITR2C_TO_SOIL1C =
  1.065062e-13, 1.067938e-13, 1.067379e-13, 1.069696e-13, 1.068412e-13, 
    1.069928e-13, 1.065646e-13, 1.068051e-13, 1.066516e-13, 1.065321e-13, 
    1.074187e-13, 1.0698e-13, 1.07874e-13, 1.075947e-13, 1.082958e-13, 
    1.078305e-13, 1.083896e-13, 1.082825e-13, 1.086049e-13, 1.085126e-13, 
    1.089243e-13, 1.086475e-13, 1.091376e-13, 1.088583e-13, 1.089019e-13, 
    1.086383e-13, 1.070684e-13, 1.073641e-13, 1.070509e-13, 1.070931e-13, 
    1.070741e-13, 1.068438e-13, 1.067275e-13, 1.064843e-13, 1.065285e-13, 
    1.067072e-13, 1.07112e-13, 1.069747e-13, 1.073208e-13, 1.07313e-13, 
    1.076977e-13, 1.075243e-13, 1.081701e-13, 1.079868e-13, 1.085164e-13, 
    1.083833e-13, 1.085102e-13, 1.084717e-13, 1.085107e-13, 1.083154e-13, 
    1.083991e-13, 1.082272e-13, 1.075568e-13, 1.07754e-13, 1.071654e-13, 
    1.068107e-13, 1.065751e-13, 1.064077e-13, 1.064314e-13, 1.064765e-13, 
    1.067082e-13, 1.06926e-13, 1.070918e-13, 1.072027e-13, 1.073119e-13, 
    1.076419e-13, 1.078166e-13, 1.082072e-13, 1.081368e-13, 1.082561e-13, 
    1.083701e-13, 1.085613e-13, 1.085298e-13, 1.08614e-13, 1.08253e-13, 
    1.084929e-13, 1.080967e-13, 1.082051e-13, 1.073412e-13, 1.070118e-13, 
    1.068714e-13, 1.067486e-13, 1.064496e-13, 1.066561e-13, 1.065747e-13, 
    1.067684e-13, 1.068914e-13, 1.068306e-13, 1.072057e-13, 1.070599e-13, 
    1.078269e-13, 1.074968e-13, 1.083568e-13, 1.081512e-13, 1.08406e-13, 
    1.082761e-13, 1.084987e-13, 1.082983e-13, 1.086453e-13, 1.087208e-13, 
    1.086692e-13, 1.088674e-13, 1.082872e-13, 1.085101e-13, 1.068289e-13, 
    1.068388e-13, 1.06885e-13, 1.066818e-13, 1.066693e-13, 1.06483e-13, 
    1.066488e-13, 1.067194e-13, 1.068985e-13, 1.070044e-13, 1.07105e-13, 
    1.073261e-13, 1.075727e-13, 1.079173e-13, 1.081646e-13, 1.083302e-13, 
    1.082287e-13, 1.083183e-13, 1.082181e-13, 1.081711e-13, 1.086925e-13, 
    1.083998e-13, 1.088389e-13, 1.088146e-13, 1.08616e-13, 1.088174e-13, 
    1.068457e-13, 1.067887e-13, 1.065903e-13, 1.067456e-13, 1.064627e-13, 
    1.066211e-13, 1.06712e-13, 1.070629e-13, 1.0714e-13, 1.072114e-13, 
    1.073524e-13, 1.075332e-13, 1.078501e-13, 1.081255e-13, 1.083767e-13, 
    1.083583e-13, 1.083648e-13, 1.084209e-13, 1.082819e-13, 1.084437e-13, 
    1.084708e-13, 1.083998e-13, 1.088114e-13, 1.086939e-13, 1.088141e-13, 
    1.087376e-13, 1.068072e-13, 1.069033e-13, 1.068514e-13, 1.069489e-13, 
    1.068802e-13, 1.071856e-13, 1.072772e-13, 1.077051e-13, 1.075296e-13, 
    1.078089e-13, 1.07558e-13, 1.076025e-13, 1.078179e-13, 1.075716e-13, 
    1.081102e-13, 1.077451e-13, 1.08423e-13, 1.080587e-13, 1.084459e-13, 
    1.083756e-13, 1.084919e-13, 1.08596e-13, 1.087269e-13, 1.089682e-13, 
    1.089124e-13, 1.091141e-13, 1.070464e-13, 1.071708e-13, 1.071599e-13, 
    1.072901e-13, 1.073863e-13, 1.075948e-13, 1.079289e-13, 1.078033e-13, 
    1.080338e-13, 1.0808e-13, 1.077299e-13, 1.079449e-13, 1.072541e-13, 
    1.073657e-13, 1.072993e-13, 1.070562e-13, 1.078322e-13, 1.074342e-13, 
    1.081686e-13, 1.079534e-13, 1.085811e-13, 1.082691e-13, 1.088816e-13, 
    1.091429e-13, 1.093888e-13, 1.096756e-13, 1.072387e-13, 1.071542e-13, 
    1.073056e-13, 1.075147e-13, 1.077088e-13, 1.079666e-13, 1.07993e-13, 
    1.080412e-13, 1.081661e-13, 1.082711e-13, 1.080564e-13, 1.082974e-13, 
    1.073915e-13, 1.078667e-13, 1.071222e-13, 1.073465e-13, 1.075024e-13, 
    1.074341e-13, 1.07789e-13, 1.078725e-13, 1.082117e-13, 1.080365e-13, 
    1.090784e-13, 1.086179e-13, 1.098939e-13, 1.095379e-13, 1.071247e-13, 
    1.072385e-13, 1.076341e-13, 1.074459e-13, 1.079838e-13, 1.081159e-13, 
    1.082234e-13, 1.083606e-13, 1.083755e-13, 1.084568e-13, 1.083236e-13, 
    1.084515e-13, 1.079671e-13, 1.081837e-13, 1.07589e-13, 1.077338e-13, 
    1.076672e-13, 1.075941e-13, 1.078197e-13, 1.080597e-13, 1.08065e-13, 
    1.081418e-13, 1.083583e-13, 1.07986e-13, 1.091375e-13, 1.084267e-13, 
    1.073625e-13, 1.075813e-13, 1.076127e-13, 1.075279e-13, 1.081027e-13, 
    1.078946e-13, 1.084548e-13, 1.083035e-13, 1.085514e-13, 1.084282e-13, 
    1.084101e-13, 1.082519e-13, 1.081533e-13, 1.079041e-13, 1.077012e-13, 
    1.075402e-13, 1.075777e-13, 1.077545e-13, 1.080744e-13, 1.083768e-13, 
    1.083106e-13, 1.085326e-13, 1.079448e-13, 1.081913e-13, 1.080961e-13, 
    1.083445e-13, 1.078e-13, 1.082634e-13, 1.076813e-13, 1.077324e-13, 
    1.078905e-13, 1.08208e-13, 1.082784e-13, 1.083533e-13, 1.083071e-13, 
    1.080826e-13, 1.080458e-13, 1.078866e-13, 1.078426e-13, 1.077213e-13, 
    1.076208e-13, 1.077126e-13, 1.07809e-13, 1.080827e-13, 1.08329e-13, 
    1.085975e-13, 1.086631e-13, 1.089761e-13, 1.087212e-13, 1.091415e-13, 
    1.08784e-13, 1.094026e-13, 1.082904e-13, 1.087737e-13, 1.078977e-13, 
    1.079922e-13, 1.08163e-13, 1.085545e-13, 1.083433e-13, 1.085904e-13, 
    1.080444e-13, 1.077605e-13, 1.076872e-13, 1.0755e-13, 1.076903e-13, 
    1.076789e-13, 1.078131e-13, 1.077699e-13, 1.080918e-13, 1.07919e-13, 
    1.084096e-13, 1.085885e-13, 1.090929e-13, 1.094016e-13, 1.097157e-13, 
    1.098541e-13, 1.098963e-13, 1.099139e-13 ;

 LITR2C_vr =
  0.001107531, 0.00110753, 0.001107531, 0.00110753, 0.00110753, 0.00110753, 
    0.001107531, 0.00110753, 0.001107531, 0.001107531, 0.001107528, 
    0.00110753, 0.001107526, 0.001107527, 0.001107525, 0.001107526, 
    0.001107524, 0.001107525, 0.001107523, 0.001107524, 0.001107522, 
    0.001107523, 0.001107521, 0.001107522, 0.001107522, 0.001107523, 
    0.001107529, 0.001107528, 0.001107529, 0.001107529, 0.001107529, 
    0.00110753, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107529, 0.00110753, 0.001107528, 0.001107528, 0.001107527, 
    0.001107528, 0.001107525, 0.001107526, 0.001107524, 0.001107524, 
    0.001107524, 0.001107524, 0.001107524, 0.001107524, 0.001107524, 
    0.001107525, 0.001107527, 0.001107527, 0.001107529, 0.00110753, 
    0.001107531, 0.001107532, 0.001107532, 0.001107532, 0.001107531, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107527, 
    0.001107526, 0.001107525, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107523, 0.001107525, 0.001107524, 
    0.001107525, 0.001107525, 0.001107528, 0.00110753, 0.00110753, 
    0.001107531, 0.001107532, 0.001107531, 0.001107531, 0.00110753, 
    0.00110753, 0.00110753, 0.001107529, 0.001107529, 0.001107526, 
    0.001107528, 0.001107524, 0.001107525, 0.001107524, 0.001107525, 
    0.001107524, 0.001107525, 0.001107523, 0.001107523, 0.001107523, 
    0.001107522, 0.001107525, 0.001107524, 0.00110753, 0.00110753, 
    0.00110753, 0.001107531, 0.001107531, 0.001107532, 0.001107531, 
    0.001107531, 0.00110753, 0.00110753, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107525, 0.001107524, 0.001107525, 
    0.001107524, 0.001107525, 0.001107525, 0.001107523, 0.001107524, 
    0.001107523, 0.001107523, 0.001107523, 0.001107523, 0.00110753, 
    0.00110753, 0.001107531, 0.001107531, 0.001107532, 0.001107531, 
    0.001107531, 0.001107529, 0.001107529, 0.001107529, 0.001107528, 
    0.001107528, 0.001107526, 0.001107525, 0.001107524, 0.001107524, 
    0.001107524, 0.001107524, 0.001107525, 0.001107524, 0.001107524, 
    0.001107524, 0.001107523, 0.001107523, 0.001107523, 0.001107523, 
    0.00110753, 0.00110753, 0.00110753, 0.00110753, 0.00110753, 0.001107529, 
    0.001107529, 0.001107527, 0.001107528, 0.001107526, 0.001107527, 
    0.001107527, 0.001107526, 0.001107527, 0.001107525, 0.001107527, 
    0.001107524, 0.001107526, 0.001107524, 0.001107524, 0.001107524, 
    0.001107523, 0.001107523, 0.001107522, 0.001107522, 0.001107521, 
    0.001107529, 0.001107529, 0.001107529, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107525, 
    0.001107527, 0.001107526, 0.001107529, 0.001107528, 0.001107528, 
    0.001107529, 0.001107526, 0.001107528, 0.001107525, 0.001107526, 
    0.001107523, 0.001107525, 0.001107522, 0.001107521, 0.00110752, 
    0.001107519, 0.001107529, 0.001107529, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107525, 
    0.001107525, 0.001107526, 0.001107525, 0.001107528, 0.001107526, 
    0.001107529, 0.001107528, 0.001107528, 0.001107528, 0.001107527, 
    0.001107526, 0.001107525, 0.001107526, 0.001107522, 0.001107523, 
    0.001107518, 0.00110752, 0.001107529, 0.001107529, 0.001107527, 
    0.001107528, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107524, 0.001107524, 0.001107526, 
    0.001107525, 0.001107527, 0.001107527, 0.001107527, 0.001107527, 
    0.001107526, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107526, 0.001107521, 0.001107524, 0.001107528, 0.001107527, 
    0.001107527, 0.001107528, 0.001107525, 0.001107526, 0.001107524, 
    0.001107524, 0.001107524, 0.001107524, 0.001107524, 0.001107525, 
    0.001107525, 0.001107526, 0.001107527, 0.001107528, 0.001107527, 
    0.001107527, 0.001107525, 0.001107524, 0.001107524, 0.001107524, 
    0.001107526, 0.001107525, 0.001107525, 0.001107524, 0.001107526, 
    0.001107525, 0.001107527, 0.001107527, 0.001107526, 0.001107525, 
    0.001107525, 0.001107524, 0.001107524, 0.001107525, 0.001107526, 
    0.001107526, 0.001107526, 0.001107527, 0.001107527, 0.001107527, 
    0.001107526, 0.001107525, 0.001107524, 0.001107523, 0.001107523, 
    0.001107522, 0.001107523, 0.001107521, 0.001107523, 0.00110752, 
    0.001107525, 0.001107523, 0.001107526, 0.001107526, 0.001107525, 
    0.001107524, 0.001107524, 0.001107523, 0.001107526, 0.001107527, 
    0.001107527, 0.001107528, 0.001107527, 0.001107527, 0.001107526, 
    0.001107527, 0.001107525, 0.001107526, 0.001107524, 0.001107523, 
    0.001107521, 0.00110752, 0.001107519, 0.001107519, 0.001107518, 
    0.001107518,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684263e-07, 2.684261e-07, 2.684261e-07, 2.684259e-07, 2.68426e-07, 
    2.684259e-07, 2.684263e-07, 2.684261e-07, 2.684262e-07, 2.684263e-07, 
    2.684255e-07, 2.684259e-07, 2.684251e-07, 2.684253e-07, 2.684247e-07, 
    2.684251e-07, 2.684246e-07, 2.684247e-07, 2.684244e-07, 2.684245e-07, 
    2.684241e-07, 2.684243e-07, 2.684239e-07, 2.684241e-07, 2.684241e-07, 
    2.684243e-07, 2.684258e-07, 2.684255e-07, 2.684258e-07, 2.684258e-07, 
    2.684258e-07, 2.68426e-07, 2.684261e-07, 2.684264e-07, 2.684263e-07, 
    2.684262e-07, 2.684258e-07, 2.684259e-07, 2.684256e-07, 2.684256e-07, 
    2.684252e-07, 2.684254e-07, 2.684248e-07, 2.684249e-07, 2.684245e-07, 
    2.684246e-07, 2.684245e-07, 2.684245e-07, 2.684245e-07, 2.684247e-07, 
    2.684246e-07, 2.684247e-07, 2.684254e-07, 2.684252e-07, 2.684257e-07, 
    2.68426e-07, 2.684263e-07, 2.684264e-07, 2.684264e-07, 2.684264e-07, 
    2.684262e-07, 2.68426e-07, 2.684258e-07, 2.684257e-07, 2.684256e-07, 
    2.684253e-07, 2.684251e-07, 2.684247e-07, 2.684248e-07, 2.684247e-07, 
    2.684246e-07, 2.684244e-07, 2.684245e-07, 2.684244e-07, 2.684247e-07, 
    2.684245e-07, 2.684249e-07, 2.684247e-07, 2.684256e-07, 2.684259e-07, 
    2.68426e-07, 2.684261e-07, 2.684264e-07, 2.684262e-07, 2.684263e-07, 
    2.684261e-07, 2.68426e-07, 2.68426e-07, 2.684257e-07, 2.684258e-07, 
    2.684251e-07, 2.684254e-07, 2.684246e-07, 2.684248e-07, 2.684246e-07, 
    2.684247e-07, 2.684245e-07, 2.684247e-07, 2.684243e-07, 2.684243e-07, 
    2.684243e-07, 2.684241e-07, 2.684247e-07, 2.684245e-07, 2.68426e-07, 
    2.68426e-07, 2.68426e-07, 2.684262e-07, 2.684262e-07, 2.684264e-07, 
    2.684262e-07, 2.684261e-07, 2.68426e-07, 2.684259e-07, 2.684258e-07, 
    2.684256e-07, 2.684253e-07, 2.68425e-07, 2.684248e-07, 2.684246e-07, 
    2.684247e-07, 2.684247e-07, 2.684247e-07, 2.684248e-07, 2.684243e-07, 
    2.684246e-07, 2.684241e-07, 2.684242e-07, 2.684244e-07, 2.684242e-07, 
    2.68426e-07, 2.684261e-07, 2.684263e-07, 2.684261e-07, 2.684264e-07, 
    2.684262e-07, 2.684262e-07, 2.684258e-07, 2.684257e-07, 2.684257e-07, 
    2.684255e-07, 2.684254e-07, 2.684251e-07, 2.684248e-07, 2.684246e-07, 
    2.684246e-07, 2.684246e-07, 2.684245e-07, 2.684247e-07, 2.684245e-07, 
    2.684245e-07, 2.684246e-07, 2.684242e-07, 2.684243e-07, 2.684242e-07, 
    2.684243e-07, 2.68426e-07, 2.68426e-07, 2.68426e-07, 2.684259e-07, 
    2.68426e-07, 2.684257e-07, 2.684256e-07, 2.684252e-07, 2.684254e-07, 
    2.684251e-07, 2.684254e-07, 2.684253e-07, 2.684251e-07, 2.684253e-07, 
    2.684248e-07, 2.684252e-07, 2.684245e-07, 2.684249e-07, 2.684245e-07, 
    2.684246e-07, 2.684245e-07, 2.684244e-07, 2.684243e-07, 2.68424e-07, 
    2.684241e-07, 2.684239e-07, 2.684259e-07, 2.684257e-07, 2.684257e-07, 
    2.684256e-07, 2.684255e-07, 2.684253e-07, 2.68425e-07, 2.684251e-07, 
    2.684249e-07, 2.684249e-07, 2.684252e-07, 2.68425e-07, 2.684257e-07, 
    2.684255e-07, 2.684256e-07, 2.684258e-07, 2.684251e-07, 2.684255e-07, 
    2.684248e-07, 2.68425e-07, 2.684244e-07, 2.684247e-07, 2.684241e-07, 
    2.684239e-07, 2.684236e-07, 2.684234e-07, 2.684257e-07, 2.684257e-07, 
    2.684256e-07, 2.684254e-07, 2.684252e-07, 2.68425e-07, 2.684249e-07, 
    2.684249e-07, 2.684248e-07, 2.684247e-07, 2.684249e-07, 2.684247e-07, 
    2.684255e-07, 2.684251e-07, 2.684258e-07, 2.684256e-07, 2.684254e-07, 
    2.684255e-07, 2.684251e-07, 2.684251e-07, 2.684247e-07, 2.684249e-07, 
    2.684239e-07, 2.684244e-07, 2.684232e-07, 2.684235e-07, 2.684258e-07, 
    2.684257e-07, 2.684253e-07, 2.684255e-07, 2.68425e-07, 2.684248e-07, 
    2.684247e-07, 2.684246e-07, 2.684246e-07, 2.684245e-07, 2.684246e-07, 
    2.684245e-07, 2.68425e-07, 2.684248e-07, 2.684253e-07, 2.684252e-07, 
    2.684253e-07, 2.684253e-07, 2.684251e-07, 2.684249e-07, 2.684249e-07, 
    2.684248e-07, 2.684246e-07, 2.68425e-07, 2.684239e-07, 2.684245e-07, 
    2.684255e-07, 2.684253e-07, 2.684253e-07, 2.684254e-07, 2.684249e-07, 
    2.684251e-07, 2.684245e-07, 2.684247e-07, 2.684244e-07, 2.684245e-07, 
    2.684246e-07, 2.684247e-07, 2.684248e-07, 2.68425e-07, 2.684252e-07, 
    2.684254e-07, 2.684253e-07, 2.684252e-07, 2.684249e-07, 2.684246e-07, 
    2.684247e-07, 2.684244e-07, 2.68425e-07, 2.684248e-07, 2.684249e-07, 
    2.684246e-07, 2.684251e-07, 2.684247e-07, 2.684253e-07, 2.684252e-07, 
    2.684251e-07, 2.684247e-07, 2.684247e-07, 2.684246e-07, 2.684247e-07, 
    2.684249e-07, 2.684249e-07, 2.684251e-07, 2.684251e-07, 2.684252e-07, 
    2.684253e-07, 2.684252e-07, 2.684251e-07, 2.684249e-07, 2.684246e-07, 
    2.684244e-07, 2.684243e-07, 2.68424e-07, 2.684243e-07, 2.684239e-07, 
    2.684242e-07, 2.684236e-07, 2.684247e-07, 2.684242e-07, 2.68425e-07, 
    2.684249e-07, 2.684248e-07, 2.684244e-07, 2.684246e-07, 2.684244e-07, 
    2.684249e-07, 2.684252e-07, 2.684252e-07, 2.684254e-07, 2.684252e-07, 
    2.684253e-07, 2.684251e-07, 2.684252e-07, 2.684249e-07, 2.68425e-07, 
    2.684246e-07, 2.684244e-07, 2.684239e-07, 2.684236e-07, 2.684233e-07, 
    2.684232e-07, 2.684232e-07, 2.684232e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -5.882173e-26, -2.59796e-25, -9.803622e-26, -2.695996e-26, 1.960724e-26, 
    -1.29898e-25, -2.450906e-27, -1.347998e-25, -2.941087e-26, -9.313441e-26, 
    -6.372354e-26, 6.862535e-26, -1.617598e-25, 3.921449e-26, 1.004871e-25, 
    -2.034252e-25, 2.695996e-26, -1.495052e-25, 9.068351e-26, -7.597807e-26, 
    -2.941087e-26, -6.617445e-26, -7.597807e-26, -8.333079e-26, 
    -1.960724e-26, 0, -4.65672e-26, -8.087988e-26, 1.519561e-25, 
    2.377378e-25, -3.431268e-26, 5.146902e-26, 9.313441e-26, 3.676358e-26, 
    -2.450905e-26, -6.372354e-26, 8.333079e-26, 1.789161e-25, 6.372354e-26, 
    -7.842898e-26, 1.176435e-25, 7.107626e-26, 1.838179e-25, 7.107626e-26, 
    9.803622e-26, 1.960724e-26, 1.642107e-25, -7.352717e-26, 1.666616e-25, 
    -1.274471e-25, -1.617598e-25, -1.495052e-25, 1.519561e-25, -9.313441e-26, 
    1.176435e-25, 2.107779e-25, 1.960724e-26, -8.82326e-26, -1.715634e-26, 
    -1.004871e-25, -2.08327e-25, -2.450906e-27, -2.377378e-25, -3.676358e-26, 
    -1.911706e-25, -6.372354e-26, 1.29898e-25, -1.176435e-25, 1.862688e-25, 
    6.617445e-26, -1.740143e-25, -1.102908e-25, -6.862535e-26, 2.450906e-27, 
    -4.41163e-26, -1.642107e-25, 2.181306e-25, 1.470543e-26, 1.530638e-41, 
    2.548942e-25, -1.470543e-26, -1.911706e-25, 2.401887e-25, -4.901811e-26, 
    1.838179e-25, 5.637083e-26, -2.08327e-25, 1.249962e-25, 2.695996e-26, 
    -6.372354e-26, -1.764652e-25, -3.431268e-26, -1.715634e-25, 8.087988e-26, 
    -1.862688e-25, -3.676358e-26, -2.941087e-25, 1.642107e-25, -1.789161e-25, 
    -7.352717e-26, 7.352717e-27, -2.401887e-25, 1.960724e-26, -3.357741e-25, 
    -9.558531e-26, 4.65672e-26, -1.960724e-26, -5.637083e-26, -7.842898e-26, 
    -1.960724e-26, 3.186177e-26, -2.181306e-25, 1.151926e-25, -1.151926e-25, 
    -1.862688e-25, 8.82326e-26, 4.166539e-26, 1.530638e-41, -2.695996e-25, 
    2.695996e-25, -4.41163e-26, 1.593089e-25, 5.637083e-26, -1.911706e-25, 
    -1.960724e-25, -4.41163e-26, 4.41163e-26, 8.087988e-26, -2.08327e-25, 
    5.146902e-26, 3.676358e-26, 3.406759e-25, 1.102908e-25, 7.352717e-26, 
    -1.151926e-25, 1.127417e-25, -1.323489e-25, 3.161668e-25, 2.450905e-26, 
    9.558531e-26, 5.882173e-26, -5.882173e-26, 3.921449e-26, -1.691125e-25, 
    -8.82326e-26, 3.921449e-26, 3.186177e-26, -1.715634e-26, 2.941087e-25, 
    1.200944e-25, 6.617445e-26, 1.862688e-25, 4.41163e-26, -9.803622e-27, 
    -1.421525e-25, 1.789161e-25, 1.446034e-25, 8.087988e-26, 1.470543e-26, 
    9.068351e-26, 2.622469e-25, -1.54407e-25, 2.107779e-25, -1.470543e-26, 
    -3.259704e-25, 1.02938e-25, -1.397016e-25, 6.372354e-26, 1.715634e-26, 
    -7.352717e-27, -8.578169e-26, 1.053889e-25, -5.391992e-26, -7.107626e-26, 
    1.691125e-25, -1.004871e-25, 2.279342e-25, -1.495052e-25, -1.691125e-25, 
    3.186177e-26, 1.617598e-25, -1.29898e-25, 2.009742e-25, -2.156797e-25, 
    6.372354e-26, 1.519561e-25, -1.642107e-25, -2.450906e-27, -9.803622e-27, 
    -1.666616e-25, 7.107626e-26, 1.078398e-25, -4.166539e-26, 1.249962e-25, 
    3.186177e-26, -1.225453e-26, -5.882173e-26, -6.127264e-26, 4.41163e-26, 
    -3.431268e-26, -1.127417e-25, 6.862535e-26, 2.695996e-26, -1.715634e-26, 
    1.530638e-41, -7.107626e-26, -1.519561e-25, 8.578169e-26, 1.02938e-25, 
    -1.666616e-25, -1.249962e-25, 1.617598e-25, -8.333079e-26, 8.333079e-26, 
    7.352717e-27, -1.372507e-25, -2.205815e-25, 1.862688e-25, 7.107626e-26, 
    -1.642107e-25, -1.078398e-25, -7.352717e-27, -7.842898e-26, 
    -6.617445e-26, -3.676358e-26, -1.838179e-25, -8.087988e-26, 
    -5.882173e-26, 1.053889e-25, -1.470543e-25, 4.901811e-26, 5.882173e-26, 
    1.225453e-25, -1.225453e-25, 1.911706e-25, -5.391992e-26, -1.764652e-25, 
    1.151926e-25, 1.200944e-25, -2.867559e-25, 8.333079e-26, -1.29898e-25, 
    -1.960724e-26, -3.676358e-26, 4.901811e-27, -9.803622e-27, 1.838179e-25, 
    -3.186177e-26, -2.352869e-25, -2.695996e-26, -4.901811e-26, 
    -1.470543e-25, 1.764652e-25, -1.764652e-25, 7.352717e-27, -4.901811e-27, 
    -9.068351e-26, 2.107779e-25, -2.622469e-25, -8.333079e-26, -1.54407e-25, 
    4.166539e-26, -2.965596e-25, -9.558531e-26, 7.352717e-27, 1.347998e-25, 
    -1.960724e-26, 5.637083e-26, -2.08327e-25, -1.102908e-25, 1.176435e-25, 
    -9.313441e-26, 2.08327e-25, 1.470543e-26, 5.882173e-26, 1.519561e-25, 
    2.695996e-26, -1.960724e-26, -2.695996e-26, -3.186177e-26, 4.41163e-26, 
    -1.446034e-25, -2.009742e-25, -1.936215e-25, -5.391992e-26, 
    -2.303851e-25, 2.450905e-26, 1.225453e-25, 1.176435e-25, -8.578169e-26, 
    -2.450906e-27, 9.313441e-26, 2.941087e-26, -1.347998e-25, -8.333079e-26, 
    4.901811e-26, -9.803622e-26, -2.499924e-25, -7.842898e-26, -7.842898e-26, 
    -2.450905e-26, -1.764652e-25, 1.985233e-25, -7.352717e-26, 1.274471e-25, 
    2.450905e-26, -1.985233e-25, -1.666616e-25, 8.087988e-26, -1.54407e-25, 
    -5.146902e-26, 3.431268e-26, 4.166539e-26, 3.921449e-26, 2.941087e-25, 
    -2.524433e-25, -2.205815e-26, 1.936215e-25, -2.181306e-25, 2.205815e-26, 
    -2.450905e-26, -2.254833e-25, 1.446034e-25, 3.921449e-26, -3.431268e-25, 
    1.127417e-25, 1.151926e-25, -5.882173e-26, -1.960724e-26, 1.470543e-26, 
    -4.901811e-26, 0, -8.82326e-26, 4.166539e-26, 1.397016e-25, 1.838179e-25, 
    2.107779e-25, -7.597807e-26,
  2.67625e-32, 2.676247e-32, 2.676247e-32, 2.676245e-32, 2.676247e-32, 
    2.676245e-32, 2.676249e-32, 2.676247e-32, 2.676248e-32, 2.676249e-32, 
    2.676241e-32, 2.676245e-32, 2.676237e-32, 2.676239e-32, 2.676233e-32, 
    2.676237e-32, 2.676232e-32, 2.676233e-32, 2.67623e-32, 2.676231e-32, 
    2.676227e-32, 2.676229e-32, 2.676225e-32, 2.676227e-32, 2.676227e-32, 
    2.676229e-32, 2.676244e-32, 2.676242e-32, 2.676244e-32, 2.676244e-32, 
    2.676244e-32, 2.676247e-32, 2.676248e-32, 2.67625e-32, 2.676249e-32, 
    2.676248e-32, 2.676244e-32, 2.676245e-32, 2.676242e-32, 2.676242e-32, 
    2.676238e-32, 2.67624e-32, 2.676234e-32, 2.676236e-32, 2.676231e-32, 
    2.676232e-32, 2.676231e-32, 2.676231e-32, 2.676231e-32, 2.676233e-32, 
    2.676232e-32, 2.676233e-32, 2.67624e-32, 2.676238e-32, 2.676244e-32, 
    2.676247e-32, 2.676249e-32, 2.676251e-32, 2.67625e-32, 2.67625e-32, 
    2.676248e-32, 2.676246e-32, 2.676244e-32, 2.676243e-32, 2.676242e-32, 
    2.676239e-32, 2.676237e-32, 2.676234e-32, 2.676234e-32, 2.676233e-32, 
    2.676232e-32, 2.67623e-32, 2.676231e-32, 2.67623e-32, 2.676233e-32, 
    2.676231e-32, 2.676235e-32, 2.676234e-32, 2.676242e-32, 2.676245e-32, 
    2.676246e-32, 2.676247e-32, 2.67625e-32, 2.676248e-32, 2.676249e-32, 
    2.676247e-32, 2.676246e-32, 2.676247e-32, 2.676243e-32, 2.676244e-32, 
    2.676237e-32, 2.67624e-32, 2.676232e-32, 2.676234e-32, 2.676232e-32, 
    2.676233e-32, 2.676231e-32, 2.676233e-32, 2.676229e-32, 2.676229e-32, 
    2.676229e-32, 2.676227e-32, 2.676233e-32, 2.676231e-32, 2.676247e-32, 
    2.676247e-32, 2.676246e-32, 2.676248e-32, 2.676248e-32, 2.67625e-32, 
    2.676248e-32, 2.676248e-32, 2.676246e-32, 2.676245e-32, 2.676244e-32, 
    2.676242e-32, 2.676239e-32, 2.676236e-32, 2.676234e-32, 2.676232e-32, 
    2.676233e-32, 2.676233e-32, 2.676234e-32, 2.676234e-32, 2.676229e-32, 
    2.676232e-32, 2.676228e-32, 2.676228e-32, 2.67623e-32, 2.676228e-32, 
    2.676247e-32, 2.676247e-32, 2.676249e-32, 2.676247e-32, 2.67625e-32, 
    2.676249e-32, 2.676248e-32, 2.676244e-32, 2.676244e-32, 2.676243e-32, 
    2.676242e-32, 2.67624e-32, 2.676237e-32, 2.676234e-32, 2.676232e-32, 
    2.676232e-32, 2.676232e-32, 2.676232e-32, 2.676233e-32, 2.676232e-32, 
    2.676231e-32, 2.676232e-32, 2.676228e-32, 2.676229e-32, 2.676228e-32, 
    2.676229e-32, 2.676247e-32, 2.676246e-32, 2.676247e-32, 2.676245e-32, 
    2.676246e-32, 2.676243e-32, 2.676242e-32, 2.676238e-32, 2.67624e-32, 
    2.676237e-32, 2.67624e-32, 2.676239e-32, 2.676237e-32, 2.67624e-32, 
    2.676234e-32, 2.676238e-32, 2.676232e-32, 2.676235e-32, 2.676231e-32, 
    2.676232e-32, 2.676231e-32, 2.67623e-32, 2.676229e-32, 2.676227e-32, 
    2.676227e-32, 2.676225e-32, 2.676244e-32, 2.676243e-32, 2.676244e-32, 
    2.676242e-32, 2.676241e-32, 2.676239e-32, 2.676236e-32, 2.676237e-32, 
    2.676235e-32, 2.676235e-32, 2.676238e-32, 2.676236e-32, 2.676243e-32, 
    2.676242e-32, 2.676242e-32, 2.676244e-32, 2.676237e-32, 2.676241e-32, 
    2.676234e-32, 2.676236e-32, 2.67623e-32, 2.676233e-32, 2.676227e-32, 
    2.676225e-32, 2.676222e-32, 2.67622e-32, 2.676243e-32, 2.676244e-32, 
    2.676242e-32, 2.67624e-32, 2.676238e-32, 2.676236e-32, 2.676236e-32, 
    2.676235e-32, 2.676234e-32, 2.676233e-32, 2.676235e-32, 2.676233e-32, 
    2.676241e-32, 2.676237e-32, 2.676244e-32, 2.676242e-32, 2.67624e-32, 
    2.676241e-32, 2.676238e-32, 2.676237e-32, 2.676234e-32, 2.676235e-32, 
    2.676225e-32, 2.67623e-32, 2.676218e-32, 2.676221e-32, 2.676244e-32, 
    2.676243e-32, 2.676239e-32, 2.676241e-32, 2.676236e-32, 2.676234e-32, 
    2.676234e-32, 2.676232e-32, 2.676232e-32, 2.676231e-32, 2.676232e-32, 
    2.676231e-32, 2.676236e-32, 2.676234e-32, 2.676239e-32, 2.676238e-32, 
    2.676239e-32, 2.676239e-32, 2.676237e-32, 2.676235e-32, 2.676235e-32, 
    2.676234e-32, 2.676232e-32, 2.676236e-32, 2.676225e-32, 2.676232e-32, 
    2.676242e-32, 2.676239e-32, 2.676239e-32, 2.67624e-32, 2.676234e-32, 
    2.676237e-32, 2.676231e-32, 2.676233e-32, 2.67623e-32, 2.676232e-32, 
    2.676232e-32, 2.676233e-32, 2.676234e-32, 2.676237e-32, 2.676238e-32, 
    2.67624e-32, 2.676239e-32, 2.676238e-32, 2.676235e-32, 2.676232e-32, 
    2.676233e-32, 2.676231e-32, 2.676236e-32, 2.676234e-32, 2.676235e-32, 
    2.676232e-32, 2.676237e-32, 2.676233e-32, 2.676239e-32, 2.676238e-32, 
    2.676237e-32, 2.676234e-32, 2.676233e-32, 2.676232e-32, 2.676233e-32, 
    2.676235e-32, 2.676235e-32, 2.676237e-32, 2.676237e-32, 2.676238e-32, 
    2.676239e-32, 2.676238e-32, 2.676237e-32, 2.676235e-32, 2.676232e-32, 
    2.67623e-32, 2.676229e-32, 2.676226e-32, 2.676229e-32, 2.676225e-32, 
    2.676228e-32, 2.676222e-32, 2.676233e-32, 2.676228e-32, 2.676237e-32, 
    2.676236e-32, 2.676234e-32, 2.67623e-32, 2.676232e-32, 2.67623e-32, 
    2.676235e-32, 2.676238e-32, 2.676239e-32, 2.67624e-32, 2.676239e-32, 
    2.676239e-32, 2.676237e-32, 2.676238e-32, 2.676235e-32, 2.676236e-32, 
    2.676232e-32, 2.67623e-32, 2.676225e-32, 2.676222e-32, 2.676219e-32, 
    2.676218e-32, 2.676218e-32, 2.676217e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  2.947935e-15, 2.955894e-15, 2.954348e-15, 2.960762e-15, 2.957206e-15, 
    2.961404e-15, 2.94955e-15, 2.956209e-15, 2.95196e-15, 2.948653e-15, 
    2.973191e-15, 2.961049e-15, 2.985794e-15, 2.978063e-15, 2.99747e-15, 
    2.98459e-15, 3.000064e-15, 2.997101e-15, 3.006024e-15, 3.003469e-15, 
    3.014864e-15, 3.007203e-15, 3.020769e-15, 3.013037e-15, 3.014246e-15, 
    3.006949e-15, 2.963496e-15, 2.97168e-15, 2.963011e-15, 2.964178e-15, 
    2.963655e-15, 2.957279e-15, 2.954062e-15, 2.947328e-15, 2.948551e-15, 
    2.953498e-15, 2.964703e-15, 2.960903e-15, 2.970482e-15, 2.970266e-15, 
    2.980915e-15, 2.976115e-15, 2.993991e-15, 2.988916e-15, 3.003576e-15, 
    2.999891e-15, 3.003402e-15, 3.002338e-15, 3.003416e-15, 2.998011e-15, 
    3.000327e-15, 2.99557e-15, 2.977014e-15, 2.982472e-15, 2.96618e-15, 
    2.956363e-15, 2.949842e-15, 2.94521e-15, 2.945865e-15, 2.947113e-15, 
    2.953527e-15, 2.959555e-15, 2.964144e-15, 2.967213e-15, 2.970235e-15, 
    2.979369e-15, 2.984205e-15, 2.995015e-15, 2.993067e-15, 2.996369e-15, 
    2.999524e-15, 3.004816e-15, 3.003946e-15, 3.006276e-15, 2.996283e-15, 
    3.002925e-15, 2.991959e-15, 2.994958e-15, 2.971048e-15, 2.961929e-15, 
    2.958042e-15, 2.954645e-15, 2.946368e-15, 2.952085e-15, 2.949831e-15, 
    2.955193e-15, 2.958596e-15, 2.956913e-15, 2.967297e-15, 2.963261e-15, 
    2.984491e-15, 2.975354e-15, 2.999156e-15, 2.993467e-15, 3.00052e-15, 
    2.996922e-15, 3.003084e-15, 2.997539e-15, 3.007143e-15, 3.009232e-15, 
    3.007805e-15, 3.01329e-15, 2.997231e-15, 3.003401e-15, 2.956866e-15, 
    2.95714e-15, 2.95842e-15, 2.952794e-15, 2.95245e-15, 2.947294e-15, 
    2.951883e-15, 2.953836e-15, 2.958794e-15, 2.961724e-15, 2.964509e-15, 
    2.970628e-15, 2.977454e-15, 2.986992e-15, 2.993836e-15, 2.998421e-15, 
    2.995611e-15, 2.998092e-15, 2.995318e-15, 2.994018e-15, 3.008449e-15, 
    3.000348e-15, 3.012501e-15, 3.011829e-15, 3.006331e-15, 3.011905e-15, 
    2.957333e-15, 2.955754e-15, 2.950264e-15, 2.95456e-15, 2.946732e-15, 
    2.951114e-15, 2.953632e-15, 2.963344e-15, 2.965478e-15, 2.967454e-15, 
    2.971356e-15, 2.976361e-15, 2.985131e-15, 2.992754e-15, 2.999708e-15, 
    2.999199e-15, 2.999378e-15, 3.00093e-15, 2.997084e-15, 3.001561e-15, 
    3.002311e-15, 3.000348e-15, 3.011739e-15, 3.008487e-15, 3.011815e-15, 
    3.009698e-15, 2.956267e-15, 2.958925e-15, 2.957489e-15, 2.960189e-15, 
    2.958286e-15, 2.966741e-15, 2.969274e-15, 2.981118e-15, 2.976262e-15, 
    2.983992e-15, 2.977048e-15, 2.978278e-15, 2.98424e-15, 2.977424e-15, 
    2.992332e-15, 2.982225e-15, 3.00099e-15, 2.990906e-15, 3.001622e-15, 
    2.999678e-15, 3.002897e-15, 3.005777e-15, 3.009401e-15, 3.01608e-15, 
    3.014534e-15, 3.020118e-15, 2.962887e-15, 2.96633e-15, 2.966029e-15, 
    2.969632e-15, 2.972295e-15, 2.978067e-15, 2.987312e-15, 2.983837e-15, 
    2.990217e-15, 2.991497e-15, 2.981805e-15, 2.987755e-15, 2.968635e-15, 
    2.971726e-15, 2.969887e-15, 2.963157e-15, 2.984636e-15, 2.97362e-15, 
    2.993949e-15, 2.987993e-15, 3.005366e-15, 2.996729e-15, 3.013683e-15, 
    3.020914e-15, 3.027721e-15, 3.035659e-15, 2.968211e-15, 2.965871e-15, 
    2.970061e-15, 2.97585e-15, 2.981222e-15, 2.988356e-15, 2.989086e-15, 
    2.990421e-15, 2.993879e-15, 2.996785e-15, 2.990842e-15, 2.997514e-15, 
    2.972439e-15, 2.985592e-15, 2.964985e-15, 2.971194e-15, 2.97551e-15, 
    2.973619e-15, 2.98344e-15, 2.985753e-15, 2.99514e-15, 2.990291e-15, 
    3.019129e-15, 3.006383e-15, 3.041702e-15, 3.031849e-15, 2.965053e-15, 
    2.968203e-15, 2.979153e-15, 2.973945e-15, 2.988833e-15, 2.99249e-15, 
    2.995465e-15, 2.999263e-15, 2.999675e-15, 3.001924e-15, 2.998237e-15, 
    3.001779e-15, 2.988371e-15, 2.994365e-15, 2.977904e-15, 2.981913e-15, 
    2.98007e-15, 2.978046e-15, 2.98429e-15, 2.990935e-15, 2.99108e-15, 
    2.993207e-15, 2.999197e-15, 2.988893e-15, 3.020767e-15, 3.001093e-15, 
    2.971636e-15, 2.977693e-15, 2.978561e-15, 2.976215e-15, 2.992125e-15, 
    2.986364e-15, 3.00187e-15, 2.997682e-15, 3.004543e-15, 3.001134e-15, 
    3.000633e-15, 2.996253e-15, 2.993524e-15, 2.986628e-15, 2.981011e-15, 
    2.976556e-15, 2.977592e-15, 2.982486e-15, 2.991342e-15, 2.999711e-15, 
    2.997877e-15, 3.004022e-15, 2.987754e-15, 2.994577e-15, 2.991941e-15, 
    2.998816e-15, 2.983744e-15, 2.996573e-15, 2.98046e-15, 2.981875e-15, 
    2.98625e-15, 2.995038e-15, 2.996986e-15, 2.99906e-15, 2.997781e-15, 
    2.991567e-15, 2.99055e-15, 2.986144e-15, 2.984926e-15, 2.981567e-15, 
    2.978784e-15, 2.981326e-15, 2.983994e-15, 2.991571e-15, 2.998389e-15, 
    3.005818e-15, 3.007636e-15, 3.016297e-15, 3.009243e-15, 3.020876e-15, 
    3.010981e-15, 3.028103e-15, 2.997319e-15, 3.010696e-15, 2.986449e-15, 
    2.989066e-15, 2.993792e-15, 3.00463e-15, 2.998784e-15, 3.005622e-15, 
    2.99051e-15, 2.982653e-15, 2.980622e-15, 2.976826e-15, 2.980709e-15, 
    2.980393e-15, 2.984107e-15, 2.982914e-15, 2.991822e-15, 2.987038e-15, 
    3.000619e-15, 3.005569e-15, 3.019532e-15, 3.028077e-15, 3.036769e-15, 
    3.040601e-15, 3.041767e-15, 3.042255e-15 ;

 LITR2N_vr =
  1.532742e-05, 1.532741e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532742e-05, 1.53274e-05, 1.532741e-05, 1.532742e-05, 
    1.532737e-05, 1.53274e-05, 1.532735e-05, 1.532736e-05, 1.532732e-05, 
    1.532735e-05, 1.532732e-05, 1.532733e-05, 1.532731e-05, 1.532731e-05, 
    1.532729e-05, 1.532731e-05, 1.532728e-05, 1.53273e-05, 1.532729e-05, 
    1.532731e-05, 1.532739e-05, 1.532738e-05, 1.532739e-05, 1.532739e-05, 
    1.532739e-05, 1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.532739e-05, 1.53274e-05, 1.532738e-05, 1.532738e-05, 
    1.532736e-05, 1.532737e-05, 1.532733e-05, 1.532734e-05, 1.532731e-05, 
    1.532732e-05, 1.532731e-05, 1.532732e-05, 1.532731e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.532736e-05, 1.532735e-05, 1.532739e-05, 
    1.53274e-05, 1.532742e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 1.532738e-05, 
    1.532736e-05, 1.532735e-05, 1.532733e-05, 1.532733e-05, 1.532733e-05, 
    1.532732e-05, 1.532731e-05, 1.532731e-05, 1.532731e-05, 1.532733e-05, 
    1.532732e-05, 1.532734e-05, 1.532733e-05, 1.532738e-05, 1.532739e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.53274e-05, 1.532738e-05, 1.532739e-05, 
    1.532735e-05, 1.532737e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532733e-05, 1.532731e-05, 1.532732e-05, 1.532731e-05, 1.53273e-05, 
    1.53273e-05, 1.53273e-05, 1.532733e-05, 1.532731e-05, 1.53274e-05, 
    1.53274e-05, 1.53274e-05, 1.532741e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 1.532739e-05, 
    1.532738e-05, 1.532736e-05, 1.532735e-05, 1.532733e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532733e-05, 1.53273e-05, 
    1.532732e-05, 1.53273e-05, 1.53273e-05, 1.532731e-05, 1.53273e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532732e-05, 1.53273e-05, 1.53273e-05, 1.53273e-05, 
    1.53273e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532738e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532735e-05, 1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532736e-05, 
    1.532734e-05, 1.532736e-05, 1.532732e-05, 1.532734e-05, 1.532732e-05, 
    1.532732e-05, 1.532732e-05, 1.532731e-05, 1.53273e-05, 1.532729e-05, 
    1.532729e-05, 1.532728e-05, 1.532739e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 
    1.532734e-05, 1.532734e-05, 1.532736e-05, 1.532734e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532739e-05, 1.532735e-05, 1.532737e-05, 
    1.532733e-05, 1.532734e-05, 1.532731e-05, 1.532733e-05, 1.532729e-05, 
    1.532728e-05, 1.532727e-05, 1.532725e-05, 1.532738e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532733e-05, 1.532734e-05, 1.532732e-05, 
    1.532737e-05, 1.532735e-05, 1.532739e-05, 1.532738e-05, 1.532737e-05, 
    1.532737e-05, 1.532735e-05, 1.532735e-05, 1.532733e-05, 1.532734e-05, 
    1.532728e-05, 1.532731e-05, 1.532724e-05, 1.532726e-05, 1.532739e-05, 
    1.532738e-05, 1.532736e-05, 1.532737e-05, 1.532734e-05, 1.532734e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 
    1.532732e-05, 1.532734e-05, 1.532733e-05, 1.532736e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532734e-05, 
    1.532733e-05, 1.532732e-05, 1.532734e-05, 1.532728e-05, 1.532732e-05, 
    1.532738e-05, 1.532736e-05, 1.532736e-05, 1.532737e-05, 1.532734e-05, 
    1.532735e-05, 1.532732e-05, 1.532732e-05, 1.532731e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.532733e-05, 1.532735e-05, 1.532736e-05, 
    1.532737e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532732e-05, 
    1.532732e-05, 1.532731e-05, 1.532734e-05, 1.532733e-05, 1.532734e-05, 
    1.532732e-05, 1.532735e-05, 1.532733e-05, 1.532736e-05, 1.532736e-05, 
    1.532735e-05, 1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532732e-05, 
    1.532734e-05, 1.532734e-05, 1.532735e-05, 1.532735e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532732e-05, 
    1.532731e-05, 1.532731e-05, 1.532729e-05, 1.53273e-05, 1.532728e-05, 
    1.53273e-05, 1.532727e-05, 1.532733e-05, 1.53273e-05, 1.532735e-05, 
    1.532734e-05, 1.532733e-05, 1.532731e-05, 1.532732e-05, 1.532731e-05, 
    1.532734e-05, 1.532735e-05, 1.532736e-05, 1.532736e-05, 1.532736e-05, 
    1.532736e-05, 1.532735e-05, 1.532735e-05, 1.532734e-05, 1.532735e-05, 
    1.532732e-05, 1.532731e-05, 1.532728e-05, 1.532727e-05, 1.532725e-05, 
    1.532724e-05, 1.532724e-05, 1.532724e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.065062e-13, 1.067938e-13, 1.067379e-13, 1.069696e-13, 1.068412e-13, 
    1.069928e-13, 1.065646e-13, 1.068051e-13, 1.066516e-13, 1.065321e-13, 
    1.074187e-13, 1.0698e-13, 1.07874e-13, 1.075947e-13, 1.082958e-13, 
    1.078305e-13, 1.083896e-13, 1.082825e-13, 1.086049e-13, 1.085126e-13, 
    1.089243e-13, 1.086475e-13, 1.091376e-13, 1.088583e-13, 1.089019e-13, 
    1.086383e-13, 1.070684e-13, 1.073641e-13, 1.070509e-13, 1.070931e-13, 
    1.070741e-13, 1.068438e-13, 1.067275e-13, 1.064843e-13, 1.065285e-13, 
    1.067072e-13, 1.07112e-13, 1.069747e-13, 1.073208e-13, 1.07313e-13, 
    1.076977e-13, 1.075243e-13, 1.081701e-13, 1.079868e-13, 1.085164e-13, 
    1.083833e-13, 1.085102e-13, 1.084717e-13, 1.085107e-13, 1.083154e-13, 
    1.083991e-13, 1.082272e-13, 1.075568e-13, 1.07754e-13, 1.071654e-13, 
    1.068107e-13, 1.065751e-13, 1.064077e-13, 1.064314e-13, 1.064765e-13, 
    1.067082e-13, 1.06926e-13, 1.070918e-13, 1.072027e-13, 1.073119e-13, 
    1.076419e-13, 1.078166e-13, 1.082072e-13, 1.081368e-13, 1.082561e-13, 
    1.083701e-13, 1.085613e-13, 1.085298e-13, 1.08614e-13, 1.08253e-13, 
    1.084929e-13, 1.080967e-13, 1.082051e-13, 1.073412e-13, 1.070118e-13, 
    1.068714e-13, 1.067486e-13, 1.064496e-13, 1.066561e-13, 1.065747e-13, 
    1.067684e-13, 1.068914e-13, 1.068306e-13, 1.072057e-13, 1.070599e-13, 
    1.078269e-13, 1.074968e-13, 1.083568e-13, 1.081512e-13, 1.08406e-13, 
    1.082761e-13, 1.084987e-13, 1.082983e-13, 1.086453e-13, 1.087208e-13, 
    1.086692e-13, 1.088674e-13, 1.082872e-13, 1.085101e-13, 1.068289e-13, 
    1.068388e-13, 1.06885e-13, 1.066818e-13, 1.066693e-13, 1.06483e-13, 
    1.066488e-13, 1.067194e-13, 1.068985e-13, 1.070044e-13, 1.07105e-13, 
    1.073261e-13, 1.075727e-13, 1.079173e-13, 1.081646e-13, 1.083302e-13, 
    1.082287e-13, 1.083183e-13, 1.082181e-13, 1.081711e-13, 1.086925e-13, 
    1.083998e-13, 1.088389e-13, 1.088146e-13, 1.08616e-13, 1.088174e-13, 
    1.068457e-13, 1.067887e-13, 1.065903e-13, 1.067456e-13, 1.064627e-13, 
    1.066211e-13, 1.06712e-13, 1.070629e-13, 1.0714e-13, 1.072114e-13, 
    1.073524e-13, 1.075332e-13, 1.078501e-13, 1.081255e-13, 1.083767e-13, 
    1.083583e-13, 1.083648e-13, 1.084209e-13, 1.082819e-13, 1.084437e-13, 
    1.084708e-13, 1.083998e-13, 1.088114e-13, 1.086939e-13, 1.088141e-13, 
    1.087376e-13, 1.068072e-13, 1.069033e-13, 1.068514e-13, 1.069489e-13, 
    1.068802e-13, 1.071856e-13, 1.072772e-13, 1.077051e-13, 1.075296e-13, 
    1.078089e-13, 1.07558e-13, 1.076025e-13, 1.078179e-13, 1.075716e-13, 
    1.081102e-13, 1.077451e-13, 1.08423e-13, 1.080587e-13, 1.084459e-13, 
    1.083756e-13, 1.084919e-13, 1.08596e-13, 1.087269e-13, 1.089682e-13, 
    1.089124e-13, 1.091141e-13, 1.070464e-13, 1.071708e-13, 1.071599e-13, 
    1.072901e-13, 1.073863e-13, 1.075948e-13, 1.079289e-13, 1.078033e-13, 
    1.080338e-13, 1.0808e-13, 1.077299e-13, 1.079449e-13, 1.072541e-13, 
    1.073657e-13, 1.072993e-13, 1.070562e-13, 1.078322e-13, 1.074342e-13, 
    1.081686e-13, 1.079534e-13, 1.085811e-13, 1.082691e-13, 1.088816e-13, 
    1.091429e-13, 1.093888e-13, 1.096756e-13, 1.072387e-13, 1.071542e-13, 
    1.073056e-13, 1.075147e-13, 1.077088e-13, 1.079666e-13, 1.07993e-13, 
    1.080412e-13, 1.081661e-13, 1.082711e-13, 1.080564e-13, 1.082974e-13, 
    1.073915e-13, 1.078667e-13, 1.071222e-13, 1.073465e-13, 1.075024e-13, 
    1.074341e-13, 1.07789e-13, 1.078725e-13, 1.082117e-13, 1.080365e-13, 
    1.090784e-13, 1.086179e-13, 1.098939e-13, 1.095379e-13, 1.071247e-13, 
    1.072385e-13, 1.076341e-13, 1.074459e-13, 1.079838e-13, 1.081159e-13, 
    1.082234e-13, 1.083606e-13, 1.083755e-13, 1.084568e-13, 1.083236e-13, 
    1.084515e-13, 1.079671e-13, 1.081837e-13, 1.07589e-13, 1.077338e-13, 
    1.076672e-13, 1.075941e-13, 1.078197e-13, 1.080597e-13, 1.08065e-13, 
    1.081418e-13, 1.083583e-13, 1.07986e-13, 1.091375e-13, 1.084267e-13, 
    1.073625e-13, 1.075813e-13, 1.076127e-13, 1.075279e-13, 1.081027e-13, 
    1.078946e-13, 1.084548e-13, 1.083035e-13, 1.085514e-13, 1.084282e-13, 
    1.084101e-13, 1.082519e-13, 1.081533e-13, 1.079041e-13, 1.077012e-13, 
    1.075402e-13, 1.075777e-13, 1.077545e-13, 1.080744e-13, 1.083768e-13, 
    1.083106e-13, 1.085326e-13, 1.079448e-13, 1.081913e-13, 1.080961e-13, 
    1.083445e-13, 1.078e-13, 1.082634e-13, 1.076813e-13, 1.077324e-13, 
    1.078905e-13, 1.08208e-13, 1.082784e-13, 1.083533e-13, 1.083071e-13, 
    1.080826e-13, 1.080458e-13, 1.078866e-13, 1.078426e-13, 1.077213e-13, 
    1.076208e-13, 1.077126e-13, 1.07809e-13, 1.080827e-13, 1.08329e-13, 
    1.085975e-13, 1.086631e-13, 1.089761e-13, 1.087212e-13, 1.091415e-13, 
    1.08784e-13, 1.094026e-13, 1.082904e-13, 1.087737e-13, 1.078977e-13, 
    1.079922e-13, 1.08163e-13, 1.085545e-13, 1.083433e-13, 1.085904e-13, 
    1.080444e-13, 1.077605e-13, 1.076872e-13, 1.0755e-13, 1.076903e-13, 
    1.076789e-13, 1.078131e-13, 1.077699e-13, 1.080918e-13, 1.07919e-13, 
    1.084096e-13, 1.085885e-13, 1.090929e-13, 1.094016e-13, 1.097157e-13, 
    1.098541e-13, 1.098963e-13, 1.099139e-13 ;

 LITR3C =
  9.697996e-06, 9.697987e-06, 9.697988e-06, 9.69798e-06, 9.697985e-06, 
    9.697979e-06, 9.697994e-06, 9.697986e-06, 9.697991e-06, 9.697995e-06, 
    9.697965e-06, 9.69798e-06, 9.697949e-06, 9.697959e-06, 9.697936e-06, 
    9.697951e-06, 9.697932e-06, 9.697936e-06, 9.697925e-06, 9.697927e-06, 
    9.697914e-06, 9.697923e-06, 9.697907e-06, 9.697917e-06, 9.697915e-06, 
    9.697924e-06, 9.697977e-06, 9.697967e-06, 9.697977e-06, 9.697976e-06, 
    9.697977e-06, 9.697985e-06, 9.697988e-06, 9.697997e-06, 9.697995e-06, 
    9.697989e-06, 9.697976e-06, 9.69798e-06, 9.697968e-06, 9.697968e-06, 
    9.697956e-06, 9.697961e-06, 9.697939e-06, 9.697946e-06, 9.697927e-06, 
    9.697932e-06, 9.697928e-06, 9.697929e-06, 9.697928e-06, 9.697935e-06, 
    9.697932e-06, 9.697937e-06, 9.69796e-06, 9.697954e-06, 9.697974e-06, 
    9.697986e-06, 9.697994e-06, 9.697999e-06, 9.697998e-06, 9.697997e-06, 
    9.697989e-06, 9.697982e-06, 9.697976e-06, 9.697972e-06, 9.697968e-06, 
    9.697957e-06, 9.697951e-06, 9.697938e-06, 9.69794e-06, 9.697937e-06, 
    9.697933e-06, 9.697927e-06, 9.697927e-06, 9.697925e-06, 9.697937e-06, 
    9.697928e-06, 9.697942e-06, 9.697938e-06, 9.697967e-06, 9.697978e-06, 
    9.697984e-06, 9.697987e-06, 9.697997e-06, 9.697991e-06, 9.697994e-06, 
    9.697987e-06, 9.697983e-06, 9.697985e-06, 9.697972e-06, 9.697977e-06, 
    9.697951e-06, 9.697962e-06, 9.697933e-06, 9.69794e-06, 9.697931e-06, 
    9.697936e-06, 9.697928e-06, 9.697935e-06, 9.697924e-06, 9.697921e-06, 
    9.697923e-06, 9.697916e-06, 9.697936e-06, 9.697928e-06, 9.697985e-06, 
    9.697985e-06, 9.697983e-06, 9.69799e-06, 9.69799e-06, 9.697997e-06, 
    9.697991e-06, 9.697988e-06, 9.697983e-06, 9.697979e-06, 9.697976e-06, 
    9.697968e-06, 9.69796e-06, 9.697948e-06, 9.697939e-06, 9.697934e-06, 
    9.697937e-06, 9.697935e-06, 9.697937e-06, 9.697939e-06, 9.697922e-06, 
    9.697932e-06, 9.697917e-06, 9.697917e-06, 9.697925e-06, 9.697917e-06, 
    9.697985e-06, 9.697987e-06, 9.697993e-06, 9.697987e-06, 9.697997e-06, 
    9.697992e-06, 9.697989e-06, 9.697977e-06, 9.697975e-06, 9.697972e-06, 
    9.697967e-06, 9.697961e-06, 9.69795e-06, 9.697941e-06, 9.697933e-06, 
    9.697933e-06, 9.697933e-06, 9.697931e-06, 9.697936e-06, 9.69793e-06, 
    9.697929e-06, 9.697932e-06, 9.697917e-06, 9.697922e-06, 9.697917e-06, 
    9.69792e-06, 9.697986e-06, 9.697982e-06, 9.697984e-06, 9.697981e-06, 
    9.697983e-06, 9.697973e-06, 9.69797e-06, 9.697956e-06, 9.697961e-06, 
    9.697952e-06, 9.69796e-06, 9.697958e-06, 9.697951e-06, 9.69796e-06, 
    9.697941e-06, 9.697954e-06, 9.697931e-06, 9.697943e-06, 9.69793e-06, 
    9.697933e-06, 9.697928e-06, 9.697925e-06, 9.69792e-06, 9.697913e-06, 
    9.697915e-06, 9.697907e-06, 9.697977e-06, 9.697973e-06, 9.697974e-06, 
    9.697969e-06, 9.697966e-06, 9.697959e-06, 9.697947e-06, 9.697952e-06, 
    9.697944e-06, 9.697943e-06, 9.697955e-06, 9.697947e-06, 9.69797e-06, 
    9.697967e-06, 9.697969e-06, 9.697977e-06, 9.697951e-06, 9.697965e-06, 
    9.697939e-06, 9.697947e-06, 9.697926e-06, 9.697937e-06, 9.697916e-06, 
    9.697907e-06, 9.697898e-06, 9.697888e-06, 9.697971e-06, 9.697974e-06, 
    9.697968e-06, 9.697962e-06, 9.697955e-06, 9.697947e-06, 9.697946e-06, 
    9.697944e-06, 9.697939e-06, 9.697936e-06, 9.697943e-06, 9.697936e-06, 
    9.697966e-06, 9.69795e-06, 9.697975e-06, 9.697967e-06, 9.697962e-06, 
    9.697965e-06, 9.697952e-06, 9.697949e-06, 9.697938e-06, 9.697944e-06, 
    9.697908e-06, 9.697925e-06, 9.697881e-06, 9.697893e-06, 9.697975e-06, 
    9.697971e-06, 9.697957e-06, 9.697964e-06, 9.697946e-06, 9.697941e-06, 
    9.697937e-06, 9.697933e-06, 9.697933e-06, 9.69793e-06, 9.697935e-06, 
    9.69793e-06, 9.697947e-06, 9.697939e-06, 9.697959e-06, 9.697955e-06, 
    9.697957e-06, 9.697959e-06, 9.697951e-06, 9.697943e-06, 9.697943e-06, 
    9.69794e-06, 9.697933e-06, 9.697946e-06, 9.697907e-06, 9.697931e-06, 
    9.697967e-06, 9.697959e-06, 9.697958e-06, 9.697961e-06, 9.697942e-06, 
    9.697949e-06, 9.69793e-06, 9.697935e-06, 9.697927e-06, 9.697931e-06, 
    9.697931e-06, 9.697937e-06, 9.69794e-06, 9.697948e-06, 9.697956e-06, 
    9.697961e-06, 9.697959e-06, 9.697954e-06, 9.697943e-06, 9.697933e-06, 
    9.697935e-06, 9.697927e-06, 9.697947e-06, 9.697938e-06, 9.697942e-06, 
    9.697934e-06, 9.697952e-06, 9.697937e-06, 9.697956e-06, 9.697955e-06, 
    9.697949e-06, 9.697938e-06, 9.697936e-06, 9.697933e-06, 9.697935e-06, 
    9.697943e-06, 9.697944e-06, 9.697949e-06, 9.69795e-06, 9.697955e-06, 
    9.697958e-06, 9.697955e-06, 9.697952e-06, 9.697943e-06, 9.697934e-06, 
    9.697925e-06, 9.697923e-06, 9.697912e-06, 9.697921e-06, 9.697907e-06, 
    9.697918e-06, 9.697897e-06, 9.697936e-06, 9.697919e-06, 9.697948e-06, 
    9.697946e-06, 9.69794e-06, 9.697927e-06, 9.697934e-06, 9.697926e-06, 
    9.697944e-06, 9.697954e-06, 9.697956e-06, 9.69796e-06, 9.697956e-06, 
    9.697957e-06, 9.697952e-06, 9.697953e-06, 9.697942e-06, 9.697948e-06, 
    9.697931e-06, 9.697926e-06, 9.697908e-06, 9.697897e-06, 9.697887e-06, 
    9.697883e-06, 9.697881e-06, 9.69788e-06 ;

 LITR3C_TO_SOIL2C =
  5.325308e-14, 5.339687e-14, 5.336894e-14, 5.34848e-14, 5.342056e-14, 
    5.34964e-14, 5.328226e-14, 5.340255e-14, 5.332579e-14, 5.326606e-14, 
    5.370932e-14, 5.348997e-14, 5.393699e-14, 5.379734e-14, 5.41479e-14, 
    5.391524e-14, 5.419478e-14, 5.414124e-14, 5.430243e-14, 5.425628e-14, 
    5.446213e-14, 5.432373e-14, 5.456879e-14, 5.442912e-14, 5.445096e-14, 
    5.431915e-14, 5.353419e-14, 5.368202e-14, 5.352542e-14, 5.354651e-14, 
    5.353706e-14, 5.342187e-14, 5.336376e-14, 5.324212e-14, 5.326421e-14, 
    5.335357e-14, 5.3556e-14, 5.348735e-14, 5.366039e-14, 5.365648e-14, 
    5.384884e-14, 5.376214e-14, 5.408506e-14, 5.399339e-14, 5.425821e-14, 
    5.419164e-14, 5.425507e-14, 5.423584e-14, 5.425532e-14, 5.415769e-14, 
    5.419952e-14, 5.411359e-14, 5.377838e-14, 5.387697e-14, 5.358267e-14, 
    5.340533e-14, 5.328753e-14, 5.320385e-14, 5.321568e-14, 5.323823e-14, 
    5.335409e-14, 5.346298e-14, 5.35459e-14, 5.360133e-14, 5.365592e-14, 
    5.382092e-14, 5.390828e-14, 5.410357e-14, 5.406838e-14, 5.412801e-14, 
    5.418502e-14, 5.428062e-14, 5.426489e-14, 5.430698e-14, 5.412647e-14, 
    5.424645e-14, 5.404835e-14, 5.410254e-14, 5.36706e-14, 5.350588e-14, 
    5.343567e-14, 5.33743e-14, 5.322478e-14, 5.332804e-14, 5.328734e-14, 
    5.338419e-14, 5.344567e-14, 5.341527e-14, 5.360284e-14, 5.352994e-14, 
    5.391346e-14, 5.37484e-14, 5.417837e-14, 5.407561e-14, 5.4203e-14, 
    5.413802e-14, 5.424933e-14, 5.414915e-14, 5.432266e-14, 5.436039e-14, 
    5.43346e-14, 5.443368e-14, 5.414359e-14, 5.425506e-14, 5.341442e-14, 
    5.341937e-14, 5.344248e-14, 5.334086e-14, 5.333465e-14, 5.32415e-14, 
    5.33244e-14, 5.335968e-14, 5.344925e-14, 5.350217e-14, 5.355248e-14, 
    5.366301e-14, 5.378633e-14, 5.395862e-14, 5.408227e-14, 5.41651e-14, 
    5.411432e-14, 5.415915e-14, 5.410903e-14, 5.408554e-14, 5.434624e-14, 
    5.41999e-14, 5.441944e-14, 5.44073e-14, 5.430797e-14, 5.440867e-14, 
    5.342286e-14, 5.339432e-14, 5.329516e-14, 5.337277e-14, 5.323136e-14, 
    5.331051e-14, 5.335599e-14, 5.353143e-14, 5.356999e-14, 5.360568e-14, 
    5.367618e-14, 5.376658e-14, 5.392502e-14, 5.406271e-14, 5.418834e-14, 
    5.417914e-14, 5.418238e-14, 5.421041e-14, 5.414094e-14, 5.422182e-14, 
    5.423537e-14, 5.419991e-14, 5.440568e-14, 5.434692e-14, 5.440705e-14, 
    5.43688e-14, 5.34036e-14, 5.345161e-14, 5.342567e-14, 5.347445e-14, 
    5.344007e-14, 5.359281e-14, 5.363856e-14, 5.385252e-14, 5.376479e-14, 
    5.390443e-14, 5.3779e-14, 5.380122e-14, 5.390892e-14, 5.378579e-14, 
    5.405509e-14, 5.387252e-14, 5.42115e-14, 5.402933e-14, 5.422291e-14, 
    5.41878e-14, 5.424594e-14, 5.429798e-14, 5.436344e-14, 5.448409e-14, 
    5.445617e-14, 5.455704e-14, 5.352318e-14, 5.358538e-14, 5.357994e-14, 
    5.364503e-14, 5.369314e-14, 5.37974e-14, 5.396441e-14, 5.390164e-14, 
    5.401689e-14, 5.404e-14, 5.386492e-14, 5.397242e-14, 5.362702e-14, 
    5.368285e-14, 5.364964e-14, 5.352807e-14, 5.391607e-14, 5.371706e-14, 
    5.40843e-14, 5.397671e-14, 5.429055e-14, 5.413452e-14, 5.444079e-14, 
    5.457142e-14, 5.469439e-14, 5.483777e-14, 5.361935e-14, 5.357709e-14, 
    5.365277e-14, 5.375736e-14, 5.38544e-14, 5.398327e-14, 5.399646e-14, 
    5.402058e-14, 5.408304e-14, 5.413554e-14, 5.402817e-14, 5.41487e-14, 
    5.369574e-14, 5.393334e-14, 5.356109e-14, 5.367325e-14, 5.375121e-14, 
    5.371704e-14, 5.389447e-14, 5.393625e-14, 5.410582e-14, 5.401822e-14, 
    5.453916e-14, 5.430892e-14, 5.494694e-14, 5.476894e-14, 5.356232e-14, 
    5.361922e-14, 5.381702e-14, 5.372295e-14, 5.399188e-14, 5.405795e-14, 
    5.411169e-14, 5.418031e-14, 5.418774e-14, 5.422837e-14, 5.416177e-14, 
    5.422576e-14, 5.398354e-14, 5.409183e-14, 5.379446e-14, 5.386689e-14, 
    5.383359e-14, 5.379702e-14, 5.390983e-14, 5.402986e-14, 5.403247e-14, 
    5.40709e-14, 5.417911e-14, 5.399297e-14, 5.456876e-14, 5.421336e-14, 
    5.368124e-14, 5.379065e-14, 5.380633e-14, 5.376395e-14, 5.405136e-14, 
    5.394728e-14, 5.422739e-14, 5.415175e-14, 5.427568e-14, 5.42141e-14, 
    5.420504e-14, 5.412592e-14, 5.407663e-14, 5.395205e-14, 5.385059e-14, 
    5.37701e-14, 5.378882e-14, 5.387722e-14, 5.403721e-14, 5.418839e-14, 
    5.415527e-14, 5.426626e-14, 5.39724e-14, 5.409566e-14, 5.404803e-14, 
    5.417223e-14, 5.389996e-14, 5.41317e-14, 5.384064e-14, 5.38662e-14, 
    5.394522e-14, 5.410398e-14, 5.413916e-14, 5.417663e-14, 5.415352e-14, 
    5.404127e-14, 5.402289e-14, 5.394331e-14, 5.39213e-14, 5.386064e-14, 
    5.381036e-14, 5.385628e-14, 5.390448e-14, 5.404135e-14, 5.416451e-14, 
    5.429871e-14, 5.433155e-14, 5.448801e-14, 5.436059e-14, 5.457072e-14, 
    5.439199e-14, 5.470129e-14, 5.414519e-14, 5.438683e-14, 5.394883e-14, 
    5.39961e-14, 5.408147e-14, 5.427726e-14, 5.417165e-14, 5.429517e-14, 
    5.402218e-14, 5.388025e-14, 5.384356e-14, 5.377499e-14, 5.384513e-14, 
    5.383943e-14, 5.390651e-14, 5.388496e-14, 5.404589e-14, 5.395947e-14, 
    5.42048e-14, 5.429421e-14, 5.454645e-14, 5.470081e-14, 5.485782e-14, 
    5.492705e-14, 5.494812e-14, 5.495692e-14 ;

 LITR3C_vr =
  0.0005537656, 0.000553765, 0.0005537652, 0.0005537647, 0.0005537649, 
    0.0005537646, 0.0005537655, 0.000553765, 0.0005537653, 0.0005537656, 
    0.0005537638, 0.0005537647, 0.0005537629, 0.0005537635, 0.0005537621, 
    0.000553763, 0.000553762, 0.0005537621, 0.0005537616, 0.0005537617, 
    0.0005537609, 0.0005537614, 0.0005537605, 0.000553761, 0.000553761, 
    0.0005537614, 0.0005537645, 0.0005537639, 0.0005537645, 0.0005537645, 
    0.0005537645, 0.0005537649, 0.0005537652, 0.0005537656, 0.0005537656, 
    0.0005537652, 0.0005537644, 0.0005537647, 0.000553764, 0.0005537641, 
    0.0005537633, 0.0005537636, 0.0005537624, 0.0005537627, 0.0005537617, 
    0.000553762, 0.0005537617, 0.0005537618, 0.0005537617, 0.0005537621, 
    0.0005537619, 0.0005537622, 0.0005537635, 0.0005537632, 0.0005537643, 
    0.000553765, 0.0005537655, 0.0005537658, 0.0005537657, 0.0005537656, 
    0.0005537652, 0.0005537648, 0.0005537645, 0.0005537642, 0.0005537641, 
    0.0005537634, 0.0005537631, 0.0005537623, 0.0005537624, 0.0005537622, 
    0.000553762, 0.0005537616, 0.0005537617, 0.0005537615, 0.0005537622, 
    0.0005537617, 0.0005537625, 0.0005537623, 0.000553764, 0.0005537646, 
    0.0005537649, 0.0005537651, 0.0005537657, 0.0005537653, 0.0005537655, 
    0.0005537651, 0.0005537649, 0.000553765, 0.0005537642, 0.0005537645, 
    0.000553763, 0.0005537636, 0.000553762, 0.0005537624, 0.0005537619, 
    0.0005537621, 0.0005537617, 0.0005537621, 0.0005537614, 0.0005537613, 
    0.0005537614, 0.000553761, 0.0005537621, 0.0005537617, 0.000553765, 
    0.0005537649, 0.0005537649, 0.0005537653, 0.0005537653, 0.0005537656, 
    0.0005537653, 0.0005537652, 0.0005537648, 0.0005537646, 0.0005537644, 
    0.000553764, 0.0005537635, 0.0005537628, 0.0005537624, 0.0005537621, 
    0.0005537622, 0.0005537621, 0.0005537622, 0.0005537624, 0.0005537614, 
    0.0005537619, 0.0005537611, 0.0005537611, 0.0005537615, 0.0005537611, 
    0.0005537649, 0.000553765, 0.0005537655, 0.0005537651, 0.0005537657, 
    0.0005537654, 0.0005537652, 0.0005537645, 0.0005537643, 0.0005537642, 
    0.0005537639, 0.0005537636, 0.000553763, 0.0005537625, 0.000553762, 
    0.000553762, 0.000553762, 0.0005537619, 0.0005537621, 0.0005537618, 
    0.0005537618, 0.0005537619, 0.0005537611, 0.0005537614, 0.0005537611, 
    0.0005537613, 0.000553765, 0.0005537648, 0.0005537649, 0.0005537648, 
    0.0005537649, 0.0005537643, 0.0005537641, 0.0005537632, 0.0005537636, 
    0.0005537631, 0.0005537635, 0.0005537635, 0.0005537631, 0.0005537635, 
    0.0005537625, 0.0005537632, 0.0005537619, 0.0005537626, 0.0005537618, 
    0.000553762, 0.0005537617, 0.0005537616, 0.0005537613, 0.0005537608, 
    0.0005537609, 0.0005537606, 0.0005537645, 0.0005537643, 0.0005537643, 
    0.0005537641, 0.0005537639, 0.0005537635, 0.0005537628, 0.0005537631, 
    0.0005537627, 0.0005537625, 0.0005537632, 0.0005537628, 0.0005537641, 
    0.0005537639, 0.0005537641, 0.0005537645, 0.000553763, 0.0005537638, 
    0.0005537624, 0.0005537628, 0.0005537616, 0.0005537622, 0.000553761, 
    0.0005537605, 0.00055376, 0.0005537595, 0.0005537642, 0.0005537643, 
    0.0005537641, 0.0005537636, 0.0005537632, 0.0005537628, 0.0005537627, 
    0.0005537626, 0.0005537624, 0.0005537622, 0.0005537626, 0.0005537621, 
    0.0005537639, 0.0005537629, 0.0005537644, 0.0005537639, 0.0005537636, 
    0.0005537638, 0.0005537631, 0.0005537629, 0.0005537623, 0.0005537626, 
    0.0005537606, 0.0005537615, 0.000553759, 0.0005537597, 0.0005537644, 
    0.0005537642, 0.0005537634, 0.0005537638, 0.0005537627, 0.0005537625, 
    0.0005537622, 0.000553762, 0.000553762, 0.0005537618, 0.0005537621, 
    0.0005537618, 0.0005537628, 0.0005537624, 0.0005537635, 0.0005537632, 
    0.0005537634, 0.0005537635, 0.0005537631, 0.0005537626, 0.0005537626, 
    0.0005537624, 0.000553762, 0.0005537627, 0.0005537605, 0.0005537618, 
    0.0005537639, 0.0005537635, 0.0005537635, 0.0005537636, 0.0005537625, 
    0.0005537629, 0.0005537618, 0.0005537621, 0.0005537616, 0.0005537618, 
    0.0005537619, 0.0005537622, 0.0005537624, 0.0005537629, 0.0005537633, 
    0.0005537636, 0.0005537635, 0.0005537632, 0.0005537625, 0.000553762, 
    0.0005537621, 0.0005537617, 0.0005537628, 0.0005537623, 0.0005537625, 
    0.000553762, 0.0005537631, 0.0005537622, 0.0005537633, 0.0005537632, 
    0.0005537629, 0.0005537623, 0.0005537621, 0.000553762, 0.0005537621, 
    0.0005537625, 0.0005537626, 0.0005537629, 0.000553763, 0.0005537632, 
    0.0005537634, 0.0005537632, 0.0005537631, 0.0005537625, 0.0005537621, 
    0.0005537616, 0.0005537614, 0.0005537608, 0.0005537613, 0.0005537605, 
    0.0005537612, 0.00055376, 0.0005537621, 0.0005537612, 0.0005537629, 
    0.0005537627, 0.0005537624, 0.0005537616, 0.000553762, 0.0005537616, 
    0.0005537626, 0.0005537632, 0.0005537633, 0.0005537636, 0.0005537633, 
    0.0005537633, 0.0005537631, 0.0005537631, 0.0005537625, 0.0005537628, 
    0.0005537619, 0.0005537616, 0.0005537606, 0.00055376, 0.0005537594, 
    0.0005537591, 0.000553759, 0.000553759,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342132e-07, 1.34213e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 
    1.342129e-07, 1.342131e-07, 1.34213e-07, 1.342131e-07, 1.342132e-07, 
    1.342127e-07, 1.342129e-07, 1.342125e-07, 1.342127e-07, 1.342123e-07, 
    1.342125e-07, 1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342122e-07, 
    1.34212e-07, 1.342122e-07, 1.342119e-07, 1.342121e-07, 1.34212e-07, 
    1.342122e-07, 1.342129e-07, 1.342128e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 1.342128e-07, 
    1.342126e-07, 1.342127e-07, 1.342124e-07, 1.342125e-07, 1.342122e-07, 
    1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342122e-07, 1.342123e-07, 
    1.342123e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 1.342129e-07, 
    1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 
    1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342122e-07, 1.342123e-07, 
    1.342122e-07, 1.342124e-07, 1.342124e-07, 1.342128e-07, 1.342129e-07, 
    1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.34213e-07, 1.34213e-07, 1.34213e-07, 1.342128e-07, 1.342129e-07, 
    1.342125e-07, 1.342127e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342123e-07, 1.342122e-07, 1.342121e-07, 
    1.342122e-07, 1.342121e-07, 1.342123e-07, 1.342122e-07, 1.34213e-07, 
    1.34213e-07, 1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342124e-07, 1.342123e-07, 
    1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342124e-07, 1.342121e-07, 
    1.342123e-07, 1.342121e-07, 1.342121e-07, 1.342122e-07, 1.342121e-07, 
    1.34213e-07, 1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 
    1.342122e-07, 1.342123e-07, 1.342121e-07, 1.342121e-07, 1.342121e-07, 
    1.342121e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342126e-07, 1.342127e-07, 
    1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 
    1.342124e-07, 1.342126e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342121e-07, 1.34212e-07, 
    1.34212e-07, 1.342119e-07, 1.342129e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342126e-07, 1.342125e-07, 1.342128e-07, 
    1.342128e-07, 1.342128e-07, 1.342129e-07, 1.342125e-07, 1.342127e-07, 
    1.342124e-07, 1.342125e-07, 1.342122e-07, 1.342123e-07, 1.342121e-07, 
    1.342119e-07, 1.342118e-07, 1.342117e-07, 1.342128e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342125e-07, 
    1.342124e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342128e-07, 1.342125e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342124e-07, 1.342124e-07, 
    1.34212e-07, 1.342122e-07, 1.342116e-07, 1.342117e-07, 1.342129e-07, 
    1.342128e-07, 1.342126e-07, 1.342127e-07, 1.342125e-07, 1.342124e-07, 
    1.342124e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 
    1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 
    1.342124e-07, 1.342123e-07, 1.342125e-07, 1.342119e-07, 1.342123e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 1.342124e-07, 
    1.342125e-07, 1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342124e-07, 1.342125e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342125e-07, 1.342124e-07, 1.342124e-07, 
    1.342123e-07, 1.342126e-07, 1.342123e-07, 1.342126e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 
    1.342124e-07, 1.342124e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342123e-07, 
    1.342122e-07, 1.342122e-07, 1.34212e-07, 1.342121e-07, 1.342119e-07, 
    1.342121e-07, 1.342118e-07, 1.342123e-07, 1.342121e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342122e-07, 1.342123e-07, 1.342122e-07, 
    1.342124e-07, 1.342126e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 
    1.342123e-07, 1.342122e-07, 1.34212e-07, 1.342118e-07, 1.342117e-07, 
    1.342116e-07, 1.342116e-07, 1.342116e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  -2.573451e-26, -4.901811e-26, -3.186177e-26, -3.798904e-26, 4.901811e-27, 
    -1.593089e-26, 1.200944e-25, 5.391992e-26, -5.514538e-26, 6.372354e-26, 
    -9.313441e-26, 6.127264e-27, -8.210533e-26, -9.313441e-26, 3.063632e-26, 
    1.715634e-26, 9.803622e-26, 2.941087e-26, -9.068351e-26, -6.249809e-26, 
    -3.186177e-26, -4.901811e-27, -1.225453e-27, 2.695996e-26, -6.127264e-27, 
    -3.921449e-26, 1.593089e-26, -1.838179e-26, -3.798904e-26, -2.573451e-26, 
    -3.676358e-26, 1.213198e-25, 4.41163e-26, 2.695996e-26, 6.372354e-26, 
    6.73999e-26, -1.960724e-26, 5.269447e-26, 2.695996e-26, 4.65672e-26, 
    2.08327e-26, -7.230172e-26, -5.637083e-26, 4.901811e-27, 8.578169e-27, 
    -1.017126e-25, -6.127264e-26, -1.078398e-25, 0, 1.225453e-27, 
    3.553813e-26, -3.798904e-26, -1.56858e-25, -4.901811e-27, -4.41163e-26, 
    4.289085e-26, 2.450905e-26, 6.004719e-26, -6.862535e-26, -1.151926e-25, 
    1.838179e-26, -2.32836e-26, 1.102908e-26, -6.127264e-27, 3.308722e-26, 
    1.985233e-25, -5.882173e-26, -5.637083e-26, -1.127417e-25, 4.043994e-26, 
    -2.32836e-26, 5.514538e-26, 8.087988e-26, 7.597807e-26, 1.225453e-26, 
    -5.514538e-26, 1.825925e-25, -1.115162e-25, -3.676358e-26, -5.146902e-26, 
    3.553813e-26, -8.087988e-26, -4.65672e-26, 4.41163e-26, -6.127264e-27, 
    -4.901811e-27, -1.960724e-26, -1.715634e-26, -1.115162e-25, 
    -4.901811e-27, 9.068351e-26, -8.087988e-26, -3.308722e-26, 1.102908e-26, 
    2.205815e-26, -4.534175e-26, 4.043994e-26, -1.017126e-25, 1.703379e-25, 
    4.901811e-26, -1.176435e-25, -9.313441e-26, -1.102908e-26, -3.063632e-26, 
    -4.043994e-26, -1.911706e-25, 4.901811e-27, 1.470543e-26, 6.617445e-26, 
    5.759628e-26, -6.127264e-27, -9.558531e-26, -2.450906e-27, -1.311234e-25, 
    -1.151926e-25, 1.715634e-26, 1.593089e-26, 3.798904e-26, 1.347998e-26, 
    -6.004719e-26, 2.205815e-26, 9.558531e-26, 1.225453e-26, 7.965443e-26, 
    4.901811e-27, -7.230172e-26, 7.352717e-27, 7.107626e-26, 8.455624e-26, 
    6.617445e-26, 2.08327e-26, -1.372507e-25, 3.553813e-26, 6.004719e-26, 
    -6.249809e-26, 3.921449e-26, -4.289085e-26, 8.700715e-26, 1.225453e-26, 
    -5.024356e-26, -9.803622e-27, -6.372354e-26, 4.65672e-26, 4.901811e-27, 
    -9.803622e-26, 2.450906e-27, 6.249809e-26, 4.41163e-26, 5.637083e-26, 
    -9.313441e-26, -2.205815e-26, -1.188689e-25, 1.715634e-26, 0, 
    9.313441e-26, 6.127264e-26, 6.862535e-26, -5.391992e-26, -7.352717e-27, 
    2.941087e-26, -2.573451e-26, -1.347998e-26, 4.65672e-26, -7.475262e-26, 
    2.32836e-26, -8.578169e-26, 8.455624e-26, -1.017126e-25, 4.043994e-26, 
    1.041635e-25, -6.127264e-26, -8.700715e-26, 1.02938e-25, 6.127264e-26, 
    1.004871e-25, 2.695996e-26, 5.391992e-26, -6.617445e-26, -1.004871e-25, 
    -2.205815e-26, 3.431268e-26, 7.107626e-26, 1.225453e-27, -6.127264e-27, 
    2.695996e-26, -2.573451e-26, 7.475262e-26, -4.41163e-26, 4.41163e-26, 
    -5.514538e-26, -1.102908e-25, 1.838179e-26, -5.269447e-26, 7.352717e-27, 
    -1.495052e-25, 5.514538e-26, 7.842898e-26, 1.347998e-25, 2.573451e-26, 
    1.556325e-25, 3.798904e-26, 2.08327e-26, 5.146902e-26, 1.470543e-26, 
    1.004871e-25, -1.102908e-25, -5.759628e-26, 9.068351e-26, -9.681077e-26, 
    -8.210533e-26, -4.534175e-26, 8.700715e-26, 9.190896e-26, -8.945805e-26, 
    1.593089e-26, -6.98508e-26, 3.676358e-27, -5.269447e-26, -2.818541e-26, 
    7.352717e-26, 1.347998e-26, -7.107626e-26, 9.803622e-27, 1.102908e-26, 
    4.043994e-26, -4.41163e-26, 1.02938e-25, 1.225453e-26, -1.225453e-26, 
    -2.450905e-26, -1.102908e-26, -5.024356e-26, 1.102908e-26, -2.941087e-26, 
    8.578169e-27, 5.024356e-26, -8.455624e-26, 8.333079e-26, -1.225453e-26, 
    5.882173e-26, 5.391992e-26, 1.776906e-25, 8.700715e-26, 1.286725e-25, 
    -6.127264e-26, 1.372507e-25, -2.695996e-26, 1.43378e-25, -1.666616e-25, 
    3.553813e-26, 4.901811e-26, 1.960724e-26, -1.715634e-26, 4.534175e-26, 
    3.186177e-26, -3.063632e-26, 2.450906e-27, -4.534175e-26, 2.695996e-26, 
    5.514538e-26, 9.313441e-26, 9.803622e-26, 6.862535e-26, -3.798904e-26, 
    3.676358e-26, -7.230172e-26, 7.720352e-26, -1.29898e-25, -4.166539e-26, 
    -4.534175e-26, 7.965443e-26, -1.642107e-25, -3.431268e-26, -3.063632e-26, 
    -1.188689e-25, -3.431268e-26, -1.225453e-26, -1.507307e-25, 
    -1.347998e-26, -9.681077e-26, 5.024356e-26, 1.838179e-26, 1.715634e-26, 
    -1.838179e-26, -5.146902e-26, -2.818541e-26, 9.803622e-27, 2.573451e-26, 
    7.652491e-42, -4.043994e-26, 5.146902e-26, -6.127264e-27, -3.676358e-27, 
    -5.882173e-26, -1.715634e-26, 2.941087e-26, -1.347998e-26, 7.107626e-26, 
    -2.573451e-26, -8.578169e-26, -1.225453e-26, -6.617445e-26, 
    -1.262216e-25, -1.752397e-25, -7.230172e-26, -1.593089e-26, 
    -1.960724e-26, -2.695996e-26, 4.043994e-26, -4.534175e-26, 1.397016e-25, 
    6.249809e-26, -4.779266e-26, -4.534175e-26, -4.534175e-26, -5.391992e-26, 
    2.450906e-27, -1.838179e-26, 2.818541e-26, 5.391992e-26, -2.695996e-26, 
    6.4949e-26, 9.803622e-27, 1.446034e-25, 0, 6.73999e-26, -4.901811e-26, 
    7.597807e-26, -9.190896e-26, 1.053889e-25, 6.004719e-26, 4.166539e-26, 
    6.4949e-26, -3.431268e-26, 2.450906e-27, -1.102908e-26, -1.151926e-25, 
    7.352717e-26,
  1.338125e-32, 1.338123e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338124e-32, 1.338123e-32, 1.338124e-32, 1.338125e-32, 
    1.33812e-32, 1.338123e-32, 1.338118e-32, 1.33812e-32, 1.338116e-32, 
    1.338119e-32, 1.338116e-32, 1.338116e-32, 1.338115e-32, 1.338115e-32, 
    1.338113e-32, 1.338115e-32, 1.338112e-32, 1.338114e-32, 1.338113e-32, 
    1.338115e-32, 1.338122e-32, 1.338121e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338122e-32, 1.338123e-32, 1.338121e-32, 1.338121e-32, 
    1.338119e-32, 1.33812e-32, 1.338117e-32, 1.338118e-32, 1.338115e-32, 
    1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338115e-32, 1.338116e-32, 
    1.338116e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 1.338122e-32, 
    1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 
    1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 
    1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338115e-32, 1.338117e-32, 
    1.338115e-32, 1.338117e-32, 1.338117e-32, 1.338121e-32, 1.338122e-32, 
    1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338121e-32, 1.338122e-32, 
    1.338119e-32, 1.33812e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338116e-32, 1.338115e-32, 1.338114e-32, 
    1.338115e-32, 1.338114e-32, 1.338116e-32, 1.338115e-32, 1.338123e-32, 
    1.338123e-32, 1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338117e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338117e-32, 1.338114e-32, 
    1.338116e-32, 1.338114e-32, 1.338114e-32, 1.338115e-32, 1.338114e-32, 
    1.338123e-32, 1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 
    1.338115e-32, 1.338116e-32, 1.338114e-32, 1.338114e-32, 1.338114e-32, 
    1.338114e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338121e-32, 1.338121e-32, 1.338119e-32, 1.33812e-32, 
    1.338119e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 1.33812e-32, 
    1.338117e-32, 1.338119e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338114e-32, 1.338113e-32, 
    1.338113e-32, 1.338113e-32, 1.338122e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338119e-32, 
    1.338118e-32, 1.338117e-32, 1.338119e-32, 1.338118e-32, 1.338121e-32, 
    1.338121e-32, 1.338121e-32, 1.338122e-32, 1.338119e-32, 1.33812e-32, 
    1.338117e-32, 1.338118e-32, 1.338115e-32, 1.338117e-32, 1.338114e-32, 
    1.338112e-32, 1.338111e-32, 1.33811e-32, 1.338121e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338116e-32, 
    1.338121e-32, 1.338118e-32, 1.338122e-32, 1.338121e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 1.338118e-32, 
    1.338113e-32, 1.338115e-32, 1.338109e-32, 1.33811e-32, 1.338122e-32, 
    1.338121e-32, 1.338119e-32, 1.33812e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 
    1.338116e-32, 1.338118e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338118e-32, 1.338112e-32, 1.338116e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338117e-32, 
    1.338118e-32, 1.338116e-32, 1.338116e-32, 1.338115e-32, 1.338116e-32, 
    1.338116e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338119e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338118e-32, 1.338117e-32, 1.338117e-32, 
    1.338116e-32, 1.338119e-32, 1.338117e-32, 1.338119e-32, 1.338119e-32, 
    1.338118e-32, 1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 
    1.338117e-32, 1.338118e-32, 1.338118e-32, 1.338118e-32, 1.338119e-32, 
    1.33812e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338116e-32, 
    1.338115e-32, 1.338115e-32, 1.338113e-32, 1.338114e-32, 1.338112e-32, 
    1.338114e-32, 1.338111e-32, 1.338116e-32, 1.338114e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338115e-32, 1.338116e-32, 1.338115e-32, 
    1.338118e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338116e-32, 1.338115e-32, 1.338113e-32, 1.338111e-32, 1.33811e-32, 
    1.338109e-32, 1.338109e-32, 1.338109e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.473967e-15, 1.477947e-15, 1.477174e-15, 1.480381e-15, 1.478603e-15, 
    1.480702e-15, 1.474775e-15, 1.478105e-15, 1.47598e-15, 1.474327e-15, 
    1.486596e-15, 1.480524e-15, 1.492897e-15, 1.489032e-15, 1.498735e-15, 
    1.492295e-15, 1.500032e-15, 1.49855e-15, 1.503012e-15, 1.501734e-15, 
    1.507432e-15, 1.503601e-15, 1.510384e-15, 1.506518e-15, 1.507123e-15, 
    1.503475e-15, 1.481748e-15, 1.48584e-15, 1.481505e-15, 1.482089e-15, 
    1.481827e-15, 1.478639e-15, 1.477031e-15, 1.473664e-15, 1.474276e-15, 
    1.476749e-15, 1.482352e-15, 1.480451e-15, 1.485241e-15, 1.485133e-15, 
    1.490457e-15, 1.488058e-15, 1.496995e-15, 1.494458e-15, 1.501788e-15, 
    1.499945e-15, 1.501701e-15, 1.501169e-15, 1.501708e-15, 1.499006e-15, 
    1.500164e-15, 1.497785e-15, 1.488507e-15, 1.491236e-15, 1.48309e-15, 
    1.478181e-15, 1.474921e-15, 1.472605e-15, 1.472932e-15, 1.473556e-15, 
    1.476763e-15, 1.479777e-15, 1.482072e-15, 1.483606e-15, 1.485117e-15, 
    1.489684e-15, 1.492102e-15, 1.497508e-15, 1.496534e-15, 1.498184e-15, 
    1.499762e-15, 1.502408e-15, 1.501973e-15, 1.503138e-15, 1.498142e-15, 
    1.501462e-15, 1.495979e-15, 1.497479e-15, 1.485524e-15, 1.480964e-15, 
    1.479021e-15, 1.477323e-15, 1.473184e-15, 1.476042e-15, 1.474916e-15, 
    1.477596e-15, 1.479298e-15, 1.478457e-15, 1.483648e-15, 1.481631e-15, 
    1.492246e-15, 1.487677e-15, 1.499578e-15, 1.496734e-15, 1.50026e-15, 
    1.498461e-15, 1.501542e-15, 1.498769e-15, 1.503572e-15, 1.504616e-15, 
    1.503902e-15, 1.506645e-15, 1.498615e-15, 1.501701e-15, 1.478433e-15, 
    1.47857e-15, 1.47921e-15, 1.476397e-15, 1.476225e-15, 1.473647e-15, 
    1.475941e-15, 1.476918e-15, 1.479397e-15, 1.480862e-15, 1.482254e-15, 
    1.485314e-15, 1.488727e-15, 1.493496e-15, 1.496918e-15, 1.499211e-15, 
    1.497805e-15, 1.499046e-15, 1.497659e-15, 1.497009e-15, 1.504224e-15, 
    1.500174e-15, 1.50625e-15, 1.505915e-15, 1.503165e-15, 1.505952e-15, 
    1.478666e-15, 1.477877e-15, 1.475132e-15, 1.47728e-15, 1.473366e-15, 
    1.475557e-15, 1.476816e-15, 1.481672e-15, 1.482739e-15, 1.483727e-15, 
    1.485678e-15, 1.48818e-15, 1.492566e-15, 1.496377e-15, 1.499854e-15, 
    1.4996e-15, 1.499689e-15, 1.500465e-15, 1.498542e-15, 1.500781e-15, 
    1.501156e-15, 1.500174e-15, 1.50587e-15, 1.504243e-15, 1.505907e-15, 
    1.504849e-15, 1.478134e-15, 1.479463e-15, 1.478744e-15, 1.480094e-15, 
    1.479143e-15, 1.48337e-15, 1.484637e-15, 1.490559e-15, 1.488131e-15, 
    1.491996e-15, 1.488524e-15, 1.489139e-15, 1.49212e-15, 1.488712e-15, 
    1.496166e-15, 1.491113e-15, 1.500495e-15, 1.495453e-15, 1.500811e-15, 
    1.499839e-15, 1.501448e-15, 1.502889e-15, 1.5047e-15, 1.50804e-15, 
    1.507267e-15, 1.510059e-15, 1.481443e-15, 1.483165e-15, 1.483014e-15, 
    1.484816e-15, 1.486148e-15, 1.489033e-15, 1.493656e-15, 1.491919e-15, 
    1.495108e-15, 1.495748e-15, 1.490902e-15, 1.493877e-15, 1.484317e-15, 
    1.485863e-15, 1.484943e-15, 1.481579e-15, 1.492318e-15, 1.48681e-15, 
    1.496974e-15, 1.493996e-15, 1.502683e-15, 1.498364e-15, 1.506841e-15, 
    1.510457e-15, 1.513861e-15, 1.517829e-15, 1.484105e-15, 1.482936e-15, 
    1.48503e-15, 1.487925e-15, 1.490611e-15, 1.494178e-15, 1.494543e-15, 
    1.495211e-15, 1.496939e-15, 1.498392e-15, 1.495421e-15, 1.498757e-15, 
    1.486219e-15, 1.492796e-15, 1.482493e-15, 1.485597e-15, 1.487755e-15, 
    1.486809e-15, 1.49172e-15, 1.492876e-15, 1.49757e-15, 1.495145e-15, 
    1.509564e-15, 1.503191e-15, 1.520851e-15, 1.515924e-15, 1.482527e-15, 
    1.484102e-15, 1.489576e-15, 1.486973e-15, 1.494416e-15, 1.496245e-15, 
    1.497733e-15, 1.499632e-15, 1.499837e-15, 1.500962e-15, 1.499119e-15, 
    1.50089e-15, 1.494185e-15, 1.497183e-15, 1.488952e-15, 1.490957e-15, 
    1.490035e-15, 1.489023e-15, 1.492145e-15, 1.495467e-15, 1.49554e-15, 
    1.496603e-15, 1.499599e-15, 1.494446e-15, 1.510383e-15, 1.500546e-15, 
    1.485818e-15, 1.488847e-15, 1.489281e-15, 1.488108e-15, 1.496063e-15, 
    1.493182e-15, 1.500935e-15, 1.498841e-15, 1.502271e-15, 1.500567e-15, 
    1.500316e-15, 1.498126e-15, 1.496762e-15, 1.493314e-15, 1.490505e-15, 
    1.488278e-15, 1.488796e-15, 1.491243e-15, 1.495671e-15, 1.499855e-15, 
    1.498939e-15, 1.502011e-15, 1.493877e-15, 1.497289e-15, 1.495971e-15, 
    1.499408e-15, 1.491872e-15, 1.498286e-15, 1.49023e-15, 1.490937e-15, 
    1.493125e-15, 1.497519e-15, 1.498493e-15, 1.49953e-15, 1.49889e-15, 
    1.495783e-15, 1.495275e-15, 1.493072e-15, 1.492463e-15, 1.490784e-15, 
    1.489392e-15, 1.490663e-15, 1.491997e-15, 1.495785e-15, 1.499194e-15, 
    1.502909e-15, 1.503818e-15, 1.508149e-15, 1.504622e-15, 1.510438e-15, 
    1.505491e-15, 1.514052e-15, 1.49866e-15, 1.505348e-15, 1.493225e-15, 
    1.494533e-15, 1.496896e-15, 1.502315e-15, 1.499392e-15, 1.502811e-15, 
    1.495255e-15, 1.491326e-15, 1.490311e-15, 1.488413e-15, 1.490354e-15, 
    1.490197e-15, 1.492053e-15, 1.491457e-15, 1.495911e-15, 1.493519e-15, 
    1.50031e-15, 1.502784e-15, 1.509766e-15, 1.514038e-15, 1.518384e-15, 
    1.5203e-15, 1.520884e-15, 1.521127e-15 ;

 LITR3N_vr =
  7.663711e-06, 7.663702e-06, 7.663704e-06, 7.663698e-06, 7.663702e-06, 
    7.663697e-06, 7.663709e-06, 7.663702e-06, 7.663707e-06, 7.66371e-06, 
    7.663686e-06, 7.663698e-06, 7.663673e-06, 7.663682e-06, 7.663662e-06, 
    7.663675e-06, 7.66366e-06, 7.663662e-06, 7.663654e-06, 7.663657e-06, 
    7.663646e-06, 7.663653e-06, 7.66364e-06, 7.663647e-06, 7.663646e-06, 
    7.663653e-06, 7.663695e-06, 7.663688e-06, 7.663696e-06, 7.663695e-06, 
    7.663695e-06, 7.663702e-06, 7.663704e-06, 7.663711e-06, 7.66371e-06, 
    7.663705e-06, 7.663694e-06, 7.663698e-06, 7.663689e-06, 7.663689e-06, 
    7.663679e-06, 7.663683e-06, 7.663666e-06, 7.663671e-06, 7.663657e-06, 
    7.66366e-06, 7.663657e-06, 7.663658e-06, 7.663657e-06, 7.663662e-06, 
    7.66366e-06, 7.663664e-06, 7.663682e-06, 7.663677e-06, 7.663692e-06, 
    7.663702e-06, 7.663709e-06, 7.663713e-06, 7.663712e-06, 7.663712e-06, 
    7.663705e-06, 7.663699e-06, 7.663695e-06, 7.663692e-06, 7.663689e-06, 
    7.66368e-06, 7.663675e-06, 7.663665e-06, 7.663667e-06, 7.663663e-06, 
    7.663661e-06, 7.663655e-06, 7.663656e-06, 7.663654e-06, 7.663663e-06, 
    7.663657e-06, 7.663668e-06, 7.663665e-06, 7.663688e-06, 7.663697e-06, 
    7.663701e-06, 7.663704e-06, 7.663712e-06, 7.663706e-06, 7.663709e-06, 
    7.663703e-06, 7.6637e-06, 7.663702e-06, 7.663692e-06, 7.663696e-06, 
    7.663675e-06, 7.663684e-06, 7.663661e-06, 7.663666e-06, 7.66366e-06, 
    7.663663e-06, 7.663657e-06, 7.663662e-06, 7.663653e-06, 7.663652e-06, 
    7.663652e-06, 7.663647e-06, 7.663662e-06, 7.663657e-06, 7.663702e-06, 
    7.663702e-06, 7.663701e-06, 7.663706e-06, 7.663706e-06, 7.663712e-06, 
    7.663707e-06, 7.663705e-06, 7.6637e-06, 7.663697e-06, 7.663694e-06, 
    7.663689e-06, 7.663682e-06, 7.663672e-06, 7.663666e-06, 7.663662e-06, 
    7.663664e-06, 7.663662e-06, 7.663664e-06, 7.663666e-06, 7.663652e-06, 
    7.66366e-06, 7.663648e-06, 7.663649e-06, 7.663654e-06, 7.663649e-06, 
    7.663702e-06, 7.663703e-06, 7.663708e-06, 7.663704e-06, 7.663712e-06, 
    7.663707e-06, 7.663705e-06, 7.663695e-06, 7.663693e-06, 7.663692e-06, 
    7.663688e-06, 7.663683e-06, 7.663674e-06, 7.663667e-06, 7.663661e-06, 
    7.663661e-06, 7.663661e-06, 7.663659e-06, 7.663662e-06, 7.663659e-06, 
    7.663658e-06, 7.66366e-06, 7.663649e-06, 7.663652e-06, 7.663649e-06, 
    7.663651e-06, 7.663702e-06, 7.6637e-06, 7.663702e-06, 7.663699e-06, 
    7.663701e-06, 7.663692e-06, 7.66369e-06, 7.663678e-06, 7.663683e-06, 
    7.663675e-06, 7.663682e-06, 7.663682e-06, 7.663675e-06, 7.663682e-06, 
    7.663668e-06, 7.663677e-06, 7.663659e-06, 7.663669e-06, 7.663659e-06, 
    7.663661e-06, 7.663657e-06, 7.663654e-06, 7.663651e-06, 7.663644e-06, 
    7.663646e-06, 7.663641e-06, 7.663696e-06, 7.663692e-06, 7.663693e-06, 
    7.66369e-06, 7.663687e-06, 7.663682e-06, 7.663672e-06, 7.663676e-06, 
    7.66367e-06, 7.663668e-06, 7.663678e-06, 7.663672e-06, 7.663691e-06, 
    7.663687e-06, 7.663689e-06, 7.663696e-06, 7.663675e-06, 7.663685e-06, 
    7.663666e-06, 7.663672e-06, 7.663655e-06, 7.663663e-06, 7.663647e-06, 
    7.66364e-06, 7.663633e-06, 7.663625e-06, 7.663691e-06, 7.663693e-06, 
    7.663689e-06, 7.663683e-06, 7.663678e-06, 7.663672e-06, 7.663671e-06, 
    7.66367e-06, 7.663666e-06, 7.663663e-06, 7.663669e-06, 7.663662e-06, 
    7.663687e-06, 7.663674e-06, 7.663694e-06, 7.663688e-06, 7.663683e-06, 
    7.663685e-06, 7.663676e-06, 7.663674e-06, 7.663665e-06, 7.66367e-06, 
    7.663642e-06, 7.663654e-06, 7.66362e-06, 7.663629e-06, 7.663694e-06, 
    7.663691e-06, 7.663681e-06, 7.663685e-06, 7.663671e-06, 7.663667e-06, 
    7.663664e-06, 7.663661e-06, 7.663661e-06, 7.663658e-06, 7.663662e-06, 
    7.663658e-06, 7.663672e-06, 7.663665e-06, 7.663682e-06, 7.663678e-06, 
    7.66368e-06, 7.663682e-06, 7.663675e-06, 7.663669e-06, 7.663669e-06, 
    7.663667e-06, 7.663661e-06, 7.663671e-06, 7.66364e-06, 7.663659e-06, 
    7.663688e-06, 7.663682e-06, 7.663681e-06, 7.663683e-06, 7.663668e-06, 
    7.663673e-06, 7.663658e-06, 7.663662e-06, 7.663656e-06, 7.663659e-06, 
    7.66366e-06, 7.663663e-06, 7.663666e-06, 7.663673e-06, 7.663679e-06, 
    7.663682e-06, 7.663682e-06, 7.663677e-06, 7.663669e-06, 7.663661e-06, 
    7.663662e-06, 7.663656e-06, 7.663672e-06, 7.663665e-06, 7.663668e-06, 
    7.663662e-06, 7.663676e-06, 7.663663e-06, 7.663679e-06, 7.663678e-06, 
    7.663673e-06, 7.663665e-06, 7.663663e-06, 7.663661e-06, 7.663662e-06, 
    7.663668e-06, 7.663669e-06, 7.663673e-06, 7.663674e-06, 7.663678e-06, 
    7.663681e-06, 7.663678e-06, 7.663675e-06, 7.663668e-06, 7.663662e-06, 
    7.663654e-06, 7.663652e-06, 7.663644e-06, 7.663652e-06, 7.66364e-06, 
    7.66365e-06, 7.663632e-06, 7.663662e-06, 7.66365e-06, 7.663673e-06, 
    7.663671e-06, 7.663666e-06, 7.663655e-06, 7.663662e-06, 7.663654e-06, 
    7.663669e-06, 7.663677e-06, 7.663679e-06, 7.663682e-06, 7.663679e-06, 
    7.663679e-06, 7.663675e-06, 7.663677e-06, 7.663668e-06, 7.663672e-06, 
    7.66366e-06, 7.663654e-06, 7.663642e-06, 7.663632e-06, 7.663624e-06, 
    7.663621e-06, 7.66362e-06, 7.663619e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.325308e-14, 5.339687e-14, 5.336894e-14, 5.34848e-14, 5.342056e-14, 
    5.34964e-14, 5.328226e-14, 5.340255e-14, 5.332579e-14, 5.326606e-14, 
    5.370932e-14, 5.348997e-14, 5.393699e-14, 5.379734e-14, 5.41479e-14, 
    5.391524e-14, 5.419478e-14, 5.414124e-14, 5.430243e-14, 5.425628e-14, 
    5.446213e-14, 5.432373e-14, 5.456879e-14, 5.442912e-14, 5.445096e-14, 
    5.431915e-14, 5.353419e-14, 5.368202e-14, 5.352542e-14, 5.354651e-14, 
    5.353706e-14, 5.342187e-14, 5.336376e-14, 5.324212e-14, 5.326421e-14, 
    5.335357e-14, 5.3556e-14, 5.348735e-14, 5.366039e-14, 5.365648e-14, 
    5.384884e-14, 5.376214e-14, 5.408506e-14, 5.399339e-14, 5.425821e-14, 
    5.419164e-14, 5.425507e-14, 5.423584e-14, 5.425532e-14, 5.415769e-14, 
    5.419952e-14, 5.411359e-14, 5.377838e-14, 5.387697e-14, 5.358267e-14, 
    5.340533e-14, 5.328753e-14, 5.320385e-14, 5.321568e-14, 5.323823e-14, 
    5.335409e-14, 5.346298e-14, 5.35459e-14, 5.360133e-14, 5.365592e-14, 
    5.382092e-14, 5.390828e-14, 5.410357e-14, 5.406838e-14, 5.412801e-14, 
    5.418502e-14, 5.428062e-14, 5.426489e-14, 5.430698e-14, 5.412647e-14, 
    5.424645e-14, 5.404835e-14, 5.410254e-14, 5.36706e-14, 5.350588e-14, 
    5.343567e-14, 5.33743e-14, 5.322478e-14, 5.332804e-14, 5.328734e-14, 
    5.338419e-14, 5.344567e-14, 5.341527e-14, 5.360284e-14, 5.352994e-14, 
    5.391346e-14, 5.37484e-14, 5.417837e-14, 5.407561e-14, 5.4203e-14, 
    5.413802e-14, 5.424933e-14, 5.414915e-14, 5.432266e-14, 5.436039e-14, 
    5.43346e-14, 5.443368e-14, 5.414359e-14, 5.425506e-14, 5.341442e-14, 
    5.341937e-14, 5.344248e-14, 5.334086e-14, 5.333465e-14, 5.32415e-14, 
    5.33244e-14, 5.335968e-14, 5.344925e-14, 5.350217e-14, 5.355248e-14, 
    5.366301e-14, 5.378633e-14, 5.395862e-14, 5.408227e-14, 5.41651e-14, 
    5.411432e-14, 5.415915e-14, 5.410903e-14, 5.408554e-14, 5.434624e-14, 
    5.41999e-14, 5.441944e-14, 5.44073e-14, 5.430797e-14, 5.440867e-14, 
    5.342286e-14, 5.339432e-14, 5.329516e-14, 5.337277e-14, 5.323136e-14, 
    5.331051e-14, 5.335599e-14, 5.353143e-14, 5.356999e-14, 5.360568e-14, 
    5.367618e-14, 5.376658e-14, 5.392502e-14, 5.406271e-14, 5.418834e-14, 
    5.417914e-14, 5.418238e-14, 5.421041e-14, 5.414094e-14, 5.422182e-14, 
    5.423537e-14, 5.419991e-14, 5.440568e-14, 5.434692e-14, 5.440705e-14, 
    5.43688e-14, 5.34036e-14, 5.345161e-14, 5.342567e-14, 5.347445e-14, 
    5.344007e-14, 5.359281e-14, 5.363856e-14, 5.385252e-14, 5.376479e-14, 
    5.390443e-14, 5.3779e-14, 5.380122e-14, 5.390892e-14, 5.378579e-14, 
    5.405509e-14, 5.387252e-14, 5.42115e-14, 5.402933e-14, 5.422291e-14, 
    5.41878e-14, 5.424594e-14, 5.429798e-14, 5.436344e-14, 5.448409e-14, 
    5.445617e-14, 5.455704e-14, 5.352318e-14, 5.358538e-14, 5.357994e-14, 
    5.364503e-14, 5.369314e-14, 5.37974e-14, 5.396441e-14, 5.390164e-14, 
    5.401689e-14, 5.404e-14, 5.386492e-14, 5.397242e-14, 5.362702e-14, 
    5.368285e-14, 5.364964e-14, 5.352807e-14, 5.391607e-14, 5.371706e-14, 
    5.40843e-14, 5.397671e-14, 5.429055e-14, 5.413452e-14, 5.444079e-14, 
    5.457142e-14, 5.469439e-14, 5.483777e-14, 5.361935e-14, 5.357709e-14, 
    5.365277e-14, 5.375736e-14, 5.38544e-14, 5.398327e-14, 5.399646e-14, 
    5.402058e-14, 5.408304e-14, 5.413554e-14, 5.402817e-14, 5.41487e-14, 
    5.369574e-14, 5.393334e-14, 5.356109e-14, 5.367325e-14, 5.375121e-14, 
    5.371704e-14, 5.389447e-14, 5.393625e-14, 5.410582e-14, 5.401822e-14, 
    5.453916e-14, 5.430892e-14, 5.494694e-14, 5.476894e-14, 5.356232e-14, 
    5.361922e-14, 5.381702e-14, 5.372295e-14, 5.399188e-14, 5.405795e-14, 
    5.411169e-14, 5.418031e-14, 5.418774e-14, 5.422837e-14, 5.416177e-14, 
    5.422576e-14, 5.398354e-14, 5.409183e-14, 5.379446e-14, 5.386689e-14, 
    5.383359e-14, 5.379702e-14, 5.390983e-14, 5.402986e-14, 5.403247e-14, 
    5.40709e-14, 5.417911e-14, 5.399297e-14, 5.456876e-14, 5.421336e-14, 
    5.368124e-14, 5.379065e-14, 5.380633e-14, 5.376395e-14, 5.405136e-14, 
    5.394728e-14, 5.422739e-14, 5.415175e-14, 5.427568e-14, 5.42141e-14, 
    5.420504e-14, 5.412592e-14, 5.407663e-14, 5.395205e-14, 5.385059e-14, 
    5.37701e-14, 5.378882e-14, 5.387722e-14, 5.403721e-14, 5.418839e-14, 
    5.415527e-14, 5.426626e-14, 5.39724e-14, 5.409566e-14, 5.404803e-14, 
    5.417223e-14, 5.389996e-14, 5.41317e-14, 5.384064e-14, 5.38662e-14, 
    5.394522e-14, 5.410398e-14, 5.413916e-14, 5.417663e-14, 5.415352e-14, 
    5.404127e-14, 5.402289e-14, 5.394331e-14, 5.39213e-14, 5.386064e-14, 
    5.381036e-14, 5.385628e-14, 5.390448e-14, 5.404135e-14, 5.416451e-14, 
    5.429871e-14, 5.433155e-14, 5.448801e-14, 5.436059e-14, 5.457072e-14, 
    5.439199e-14, 5.470129e-14, 5.414519e-14, 5.438683e-14, 5.394883e-14, 
    5.39961e-14, 5.408147e-14, 5.427726e-14, 5.417165e-14, 5.429517e-14, 
    5.402218e-14, 5.388025e-14, 5.384356e-14, 5.377499e-14, 5.384513e-14, 
    5.383943e-14, 5.390651e-14, 5.388496e-14, 5.404589e-14, 5.395947e-14, 
    5.42048e-14, 5.429421e-14, 5.454645e-14, 5.470081e-14, 5.485782e-14, 
    5.492705e-14, 5.494812e-14, 5.495692e-14 ;

 LITTERC =
  5.976202e-05, 5.976187e-05, 5.97619e-05, 5.976178e-05, 5.976185e-05, 
    5.976177e-05, 5.976199e-05, 5.976186e-05, 5.976194e-05, 5.9762e-05, 
    5.976155e-05, 5.976178e-05, 5.976132e-05, 5.976146e-05, 5.976111e-05, 
    5.976134e-05, 5.976106e-05, 5.976111e-05, 5.976095e-05, 5.9761e-05, 
    5.976079e-05, 5.976093e-05, 5.976068e-05, 5.976082e-05, 5.97608e-05, 
    5.976094e-05, 5.976173e-05, 5.976158e-05, 5.976174e-05, 5.976172e-05, 
    5.976173e-05, 5.976185e-05, 5.97619e-05, 5.976203e-05, 5.976201e-05, 
    5.976191e-05, 5.976171e-05, 5.976178e-05, 5.97616e-05, 5.976161e-05, 
    5.976141e-05, 5.97615e-05, 5.976117e-05, 5.976126e-05, 5.9761e-05, 
    5.976106e-05, 5.9761e-05, 5.976102e-05, 5.9761e-05, 5.97611e-05, 
    5.976106e-05, 5.976114e-05, 5.976148e-05, 5.976138e-05, 5.976168e-05, 
    5.976186e-05, 5.976198e-05, 5.976206e-05, 5.976205e-05, 5.976203e-05, 
    5.976191e-05, 5.97618e-05, 5.976172e-05, 5.976166e-05, 5.976161e-05, 
    5.976144e-05, 5.976135e-05, 5.976115e-05, 5.976119e-05, 5.976113e-05, 
    5.976107e-05, 5.976097e-05, 5.976099e-05, 5.976095e-05, 5.976113e-05, 
    5.976101e-05, 5.976121e-05, 5.976115e-05, 5.976159e-05, 5.976176e-05, 
    5.976183e-05, 5.976189e-05, 5.976205e-05, 5.976194e-05, 5.976198e-05, 
    5.976188e-05, 5.976182e-05, 5.976185e-05, 5.976166e-05, 5.976174e-05, 
    5.976135e-05, 5.976151e-05, 5.976108e-05, 5.976118e-05, 5.976105e-05, 
    5.976112e-05, 5.976101e-05, 5.976111e-05, 5.976093e-05, 5.976089e-05, 
    5.976092e-05, 5.976082e-05, 5.976111e-05, 5.9761e-05, 5.976185e-05, 
    5.976185e-05, 5.976182e-05, 5.976193e-05, 5.976193e-05, 5.976203e-05, 
    5.976194e-05, 5.976191e-05, 5.976182e-05, 5.976176e-05, 5.976171e-05, 
    5.97616e-05, 5.976147e-05, 5.97613e-05, 5.976118e-05, 5.976109e-05, 
    5.976114e-05, 5.97611e-05, 5.976115e-05, 5.976117e-05, 5.976091e-05, 
    5.976106e-05, 5.976083e-05, 5.976085e-05, 5.976095e-05, 5.976085e-05, 
    5.976184e-05, 5.976187e-05, 5.976197e-05, 5.976189e-05, 5.976204e-05, 
    5.976196e-05, 5.976191e-05, 5.976173e-05, 5.976169e-05, 5.976166e-05, 
    5.976159e-05, 5.97615e-05, 5.976133e-05, 5.976119e-05, 5.976107e-05, 
    5.976108e-05, 5.976107e-05, 5.976105e-05, 5.976111e-05, 5.976103e-05, 
    5.976102e-05, 5.976106e-05, 5.976085e-05, 5.976091e-05, 5.976085e-05, 
    5.976089e-05, 5.976186e-05, 5.976181e-05, 5.976184e-05, 5.976179e-05, 
    5.976183e-05, 5.976167e-05, 5.976162e-05, 5.976141e-05, 5.97615e-05, 
    5.976135e-05, 5.976148e-05, 5.976146e-05, 5.976135e-05, 5.976147e-05, 
    5.97612e-05, 5.976139e-05, 5.976105e-05, 5.976123e-05, 5.976103e-05, 
    5.976107e-05, 5.976101e-05, 5.976096e-05, 5.976089e-05, 5.976077e-05, 
    5.97608e-05, 5.976069e-05, 5.976174e-05, 5.976168e-05, 5.976169e-05, 
    5.976162e-05, 5.976157e-05, 5.976146e-05, 5.976129e-05, 5.976136e-05, 
    5.976124e-05, 5.976122e-05, 5.976139e-05, 5.976129e-05, 5.976163e-05, 
    5.976158e-05, 5.976161e-05, 5.976174e-05, 5.976134e-05, 5.976154e-05, 
    5.976117e-05, 5.976128e-05, 5.976097e-05, 5.976112e-05, 5.976081e-05, 
    5.976068e-05, 5.976055e-05, 5.976041e-05, 5.976165e-05, 5.976169e-05, 
    5.976161e-05, 5.97615e-05, 5.976141e-05, 5.976127e-05, 5.976126e-05, 
    5.976124e-05, 5.976117e-05, 5.976112e-05, 5.976123e-05, 5.976111e-05, 
    5.976157e-05, 5.976133e-05, 5.97617e-05, 5.976159e-05, 5.976151e-05, 
    5.976154e-05, 5.976137e-05, 5.976132e-05, 5.976115e-05, 5.976124e-05, 
    5.976071e-05, 5.976095e-05, 5.97603e-05, 5.976048e-05, 5.97617e-05, 
    5.976165e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 5.97612e-05, 
    5.976114e-05, 5.976107e-05, 5.976107e-05, 5.976103e-05, 5.97611e-05, 
    5.976103e-05, 5.976127e-05, 5.976117e-05, 5.976147e-05, 5.976139e-05, 
    5.976143e-05, 5.976146e-05, 5.976135e-05, 5.976123e-05, 5.976123e-05, 
    5.976119e-05, 5.976108e-05, 5.976127e-05, 5.976068e-05, 5.976104e-05, 
    5.976158e-05, 5.976147e-05, 5.976146e-05, 5.97615e-05, 5.976121e-05, 
    5.976131e-05, 5.976103e-05, 5.97611e-05, 5.976098e-05, 5.976104e-05, 
    5.976105e-05, 5.976113e-05, 5.976118e-05, 5.976131e-05, 5.976141e-05, 
    5.976149e-05, 5.976147e-05, 5.976138e-05, 5.976122e-05, 5.976107e-05, 
    5.97611e-05, 5.976099e-05, 5.976129e-05, 5.976116e-05, 5.976121e-05, 
    5.976109e-05, 5.976136e-05, 5.976113e-05, 5.976142e-05, 5.976139e-05, 
    5.976131e-05, 5.976115e-05, 5.976112e-05, 5.976108e-05, 5.97611e-05, 
    5.976122e-05, 5.976123e-05, 5.976131e-05, 5.976134e-05, 5.97614e-05, 
    5.976145e-05, 5.976141e-05, 5.976135e-05, 5.976122e-05, 5.976109e-05, 
    5.976095e-05, 5.976092e-05, 5.976076e-05, 5.976089e-05, 5.976068e-05, 
    5.976086e-05, 5.976055e-05, 5.976111e-05, 5.976087e-05, 5.976131e-05, 
    5.976126e-05, 5.976118e-05, 5.976098e-05, 5.976109e-05, 5.976096e-05, 
    5.976123e-05, 5.976138e-05, 5.976142e-05, 5.976149e-05, 5.976142e-05, 
    5.976142e-05, 5.976135e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976105e-05, 5.976096e-05, 5.97607e-05, 5.976055e-05, 5.976039e-05, 
    5.976032e-05, 5.97603e-05, 5.976029e-05 ;

 LITTERC_HR =
  8.591897e-13, 8.615078e-13, 8.610575e-13, 8.629254e-13, 8.618897e-13, 
    8.631123e-13, 8.596602e-13, 8.615995e-13, 8.603619e-13, 8.593989e-13, 
    8.66545e-13, 8.630088e-13, 8.702151e-13, 8.679639e-13, 8.736153e-13, 
    8.698645e-13, 8.743711e-13, 8.735079e-13, 8.761065e-13, 8.753624e-13, 
    8.78681e-13, 8.764498e-13, 8.804005e-13, 8.781488e-13, 8.785009e-13, 
    8.76376e-13, 8.637216e-13, 8.661048e-13, 8.635801e-13, 8.639202e-13, 
    8.637678e-13, 8.619109e-13, 8.60974e-13, 8.590129e-13, 8.593692e-13, 
    8.608098e-13, 8.640731e-13, 8.629664e-13, 8.65756e-13, 8.656931e-13, 
    8.687941e-13, 8.673965e-13, 8.726022e-13, 8.711244e-13, 8.753935e-13, 
    8.743204e-13, 8.75343e-13, 8.750331e-13, 8.75347e-13, 8.737731e-13, 
    8.744475e-13, 8.730623e-13, 8.676582e-13, 8.692477e-13, 8.645031e-13, 
    8.616442e-13, 8.597451e-13, 8.58396e-13, 8.585868e-13, 8.589503e-13, 
    8.608182e-13, 8.625737e-13, 8.639103e-13, 8.648039e-13, 8.65684e-13, 
    8.683441e-13, 8.697523e-13, 8.729006e-13, 8.723333e-13, 8.732947e-13, 
    8.742137e-13, 8.757548e-13, 8.755013e-13, 8.761798e-13, 8.732698e-13, 
    8.75204e-13, 8.720105e-13, 8.72884e-13, 8.659207e-13, 8.632651e-13, 
    8.621332e-13, 8.611439e-13, 8.587334e-13, 8.603982e-13, 8.59742e-13, 
    8.613034e-13, 8.622946e-13, 8.618045e-13, 8.648283e-13, 8.636531e-13, 
    8.698358e-13, 8.671749e-13, 8.741065e-13, 8.724498e-13, 8.745035e-13, 
    8.734559e-13, 8.752503e-13, 8.736355e-13, 8.764325e-13, 8.770408e-13, 
    8.766251e-13, 8.782224e-13, 8.735458e-13, 8.753427e-13, 8.617907e-13, 
    8.618706e-13, 8.622432e-13, 8.606048e-13, 8.605048e-13, 8.59003e-13, 
    8.603395e-13, 8.609082e-13, 8.623522e-13, 8.632054e-13, 8.640164e-13, 
    8.657984e-13, 8.677864e-13, 8.70564e-13, 8.725572e-13, 8.738925e-13, 
    8.73074e-13, 8.737966e-13, 8.729887e-13, 8.7261e-13, 8.768127e-13, 
    8.744536e-13, 8.779927e-13, 8.777971e-13, 8.761959e-13, 8.778192e-13, 
    8.619267e-13, 8.614667e-13, 8.598681e-13, 8.611192e-13, 8.588395e-13, 
    8.601155e-13, 8.608488e-13, 8.636771e-13, 8.642987e-13, 8.648741e-13, 
    8.660106e-13, 8.67468e-13, 8.700222e-13, 8.72242e-13, 8.742672e-13, 
    8.74119e-13, 8.741711e-13, 8.746231e-13, 8.735031e-13, 8.748069e-13, 
    8.750254e-13, 8.744537e-13, 8.777709e-13, 8.768238e-13, 8.77793e-13, 
    8.771764e-13, 8.616163e-13, 8.623903e-13, 8.619721e-13, 8.627584e-13, 
    8.622042e-13, 8.646666e-13, 8.654043e-13, 8.688535e-13, 8.674392e-13, 
    8.696903e-13, 8.676682e-13, 8.680265e-13, 8.697626e-13, 8.677777e-13, 
    8.721191e-13, 8.691759e-13, 8.746406e-13, 8.717039e-13, 8.748245e-13, 
    8.742585e-13, 8.751958e-13, 8.760347e-13, 8.7709e-13, 8.79035e-13, 
    8.785849e-13, 8.802109e-13, 8.63544e-13, 8.645469e-13, 8.644591e-13, 
    8.655085e-13, 8.66284e-13, 8.679648e-13, 8.706572e-13, 8.696453e-13, 
    8.715032e-13, 8.718759e-13, 8.690534e-13, 8.707863e-13, 8.652181e-13, 
    8.661182e-13, 8.655827e-13, 8.636229e-13, 8.698778e-13, 8.666697e-13, 
    8.725901e-13, 8.708555e-13, 8.75915e-13, 8.733995e-13, 8.783369e-13, 
    8.804428e-13, 8.824252e-13, 8.847366e-13, 8.650945e-13, 8.644133e-13, 
    8.656333e-13, 8.673193e-13, 8.688838e-13, 8.709612e-13, 8.71174e-13, 
    8.715628e-13, 8.725696e-13, 8.73416e-13, 8.716852e-13, 8.736282e-13, 
    8.663259e-13, 8.701563e-13, 8.641552e-13, 8.659634e-13, 8.672201e-13, 
    8.666694e-13, 8.695298e-13, 8.702032e-13, 8.729369e-13, 8.715247e-13, 
    8.799228e-13, 8.762111e-13, 8.864965e-13, 8.83627e-13, 8.641751e-13, 
    8.650924e-13, 8.682811e-13, 8.667646e-13, 8.711001e-13, 8.721653e-13, 
    8.730316e-13, 8.741377e-13, 8.742575e-13, 8.749126e-13, 8.738389e-13, 
    8.748704e-13, 8.709657e-13, 8.727113e-13, 8.679175e-13, 8.690851e-13, 
    8.685482e-13, 8.679588e-13, 8.697773e-13, 8.717123e-13, 8.717544e-13, 
    8.723739e-13, 8.741185e-13, 8.711177e-13, 8.803999e-13, 8.746705e-13, 
    8.660921e-13, 8.67856e-13, 8.681088e-13, 8.674256e-13, 8.720589e-13, 
    8.703811e-13, 8.748967e-13, 8.736773e-13, 8.756752e-13, 8.746825e-13, 
    8.745364e-13, 8.73261e-13, 8.724663e-13, 8.704579e-13, 8.688223e-13, 
    8.675248e-13, 8.678266e-13, 8.692517e-13, 8.718308e-13, 8.742679e-13, 
    8.737341e-13, 8.755234e-13, 8.70786e-13, 8.727731e-13, 8.720053e-13, 
    8.740076e-13, 8.696182e-13, 8.733541e-13, 8.686619e-13, 8.690739e-13, 
    8.703478e-13, 8.729073e-13, 8.734744e-13, 8.740784e-13, 8.737059e-13, 
    8.718964e-13, 8.716e-13, 8.703171e-13, 8.699623e-13, 8.689842e-13, 
    8.681738e-13, 8.689141e-13, 8.696911e-13, 8.718975e-13, 8.73883e-13, 
    8.760465e-13, 8.765759e-13, 8.790982e-13, 8.77044e-13, 8.804316e-13, 
    8.775502e-13, 8.825364e-13, 8.735716e-13, 8.77467e-13, 8.70406e-13, 
    8.711681e-13, 8.725444e-13, 8.757007e-13, 8.739981e-13, 8.759895e-13, 
    8.715886e-13, 8.693005e-13, 8.68709e-13, 8.676036e-13, 8.687343e-13, 
    8.686424e-13, 8.697238e-13, 8.693764e-13, 8.719707e-13, 8.705776e-13, 
    8.745325e-13, 8.75974e-13, 8.800403e-13, 8.825286e-13, 8.850598e-13, 
    8.861758e-13, 8.865154e-13, 8.866573e-13 ;

 LITTERC_LOSS =
  1.59121e-12, 1.595503e-12, 1.594669e-12, 1.598129e-12, 1.596211e-12, 
    1.598475e-12, 1.592082e-12, 1.595673e-12, 1.593381e-12, 1.591598e-12, 
    1.604832e-12, 1.598283e-12, 1.61163e-12, 1.60746e-12, 1.617927e-12, 
    1.61098e-12, 1.619326e-12, 1.617728e-12, 1.62254e-12, 1.621162e-12, 
    1.627308e-12, 1.623176e-12, 1.630493e-12, 1.626323e-12, 1.626975e-12, 
    1.62304e-12, 1.599603e-12, 1.604017e-12, 1.599341e-12, 1.599971e-12, 
    1.599689e-12, 1.59625e-12, 1.594515e-12, 1.590883e-12, 1.591543e-12, 
    1.594211e-12, 1.600254e-12, 1.598205e-12, 1.603371e-12, 1.603255e-12, 
    1.608998e-12, 1.606409e-12, 1.61605e-12, 1.613314e-12, 1.62122e-12, 
    1.619233e-12, 1.621126e-12, 1.620552e-12, 1.621134e-12, 1.618219e-12, 
    1.619468e-12, 1.616902e-12, 1.606894e-12, 1.609838e-12, 1.601051e-12, 
    1.595756e-12, 1.592239e-12, 1.58974e-12, 1.590094e-12, 1.590767e-12, 
    1.594226e-12, 1.597477e-12, 1.599953e-12, 1.601608e-12, 1.603238e-12, 
    1.608164e-12, 1.610772e-12, 1.616603e-12, 1.615552e-12, 1.617333e-12, 
    1.619035e-12, 1.621889e-12, 1.62142e-12, 1.622676e-12, 1.617287e-12, 
    1.620869e-12, 1.614954e-12, 1.616572e-12, 1.603676e-12, 1.598758e-12, 
    1.596662e-12, 1.59483e-12, 1.590365e-12, 1.593448e-12, 1.592233e-12, 
    1.595125e-12, 1.596961e-12, 1.596053e-12, 1.601653e-12, 1.599477e-12, 
    1.610927e-12, 1.605999e-12, 1.618836e-12, 1.615768e-12, 1.619572e-12, 
    1.617631e-12, 1.620955e-12, 1.617964e-12, 1.623144e-12, 1.624271e-12, 
    1.623501e-12, 1.626459e-12, 1.617798e-12, 1.621126e-12, 1.596027e-12, 
    1.596175e-12, 1.596865e-12, 1.593831e-12, 1.593646e-12, 1.590864e-12, 
    1.59334e-12, 1.594393e-12, 1.597067e-12, 1.598647e-12, 1.600149e-12, 
    1.60345e-12, 1.607131e-12, 1.612276e-12, 1.615967e-12, 1.61844e-12, 
    1.616924e-12, 1.618262e-12, 1.616766e-12, 1.616065e-12, 1.623848e-12, 
    1.619479e-12, 1.626034e-12, 1.625671e-12, 1.622706e-12, 1.625712e-12, 
    1.596279e-12, 1.595427e-12, 1.592467e-12, 1.594784e-12, 1.590562e-12, 
    1.592925e-12, 1.594283e-12, 1.599521e-12, 1.600672e-12, 1.601738e-12, 
    1.603843e-12, 1.606542e-12, 1.611272e-12, 1.615383e-12, 1.619134e-12, 
    1.618859e-12, 1.618956e-12, 1.619793e-12, 1.617719e-12, 1.620133e-12, 
    1.620538e-12, 1.619479e-12, 1.625623e-12, 1.623869e-12, 1.625664e-12, 
    1.624522e-12, 1.595704e-12, 1.597138e-12, 1.596363e-12, 1.59782e-12, 
    1.596793e-12, 1.601353e-12, 1.60272e-12, 1.609108e-12, 1.606488e-12, 
    1.610658e-12, 1.606913e-12, 1.607576e-12, 1.610791e-12, 1.607115e-12, 
    1.615156e-12, 1.609705e-12, 1.619826e-12, 1.614387e-12, 1.620166e-12, 
    1.619118e-12, 1.620854e-12, 1.622407e-12, 1.624362e-12, 1.627964e-12, 
    1.62713e-12, 1.630142e-12, 1.599275e-12, 1.601132e-12, 1.600969e-12, 
    1.602913e-12, 1.604349e-12, 1.607462e-12, 1.612448e-12, 1.610574e-12, 
    1.614015e-12, 1.614705e-12, 1.609478e-12, 1.612687e-12, 1.602375e-12, 
    1.604042e-12, 1.60305e-12, 1.599421e-12, 1.611005e-12, 1.605063e-12, 
    1.616028e-12, 1.612815e-12, 1.622186e-12, 1.617527e-12, 1.626671e-12, 
    1.630571e-12, 1.634243e-12, 1.638524e-12, 1.602146e-12, 1.600884e-12, 
    1.603144e-12, 1.606266e-12, 1.609164e-12, 1.613011e-12, 1.613405e-12, 
    1.614125e-12, 1.61599e-12, 1.617558e-12, 1.614352e-12, 1.61795e-12, 
    1.604427e-12, 1.611521e-12, 1.600406e-12, 1.603755e-12, 1.606083e-12, 
    1.605063e-12, 1.61036e-12, 1.611607e-12, 1.61667e-12, 1.614055e-12, 
    1.629608e-12, 1.622734e-12, 1.641783e-12, 1.636469e-12, 1.600443e-12, 
    1.602142e-12, 1.608048e-12, 1.605239e-12, 1.613269e-12, 1.615241e-12, 
    1.616846e-12, 1.618894e-12, 1.619116e-12, 1.620329e-12, 1.618341e-12, 
    1.620251e-12, 1.61302e-12, 1.616252e-12, 1.607374e-12, 1.609537e-12, 
    1.608542e-12, 1.607451e-12, 1.610819e-12, 1.614402e-12, 1.61448e-12, 
    1.615628e-12, 1.618859e-12, 1.613301e-12, 1.630492e-12, 1.619881e-12, 
    1.603994e-12, 1.60726e-12, 1.607728e-12, 1.606463e-12, 1.615044e-12, 
    1.611937e-12, 1.6203e-12, 1.618042e-12, 1.621742e-12, 1.619903e-12, 
    1.619633e-12, 1.617271e-12, 1.615799e-12, 1.612079e-12, 1.60905e-12, 
    1.606647e-12, 1.607206e-12, 1.609845e-12, 1.614622e-12, 1.619135e-12, 
    1.618147e-12, 1.621461e-12, 1.612687e-12, 1.616367e-12, 1.614945e-12, 
    1.618653e-12, 1.610524e-12, 1.617443e-12, 1.608753e-12, 1.609516e-12, 
    1.611875e-12, 1.616615e-12, 1.617666e-12, 1.618784e-12, 1.618094e-12, 
    1.614743e-12, 1.614194e-12, 1.611818e-12, 1.611161e-12, 1.60935e-12, 
    1.607849e-12, 1.60922e-12, 1.610659e-12, 1.614745e-12, 1.618422e-12, 
    1.622429e-12, 1.62341e-12, 1.628081e-12, 1.624277e-12, 1.630551e-12, 
    1.625214e-12, 1.634449e-12, 1.617846e-12, 1.62506e-12, 1.611983e-12, 
    1.613394e-12, 1.615943e-12, 1.621789e-12, 1.618636e-12, 1.622324e-12, 
    1.614173e-12, 1.609935e-12, 1.60884e-12, 1.606793e-12, 1.608887e-12, 
    1.608717e-12, 1.61072e-12, 1.610076e-12, 1.614881e-12, 1.612301e-12, 
    1.619625e-12, 1.622295e-12, 1.629826e-12, 1.634434e-12, 1.639122e-12, 
    1.641189e-12, 1.641818e-12, 1.642081e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  3.91629e-18, 3.914856e-18, 3.915128e-18, 3.913988e-18, 3.91461e-18, 
    3.913871e-18, 3.915987e-18, 3.91481e-18, 3.915554e-18, 3.916144e-18, 
    3.911814e-18, 3.913934e-18, 3.909504e-18, 3.91087e-18, 3.907406e-18, 
    3.909732e-18, 3.906933e-18, 3.907446e-18, 3.905837e-18, 3.906296e-18, 
    3.904299e-18, 3.905625e-18, 3.903221e-18, 3.904601e-18, 3.904395e-18, 
    3.905673e-18, 3.913481e-18, 3.912086e-18, 3.91357e-18, 3.913369e-18, 
    3.913454e-18, 3.914607e-18, 3.915207e-18, 3.91638e-18, 3.916163e-18, 
    3.91529e-18, 3.913279e-18, 3.913943e-18, 3.912217e-18, 3.912255e-18, 
    3.910355e-18, 3.911212e-18, 3.908005e-18, 3.908909e-18, 3.906277e-18, 
    3.906942e-18, 3.906312e-18, 3.9065e-18, 3.90631e-18, 3.907284e-18, 
    3.906868e-18, 3.907717e-18, 3.911057e-18, 3.910083e-18, 3.913005e-18, 
    3.914808e-18, 3.91594e-18, 3.916765e-18, 3.916649e-18, 3.916431e-18, 
    3.915285e-18, 3.914186e-18, 3.913356e-18, 3.912806e-18, 3.912261e-18, 
    3.910682e-18, 3.909789e-18, 3.907836e-18, 3.908165e-18, 3.907589e-18, 
    3.907007e-18, 3.906062e-18, 3.906214e-18, 3.905803e-18, 3.907588e-18, 
    3.906409e-18, 3.908358e-18, 3.907827e-18, 3.912205e-18, 3.913759e-18, 
    3.9145e-18, 3.915079e-18, 3.91656e-18, 3.915543e-18, 3.915946e-18, 
    3.914967e-18, 3.914359e-18, 3.914655e-18, 3.912791e-18, 3.913519e-18, 
    3.909736e-18, 3.911363e-18, 3.907075e-18, 3.908095e-18, 3.906827e-18, 
    3.907469e-18, 3.906377e-18, 3.90736e-18, 3.905642e-18, 3.905279e-18, 
    3.90553e-18, 3.904539e-18, 3.907417e-18, 3.906321e-18, 3.914668e-18, 
    3.914621e-18, 3.914387e-18, 3.915416e-18, 3.915475e-18, 3.916391e-18, 
    3.915567e-18, 3.915224e-18, 3.914316e-18, 3.913797e-18, 3.913298e-18, 
    3.9122e-18, 3.91099e-18, 3.909275e-18, 3.90803e-18, 3.907201e-18, 
    3.907703e-18, 3.90726e-18, 3.907759e-18, 3.907988e-18, 3.905422e-18, 
    3.90687e-18, 3.904681e-18, 3.904799e-18, 3.905796e-18, 3.904786e-18, 
    3.914586e-18, 3.914864e-18, 3.915861e-18, 3.91508e-18, 3.91649e-18, 
    3.915713e-18, 3.915272e-18, 3.913524e-18, 3.913118e-18, 3.912771e-18, 
    3.912064e-18, 3.911169e-18, 3.909606e-18, 3.908234e-18, 3.906969e-18, 
    3.90706e-18, 3.907029e-18, 3.906756e-18, 3.907444e-18, 3.906643e-18, 
    3.906517e-18, 3.906859e-18, 3.904815e-18, 3.905398e-18, 3.904802e-18, 
    3.905178e-18, 3.914771e-18, 3.914298e-18, 3.914555e-18, 3.914077e-18, 
    3.914421e-18, 3.912919e-18, 3.912469e-18, 3.910342e-18, 3.911191e-18, 
    3.909814e-18, 3.911044e-18, 3.910831e-18, 3.909808e-18, 3.910972e-18, 
    3.908327e-18, 3.910153e-18, 3.906746e-18, 3.908603e-18, 3.906631e-18, 
    3.906975e-18, 3.906397e-18, 3.90589e-18, 3.905235e-18, 3.904056e-18, 
    3.904325e-18, 3.903324e-18, 3.913585e-18, 3.912982e-18, 3.913018e-18, 
    3.912374e-18, 3.911902e-18, 3.910858e-18, 3.909207e-18, 3.909822e-18, 
    3.908674e-18, 3.90845e-18, 3.910183e-18, 3.909135e-18, 3.912564e-18, 
    3.912027e-18, 3.912334e-18, 3.913547e-18, 3.909704e-18, 3.911685e-18, 
    3.908013e-18, 3.90908e-18, 3.905965e-18, 3.90753e-18, 3.904477e-18, 
    3.903219e-18, 3.901958e-18, 3.900578e-18, 3.912633e-18, 3.913045e-18, 
    3.912292e-18, 3.911283e-18, 3.910298e-18, 3.909019e-18, 3.908878e-18, 
    3.908644e-18, 3.908015e-18, 3.907495e-18, 3.908586e-18, 3.907364e-18, 
    3.911937e-18, 3.909524e-18, 3.913217e-18, 3.912127e-18, 3.911335e-18, 
    3.911665e-18, 3.909888e-18, 3.909476e-18, 3.907808e-18, 3.90866e-18, 
    3.903545e-18, 3.905807e-18, 3.899472e-18, 3.901249e-18, 3.913193e-18, 
    3.912626e-18, 3.910681e-18, 3.911604e-18, 3.908924e-18, 3.908273e-18, 
    3.907729e-18, 3.907063e-18, 3.906978e-18, 3.906582e-18, 3.907234e-18, 
    3.906601e-18, 3.909016e-18, 3.907933e-18, 3.910882e-18, 3.910174e-18, 
    3.910494e-18, 3.910858e-18, 3.909737e-18, 3.908574e-18, 3.908521e-18, 
    3.908152e-18, 3.907165e-18, 3.908912e-18, 3.903304e-18, 3.906811e-18, 
    3.91201e-18, 3.910958e-18, 3.910774e-18, 3.911187e-18, 3.908339e-18, 
    3.909374e-18, 3.906588e-18, 3.907334e-18, 3.906104e-18, 3.906717e-18, 
    3.906809e-18, 3.90759e-18, 3.908086e-18, 3.909332e-18, 3.910339e-18, 
    3.911124e-18, 3.910939e-18, 3.910076e-18, 3.908496e-18, 3.906983e-18, 
    3.907318e-18, 3.906197e-18, 3.909119e-18, 3.907907e-18, 3.908384e-18, 
    3.907135e-18, 3.909844e-18, 3.907621e-18, 3.910423e-18, 3.910171e-18, 
    3.909394e-18, 3.907844e-18, 3.907459e-18, 3.9071e-18, 3.907316e-18, 
    3.90845e-18, 3.908624e-18, 3.909406e-18, 3.909636e-18, 3.910224e-18, 
    3.910724e-18, 3.910274e-18, 3.909807e-18, 3.908439e-18, 3.907221e-18, 
    3.905887e-18, 3.90555e-18, 3.904063e-18, 3.905311e-18, 3.90329e-18, 
    3.905064e-18, 3.901965e-18, 3.907451e-18, 3.905062e-18, 3.909349e-18, 
    3.90888e-18, 3.90806e-18, 3.906126e-18, 3.90714e-18, 3.90594e-18, 
    3.908629e-18, 3.91006e-18, 3.910397e-18, 3.911081e-18, 3.910381e-18, 
    3.910436e-18, 3.909769e-18, 3.909981e-18, 3.908393e-18, 3.909245e-18, 
    3.906818e-18, 3.905942e-18, 3.903438e-18, 3.901924e-18, 3.900341e-18, 
    3.899658e-18, 3.899447e-18, 3.899361e-18 ;

 MEG_acetic_acid =
  5.874434e-19, 5.872284e-19, 5.872692e-19, 5.870982e-19, 5.871915e-19, 
    5.870807e-19, 5.87398e-19, 5.872215e-19, 5.873331e-19, 5.874216e-19, 
    5.867721e-19, 5.8709e-19, 5.864256e-19, 5.866305e-19, 5.86111e-19, 
    5.864597e-19, 5.8604e-19, 5.861169e-19, 5.858756e-19, 5.859444e-19, 
    5.856448e-19, 5.858437e-19, 5.854831e-19, 5.8569e-19, 5.856592e-19, 
    5.85851e-19, 5.870221e-19, 5.868129e-19, 5.870354e-19, 5.870054e-19, 
    5.87018e-19, 5.87191e-19, 5.87281e-19, 5.874571e-19, 5.874243e-19, 
    5.872934e-19, 5.869918e-19, 5.870914e-19, 5.868325e-19, 5.868382e-19, 
    5.865533e-19, 5.866818e-19, 5.862007e-19, 5.863364e-19, 5.859415e-19, 
    5.860413e-19, 5.859468e-19, 5.85975e-19, 5.859465e-19, 5.860926e-19, 
    5.860302e-19, 5.861576e-19, 5.866585e-19, 5.865124e-19, 5.869508e-19, 
    5.872212e-19, 5.87391e-19, 5.875147e-19, 5.874972e-19, 5.874647e-19, 
    5.872928e-19, 5.871278e-19, 5.870034e-19, 5.869209e-19, 5.868391e-19, 
    5.866024e-19, 5.864683e-19, 5.861753e-19, 5.862247e-19, 5.861384e-19, 
    5.86051e-19, 5.859092e-19, 5.85932e-19, 5.858704e-19, 5.861381e-19, 
    5.859614e-19, 5.862537e-19, 5.861741e-19, 5.868307e-19, 5.870638e-19, 
    5.87175e-19, 5.872618e-19, 5.87484e-19, 5.873314e-19, 5.873919e-19, 
    5.87245e-19, 5.871538e-19, 5.871983e-19, 5.869187e-19, 5.870279e-19, 
    5.864604e-19, 5.867044e-19, 5.860612e-19, 5.862143e-19, 5.860241e-19, 
    5.861204e-19, 5.859564e-19, 5.861039e-19, 5.858464e-19, 5.857919e-19, 
    5.858294e-19, 5.856808e-19, 5.861125e-19, 5.859482e-19, 5.872002e-19, 
    5.871931e-19, 5.87158e-19, 5.873125e-19, 5.873212e-19, 5.874587e-19, 
    5.87335e-19, 5.872836e-19, 5.871474e-19, 5.870696e-19, 5.869946e-19, 
    5.868299e-19, 5.866485e-19, 5.863912e-19, 5.862045e-19, 5.860801e-19, 
    5.861554e-19, 5.860891e-19, 5.861638e-19, 5.861982e-19, 5.858132e-19, 
    5.860304e-19, 5.857022e-19, 5.857198e-19, 5.858694e-19, 5.857179e-19, 
    5.871878e-19, 5.872295e-19, 5.873791e-19, 5.87262e-19, 5.874735e-19, 
    5.873569e-19, 5.872908e-19, 5.870286e-19, 5.869677e-19, 5.869156e-19, 
    5.868096e-19, 5.866753e-19, 5.864409e-19, 5.86235e-19, 5.860454e-19, 
    5.86059e-19, 5.860543e-19, 5.860134e-19, 5.861167e-19, 5.859964e-19, 
    5.859775e-19, 5.860289e-19, 5.857223e-19, 5.858096e-19, 5.857202e-19, 
    5.857767e-19, 5.872156e-19, 5.871447e-19, 5.871832e-19, 5.871116e-19, 
    5.871631e-19, 5.869378e-19, 5.868704e-19, 5.865513e-19, 5.866787e-19, 
    5.864721e-19, 5.866566e-19, 5.866247e-19, 5.864712e-19, 5.866457e-19, 
    5.86249e-19, 5.86523e-19, 5.860119e-19, 5.862905e-19, 5.859947e-19, 
    5.860462e-19, 5.859595e-19, 5.858835e-19, 5.857853e-19, 5.856083e-19, 
    5.856487e-19, 5.854986e-19, 5.870378e-19, 5.869472e-19, 5.869526e-19, 
    5.868561e-19, 5.867852e-19, 5.866287e-19, 5.86381e-19, 5.864732e-19, 
    5.863011e-19, 5.862675e-19, 5.865275e-19, 5.863702e-19, 5.868846e-19, 
    5.868041e-19, 5.868502e-19, 5.870321e-19, 5.864556e-19, 5.867527e-19, 
    5.862019e-19, 5.86362e-19, 5.858947e-19, 5.861295e-19, 5.856715e-19, 
    5.854829e-19, 5.852936e-19, 5.850867e-19, 5.86895e-19, 5.869568e-19, 
    5.868438e-19, 5.866924e-19, 5.865447e-19, 5.863528e-19, 5.863317e-19, 
    5.862965e-19, 5.862022e-19, 5.861243e-19, 5.862879e-19, 5.861046e-19, 
    5.867906e-19, 5.864286e-19, 5.869825e-19, 5.86819e-19, 5.867002e-19, 
    5.867497e-19, 5.864832e-19, 5.864213e-19, 5.861712e-19, 5.86299e-19, 
    5.855317e-19, 5.85871e-19, 5.849208e-19, 5.851874e-19, 5.86979e-19, 
    5.86894e-19, 5.866021e-19, 5.867405e-19, 5.863386e-19, 5.862409e-19, 
    5.861594e-19, 5.860594e-19, 5.860467e-19, 5.859872e-19, 5.860851e-19, 
    5.859901e-19, 5.863524e-19, 5.8619e-19, 5.866324e-19, 5.865261e-19, 
    5.865741e-19, 5.866286e-19, 5.864606e-19, 5.86286e-19, 5.862781e-19, 
    5.862228e-19, 5.860747e-19, 5.863368e-19, 5.854955e-19, 5.860216e-19, 
    5.868015e-19, 5.866437e-19, 5.866161e-19, 5.866781e-19, 5.862509e-19, 
    5.864061e-19, 5.859881e-19, 5.861e-19, 5.859156e-19, 5.860076e-19, 
    5.860213e-19, 5.861386e-19, 5.862128e-19, 5.863997e-19, 5.865508e-19, 
    5.866685e-19, 5.866408e-19, 5.865114e-19, 5.862743e-19, 5.860475e-19, 
    5.860977e-19, 5.859296e-19, 5.863678e-19, 5.86186e-19, 5.862576e-19, 
    5.860702e-19, 5.864766e-19, 5.861431e-19, 5.865634e-19, 5.865257e-19, 
    5.864091e-19, 5.861765e-19, 5.861189e-19, 5.860649e-19, 5.860974e-19, 
    5.862675e-19, 5.862936e-19, 5.864109e-19, 5.864454e-19, 5.865336e-19, 
    5.866086e-19, 5.865411e-19, 5.864711e-19, 5.862658e-19, 5.860832e-19, 
    5.85883e-19, 5.858324e-19, 5.856093e-19, 5.857966e-19, 5.854934e-19, 
    5.857596e-19, 5.852948e-19, 5.861175e-19, 5.857593e-19, 5.864024e-19, 
    5.86332e-19, 5.86209e-19, 5.859188e-19, 5.860711e-19, 5.85891e-19, 
    5.862943e-19, 5.86509e-19, 5.865595e-19, 5.866621e-19, 5.865571e-19, 
    5.865655e-19, 5.864653e-19, 5.864972e-19, 5.862589e-19, 5.863867e-19, 
    5.860228e-19, 5.858914e-19, 5.855158e-19, 5.852887e-19, 5.850512e-19, 
    5.849486e-19, 5.849171e-19, 5.849041e-19 ;

 MEG_acetone =
  1.22078e-16, 1.220548e-16, 1.220592e-16, 1.220408e-16, 1.220508e-16, 
    1.220389e-16, 1.220731e-16, 1.220541e-16, 1.220661e-16, 1.220757e-16, 
    1.220056e-16, 1.220399e-16, 1.219683e-16, 1.219904e-16, 1.219344e-16, 
    1.21972e-16, 1.219267e-16, 1.21935e-16, 1.21909e-16, 1.219164e-16, 
    1.218842e-16, 1.219056e-16, 1.218668e-16, 1.218891e-16, 1.218857e-16, 
    1.219064e-16, 1.220326e-16, 1.2201e-16, 1.22034e-16, 1.220308e-16, 
    1.220321e-16, 1.220508e-16, 1.220605e-16, 1.220795e-16, 1.22076e-16, 
    1.220618e-16, 1.220293e-16, 1.220401e-16, 1.220121e-16, 1.220128e-16, 
    1.21982e-16, 1.219959e-16, 1.21944e-16, 1.219587e-16, 1.219161e-16, 
    1.219269e-16, 1.219167e-16, 1.219197e-16, 1.219167e-16, 1.219324e-16, 
    1.219257e-16, 1.219394e-16, 1.219934e-16, 1.219776e-16, 1.220249e-16, 
    1.22054e-16, 1.220724e-16, 1.220857e-16, 1.220838e-16, 1.220803e-16, 
    1.220618e-16, 1.22044e-16, 1.220306e-16, 1.220217e-16, 1.220129e-16, 
    1.219873e-16, 1.219729e-16, 1.219413e-16, 1.219466e-16, 1.219373e-16, 
    1.219279e-16, 1.219126e-16, 1.219151e-16, 1.219085e-16, 1.219373e-16, 
    1.219183e-16, 1.219498e-16, 1.219412e-16, 1.220119e-16, 1.220371e-16, 
    1.220491e-16, 1.220584e-16, 1.220824e-16, 1.220659e-16, 1.220725e-16, 
    1.220566e-16, 1.220468e-16, 1.220516e-16, 1.220214e-16, 1.220332e-16, 
    1.21972e-16, 1.219983e-16, 1.21929e-16, 1.219455e-16, 1.21925e-16, 
    1.219354e-16, 1.219177e-16, 1.219336e-16, 1.219059e-16, 1.219e-16, 
    1.219041e-16, 1.218881e-16, 1.219345e-16, 1.219168e-16, 1.220518e-16, 
    1.22051e-16, 1.220472e-16, 1.220639e-16, 1.220648e-16, 1.220797e-16, 
    1.220663e-16, 1.220608e-16, 1.220461e-16, 1.220377e-16, 1.220296e-16, 
    1.220119e-16, 1.219923e-16, 1.219646e-16, 1.219444e-16, 1.21931e-16, 
    1.219392e-16, 1.21932e-16, 1.219401e-16, 1.219438e-16, 1.219023e-16, 
    1.219257e-16, 1.218904e-16, 1.218923e-16, 1.219084e-16, 1.218921e-16, 
    1.220504e-16, 1.22055e-16, 1.220711e-16, 1.220585e-16, 1.220813e-16, 
    1.220687e-16, 1.220616e-16, 1.220333e-16, 1.220267e-16, 1.220211e-16, 
    1.220097e-16, 1.219952e-16, 1.219699e-16, 1.219477e-16, 1.219273e-16, 
    1.219288e-16, 1.219283e-16, 1.219239e-16, 1.21935e-16, 1.21922e-16, 
    1.2192e-16, 1.219255e-16, 1.218925e-16, 1.219019e-16, 1.218923e-16, 
    1.218984e-16, 1.220535e-16, 1.220458e-16, 1.2205e-16, 1.220422e-16, 
    1.220478e-16, 1.220235e-16, 1.220162e-16, 1.219818e-16, 1.219956e-16, 
    1.219733e-16, 1.219932e-16, 1.219897e-16, 1.219732e-16, 1.21992e-16, 
    1.219492e-16, 1.219788e-16, 1.219237e-16, 1.219537e-16, 1.219218e-16, 
    1.219274e-16, 1.219181e-16, 1.219099e-16, 1.218993e-16, 1.218803e-16, 
    1.218846e-16, 1.218685e-16, 1.220343e-16, 1.220245e-16, 1.220251e-16, 
    1.220147e-16, 1.22007e-16, 1.219902e-16, 1.219635e-16, 1.219734e-16, 
    1.219549e-16, 1.219512e-16, 1.219793e-16, 1.219623e-16, 1.220178e-16, 
    1.220091e-16, 1.22014e-16, 1.220337e-16, 1.219715e-16, 1.220035e-16, 
    1.219442e-16, 1.219614e-16, 1.219111e-16, 1.219363e-16, 1.218871e-16, 
    1.218668e-16, 1.218464e-16, 1.218242e-16, 1.220189e-16, 1.220255e-16, 
    1.220134e-16, 1.21997e-16, 1.219811e-16, 1.219604e-16, 1.219582e-16, 
    1.219544e-16, 1.219442e-16, 1.219358e-16, 1.219534e-16, 1.219337e-16, 
    1.220076e-16, 1.219686e-16, 1.220283e-16, 1.220107e-16, 1.219979e-16, 
    1.220032e-16, 1.219745e-16, 1.219678e-16, 1.219408e-16, 1.219546e-16, 
    1.21872e-16, 1.219085e-16, 1.218064e-16, 1.21835e-16, 1.220279e-16, 
    1.220188e-16, 1.219873e-16, 1.220022e-16, 1.219589e-16, 1.219484e-16, 
    1.219396e-16, 1.219288e-16, 1.219274e-16, 1.21921e-16, 1.219316e-16, 
    1.219214e-16, 1.219604e-16, 1.219429e-16, 1.219906e-16, 1.219791e-16, 
    1.219843e-16, 1.219902e-16, 1.21972e-16, 1.219532e-16, 1.219524e-16, 
    1.219464e-16, 1.219304e-16, 1.219587e-16, 1.218681e-16, 1.219247e-16, 
    1.220088e-16, 1.219918e-16, 1.219888e-16, 1.219955e-16, 1.219495e-16, 
    1.219662e-16, 1.219211e-16, 1.219332e-16, 1.219133e-16, 1.219232e-16, 
    1.219247e-16, 1.219373e-16, 1.219453e-16, 1.219655e-16, 1.219818e-16, 
    1.219945e-16, 1.219915e-16, 1.219775e-16, 1.21952e-16, 1.219275e-16, 
    1.219329e-16, 1.219148e-16, 1.21962e-16, 1.219424e-16, 1.219502e-16, 
    1.2193e-16, 1.219738e-16, 1.219378e-16, 1.219831e-16, 1.219791e-16, 
    1.219665e-16, 1.219414e-16, 1.219352e-16, 1.219294e-16, 1.219329e-16, 
    1.219512e-16, 1.219541e-16, 1.219667e-16, 1.219704e-16, 1.219799e-16, 
    1.21988e-16, 1.219807e-16, 1.219732e-16, 1.219511e-16, 1.219314e-16, 
    1.219098e-16, 1.219044e-16, 1.218804e-16, 1.219005e-16, 1.218679e-16, 
    1.218965e-16, 1.218465e-16, 1.219351e-16, 1.218965e-16, 1.219658e-16, 
    1.219582e-16, 1.219449e-16, 1.219137e-16, 1.219301e-16, 1.219107e-16, 
    1.219541e-16, 1.219773e-16, 1.219827e-16, 1.219938e-16, 1.219824e-16, 
    1.219833e-16, 1.219726e-16, 1.21976e-16, 1.219503e-16, 1.219641e-16, 
    1.219249e-16, 1.219107e-16, 1.218703e-16, 1.218459e-16, 1.218204e-16, 
    1.218094e-16, 1.21806e-16, 1.218046e-16 ;

 MEG_carene_3 =
  4.842077e-17, 4.84111e-17, 4.841293e-17, 4.840524e-17, 4.840944e-17, 
    4.840446e-17, 4.841873e-17, 4.841079e-17, 4.841581e-17, 4.841979e-17, 
    4.839058e-17, 4.840488e-17, 4.8375e-17, 4.838422e-17, 4.836087e-17, 
    4.837654e-17, 4.835768e-17, 4.836113e-17, 4.83503e-17, 4.835339e-17, 
    4.833994e-17, 4.834887e-17, 4.833269e-17, 4.834197e-17, 4.834059e-17, 
    4.83492e-17, 4.840182e-17, 4.839242e-17, 4.840242e-17, 4.840107e-17, 
    4.840164e-17, 4.840942e-17, 4.841346e-17, 4.842139e-17, 4.841991e-17, 
    4.841402e-17, 4.840046e-17, 4.840494e-17, 4.83933e-17, 4.839356e-17, 
    4.838075e-17, 4.838652e-17, 4.83649e-17, 4.8371e-17, 4.835326e-17, 
    4.835774e-17, 4.83535e-17, 4.835476e-17, 4.835348e-17, 4.836004e-17, 
    4.835724e-17, 4.836296e-17, 4.838548e-17, 4.837891e-17, 4.839862e-17, 
    4.841077e-17, 4.841841e-17, 4.842398e-17, 4.842319e-17, 4.842173e-17, 
    4.841399e-17, 4.840658e-17, 4.840098e-17, 4.839728e-17, 4.83936e-17, 
    4.838295e-17, 4.837692e-17, 4.836376e-17, 4.836598e-17, 4.83621e-17, 
    4.835818e-17, 4.835181e-17, 4.835283e-17, 4.835007e-17, 4.836208e-17, 
    4.835415e-17, 4.836729e-17, 4.83637e-17, 4.839322e-17, 4.84037e-17, 
    4.84087e-17, 4.84126e-17, 4.84226e-17, 4.841573e-17, 4.841845e-17, 
    4.841185e-17, 4.840774e-17, 4.840975e-17, 4.839717e-17, 4.840208e-17, 
    4.837657e-17, 4.838754e-17, 4.835863e-17, 4.836551e-17, 4.835697e-17, 
    4.836129e-17, 4.835393e-17, 4.836055e-17, 4.834899e-17, 4.834654e-17, 
    4.834823e-17, 4.834156e-17, 4.836094e-17, 4.835356e-17, 4.840983e-17, 
    4.840951e-17, 4.840794e-17, 4.841488e-17, 4.841527e-17, 4.842146e-17, 
    4.84159e-17, 4.841358e-17, 4.840746e-17, 4.840396e-17, 4.840059e-17, 
    4.839319e-17, 4.838503e-17, 4.837347e-17, 4.836507e-17, 4.835948e-17, 
    4.836286e-17, 4.835988e-17, 4.836324e-17, 4.836479e-17, 4.83475e-17, 
    4.835725e-17, 4.834252e-17, 4.834331e-17, 4.835002e-17, 4.834322e-17, 
    4.840927e-17, 4.841115e-17, 4.841788e-17, 4.841261e-17, 4.842212e-17, 
    4.841688e-17, 4.841391e-17, 4.840212e-17, 4.839938e-17, 4.839704e-17, 
    4.839227e-17, 4.838623e-17, 4.837569e-17, 4.836644e-17, 4.835792e-17, 
    4.835853e-17, 4.835833e-17, 4.835649e-17, 4.836112e-17, 4.835572e-17, 
    4.835487e-17, 4.835718e-17, 4.834342e-17, 4.834734e-17, 4.834333e-17, 
    4.834586e-17, 4.841052e-17, 4.840734e-17, 4.840907e-17, 4.840585e-17, 
    4.840816e-17, 4.839803e-17, 4.8395e-17, 4.838066e-17, 4.838638e-17, 
    4.83771e-17, 4.838539e-17, 4.838396e-17, 4.837706e-17, 4.83849e-17, 
    4.836706e-17, 4.837939e-17, 4.835642e-17, 4.836894e-17, 4.835565e-17, 
    4.835796e-17, 4.835407e-17, 4.835065e-17, 4.834625e-17, 4.83383e-17, 
    4.834012e-17, 4.833338e-17, 4.840253e-17, 4.839846e-17, 4.83987e-17, 
    4.839436e-17, 4.839118e-17, 4.838414e-17, 4.8373e-17, 4.837715e-17, 
    4.836941e-17, 4.83679e-17, 4.837959e-17, 4.837252e-17, 4.839564e-17, 
    4.839202e-17, 4.839409e-17, 4.840227e-17, 4.837635e-17, 4.838971e-17, 
    4.836495e-17, 4.837215e-17, 4.835116e-17, 4.83617e-17, 4.834114e-17, 
    4.833268e-17, 4.83242e-17, 4.831492e-17, 4.839611e-17, 4.839889e-17, 
    4.839381e-17, 4.8387e-17, 4.838036e-17, 4.837174e-17, 4.837079e-17, 
    4.836921e-17, 4.836497e-17, 4.836147e-17, 4.836882e-17, 4.836058e-17, 
    4.839141e-17, 4.837514e-17, 4.840004e-17, 4.839269e-17, 4.838735e-17, 
    4.838958e-17, 4.83776e-17, 4.837482e-17, 4.836357e-17, 4.836932e-17, 
    4.833487e-17, 4.835009e-17, 4.830749e-17, 4.831943e-17, 4.839989e-17, 
    4.839606e-17, 4.838294e-17, 4.838916e-17, 4.83711e-17, 4.83667e-17, 
    4.836304e-17, 4.835855e-17, 4.835798e-17, 4.835531e-17, 4.83597e-17, 
    4.835544e-17, 4.837172e-17, 4.836441e-17, 4.83843e-17, 4.837952e-17, 
    4.838168e-17, 4.838414e-17, 4.837658e-17, 4.836873e-17, 4.836838e-17, 
    4.836589e-17, 4.835924e-17, 4.837102e-17, 4.833325e-17, 4.835685e-17, 
    4.839191e-17, 4.838481e-17, 4.838357e-17, 4.838636e-17, 4.836716e-17, 
    4.837413e-17, 4.835535e-17, 4.836038e-17, 4.835209e-17, 4.835622e-17, 
    4.835684e-17, 4.836211e-17, 4.836544e-17, 4.837384e-17, 4.838064e-17, 
    4.838593e-17, 4.838468e-17, 4.837887e-17, 4.836821e-17, 4.835801e-17, 
    4.836027e-17, 4.835272e-17, 4.837241e-17, 4.836423e-17, 4.836746e-17, 
    4.835904e-17, 4.83773e-17, 4.836231e-17, 4.838121e-17, 4.837951e-17, 
    4.837427e-17, 4.836381e-17, 4.836122e-17, 4.83588e-17, 4.836026e-17, 
    4.83679e-17, 4.836908e-17, 4.837435e-17, 4.83759e-17, 4.837986e-17, 
    4.838324e-17, 4.83802e-17, 4.837705e-17, 4.836783e-17, 4.835962e-17, 
    4.835063e-17, 4.834836e-17, 4.833835e-17, 4.834675e-17, 4.833315e-17, 
    4.834509e-17, 4.832424e-17, 4.836116e-17, 4.834508e-17, 4.837397e-17, 
    4.83708e-17, 4.836527e-17, 4.835224e-17, 4.835907e-17, 4.835099e-17, 
    4.836911e-17, 4.837876e-17, 4.838103e-17, 4.838564e-17, 4.838092e-17, 
    4.838129e-17, 4.837679e-17, 4.837823e-17, 4.836752e-17, 4.837326e-17, 
    4.835691e-17, 4.835101e-17, 4.833416e-17, 4.832397e-17, 4.831333e-17, 
    4.830874e-17, 4.830733e-17, 4.830675e-17 ;

 MEG_ethanol =
  3.91629e-18, 3.914856e-18, 3.915128e-18, 3.913988e-18, 3.91461e-18, 
    3.913871e-18, 3.915987e-18, 3.91481e-18, 3.915554e-18, 3.916144e-18, 
    3.911814e-18, 3.913934e-18, 3.909504e-18, 3.91087e-18, 3.907406e-18, 
    3.909732e-18, 3.906933e-18, 3.907446e-18, 3.905837e-18, 3.906296e-18, 
    3.904299e-18, 3.905625e-18, 3.903221e-18, 3.904601e-18, 3.904395e-18, 
    3.905673e-18, 3.913481e-18, 3.912086e-18, 3.91357e-18, 3.913369e-18, 
    3.913454e-18, 3.914607e-18, 3.915207e-18, 3.91638e-18, 3.916163e-18, 
    3.91529e-18, 3.913279e-18, 3.913943e-18, 3.912217e-18, 3.912255e-18, 
    3.910355e-18, 3.911212e-18, 3.908005e-18, 3.908909e-18, 3.906277e-18, 
    3.906942e-18, 3.906312e-18, 3.9065e-18, 3.90631e-18, 3.907284e-18, 
    3.906868e-18, 3.907717e-18, 3.911057e-18, 3.910083e-18, 3.913005e-18, 
    3.914808e-18, 3.91594e-18, 3.916765e-18, 3.916649e-18, 3.916431e-18, 
    3.915285e-18, 3.914186e-18, 3.913356e-18, 3.912806e-18, 3.912261e-18, 
    3.910682e-18, 3.909789e-18, 3.907836e-18, 3.908165e-18, 3.907589e-18, 
    3.907007e-18, 3.906062e-18, 3.906214e-18, 3.905803e-18, 3.907588e-18, 
    3.906409e-18, 3.908358e-18, 3.907827e-18, 3.912205e-18, 3.913759e-18, 
    3.9145e-18, 3.915079e-18, 3.91656e-18, 3.915543e-18, 3.915946e-18, 
    3.914967e-18, 3.914359e-18, 3.914655e-18, 3.912791e-18, 3.913519e-18, 
    3.909736e-18, 3.911363e-18, 3.907075e-18, 3.908095e-18, 3.906827e-18, 
    3.907469e-18, 3.906377e-18, 3.90736e-18, 3.905642e-18, 3.905279e-18, 
    3.90553e-18, 3.904539e-18, 3.907417e-18, 3.906321e-18, 3.914668e-18, 
    3.914621e-18, 3.914387e-18, 3.915416e-18, 3.915475e-18, 3.916391e-18, 
    3.915567e-18, 3.915224e-18, 3.914316e-18, 3.913797e-18, 3.913298e-18, 
    3.9122e-18, 3.91099e-18, 3.909275e-18, 3.90803e-18, 3.907201e-18, 
    3.907703e-18, 3.90726e-18, 3.907759e-18, 3.907988e-18, 3.905422e-18, 
    3.90687e-18, 3.904681e-18, 3.904799e-18, 3.905796e-18, 3.904786e-18, 
    3.914586e-18, 3.914864e-18, 3.915861e-18, 3.91508e-18, 3.91649e-18, 
    3.915713e-18, 3.915272e-18, 3.913524e-18, 3.913118e-18, 3.912771e-18, 
    3.912064e-18, 3.911169e-18, 3.909606e-18, 3.908234e-18, 3.906969e-18, 
    3.90706e-18, 3.907029e-18, 3.906756e-18, 3.907444e-18, 3.906643e-18, 
    3.906517e-18, 3.906859e-18, 3.904815e-18, 3.905398e-18, 3.904802e-18, 
    3.905178e-18, 3.914771e-18, 3.914298e-18, 3.914555e-18, 3.914077e-18, 
    3.914421e-18, 3.912919e-18, 3.912469e-18, 3.910342e-18, 3.911191e-18, 
    3.909814e-18, 3.911044e-18, 3.910831e-18, 3.909808e-18, 3.910972e-18, 
    3.908327e-18, 3.910153e-18, 3.906746e-18, 3.908603e-18, 3.906631e-18, 
    3.906975e-18, 3.906397e-18, 3.90589e-18, 3.905235e-18, 3.904056e-18, 
    3.904325e-18, 3.903324e-18, 3.913585e-18, 3.912982e-18, 3.913018e-18, 
    3.912374e-18, 3.911902e-18, 3.910858e-18, 3.909207e-18, 3.909822e-18, 
    3.908674e-18, 3.90845e-18, 3.910183e-18, 3.909135e-18, 3.912564e-18, 
    3.912027e-18, 3.912334e-18, 3.913547e-18, 3.909704e-18, 3.911685e-18, 
    3.908013e-18, 3.90908e-18, 3.905965e-18, 3.90753e-18, 3.904477e-18, 
    3.903219e-18, 3.901958e-18, 3.900578e-18, 3.912633e-18, 3.913045e-18, 
    3.912292e-18, 3.911283e-18, 3.910298e-18, 3.909019e-18, 3.908878e-18, 
    3.908644e-18, 3.908015e-18, 3.907495e-18, 3.908586e-18, 3.907364e-18, 
    3.911937e-18, 3.909524e-18, 3.913217e-18, 3.912127e-18, 3.911335e-18, 
    3.911665e-18, 3.909888e-18, 3.909476e-18, 3.907808e-18, 3.90866e-18, 
    3.903545e-18, 3.905807e-18, 3.899472e-18, 3.901249e-18, 3.913193e-18, 
    3.912626e-18, 3.910681e-18, 3.911604e-18, 3.908924e-18, 3.908273e-18, 
    3.907729e-18, 3.907063e-18, 3.906978e-18, 3.906582e-18, 3.907234e-18, 
    3.906601e-18, 3.909016e-18, 3.907933e-18, 3.910882e-18, 3.910174e-18, 
    3.910494e-18, 3.910858e-18, 3.909737e-18, 3.908574e-18, 3.908521e-18, 
    3.908152e-18, 3.907165e-18, 3.908912e-18, 3.903304e-18, 3.906811e-18, 
    3.91201e-18, 3.910958e-18, 3.910774e-18, 3.911187e-18, 3.908339e-18, 
    3.909374e-18, 3.906588e-18, 3.907334e-18, 3.906104e-18, 3.906717e-18, 
    3.906809e-18, 3.90759e-18, 3.908086e-18, 3.909332e-18, 3.910339e-18, 
    3.911124e-18, 3.910939e-18, 3.910076e-18, 3.908496e-18, 3.906983e-18, 
    3.907318e-18, 3.906197e-18, 3.909119e-18, 3.907907e-18, 3.908384e-18, 
    3.907135e-18, 3.909844e-18, 3.907621e-18, 3.910423e-18, 3.910171e-18, 
    3.909394e-18, 3.907844e-18, 3.907459e-18, 3.9071e-18, 3.907316e-18, 
    3.90845e-18, 3.908624e-18, 3.909406e-18, 3.909636e-18, 3.910224e-18, 
    3.910724e-18, 3.910274e-18, 3.909807e-18, 3.908439e-18, 3.907221e-18, 
    3.905887e-18, 3.90555e-18, 3.904063e-18, 3.905311e-18, 3.90329e-18, 
    3.905064e-18, 3.901965e-18, 3.907451e-18, 3.905062e-18, 3.909349e-18, 
    3.90888e-18, 3.90806e-18, 3.906126e-18, 3.90714e-18, 3.90594e-18, 
    3.908629e-18, 3.91006e-18, 3.910397e-18, 3.911081e-18, 3.910381e-18, 
    3.910436e-18, 3.909769e-18, 3.909981e-18, 3.908393e-18, 3.909245e-18, 
    3.906818e-18, 3.905942e-18, 3.903438e-18, 3.901924e-18, 3.900341e-18, 
    3.899658e-18, 3.899447e-18, 3.899361e-18 ;

 MEG_formaldehyde =
  7.832579e-19, 7.829712e-19, 7.830256e-19, 7.827976e-19, 7.82922e-19, 
    7.827742e-19, 7.831973e-19, 7.82962e-19, 7.831108e-19, 7.832288e-19, 
    7.823628e-19, 7.827867e-19, 7.819007e-19, 7.82174e-19, 7.814813e-19, 
    7.819463e-19, 7.813867e-19, 7.814892e-19, 7.811675e-19, 7.812592e-19, 
    7.808597e-19, 7.81125e-19, 7.806442e-19, 7.809201e-19, 7.80879e-19, 
    7.811347e-19, 7.826961e-19, 7.824173e-19, 7.827139e-19, 7.826738e-19, 
    7.826907e-19, 7.829213e-19, 7.830413e-19, 7.832761e-19, 7.832325e-19, 
    7.830579e-19, 7.826557e-19, 7.827885e-19, 7.824433e-19, 7.82451e-19, 
    7.820711e-19, 7.822423e-19, 7.81601e-19, 7.817818e-19, 7.812553e-19, 
    7.813884e-19, 7.812625e-19, 7.812999e-19, 7.81262e-19, 7.814568e-19, 
    7.813737e-19, 7.815435e-19, 7.822113e-19, 7.820166e-19, 7.826011e-19, 
    7.829616e-19, 7.83188e-19, 7.833529e-19, 7.833296e-19, 7.832863e-19, 
    7.83057e-19, 7.828371e-19, 7.826712e-19, 7.825612e-19, 7.824521e-19, 
    7.821365e-19, 7.819577e-19, 7.815671e-19, 7.816329e-19, 7.815178e-19, 
    7.814013e-19, 7.812123e-19, 7.812427e-19, 7.811606e-19, 7.815175e-19, 
    7.812819e-19, 7.816716e-19, 7.815654e-19, 7.824409e-19, 7.827518e-19, 
    7.829e-19, 7.830158e-19, 7.83312e-19, 7.831085e-19, 7.831891e-19, 
    7.829934e-19, 7.828717e-19, 7.829311e-19, 7.825582e-19, 7.827038e-19, 
    7.819472e-19, 7.822725e-19, 7.81415e-19, 7.81619e-19, 7.813655e-19, 
    7.814938e-19, 7.812753e-19, 7.814719e-19, 7.811285e-19, 7.810559e-19, 
    7.811059e-19, 7.809078e-19, 7.814833e-19, 7.812642e-19, 7.829336e-19, 
    7.829241e-19, 7.828774e-19, 7.830833e-19, 7.830949e-19, 7.832782e-19, 
    7.831133e-19, 7.830447e-19, 7.828632e-19, 7.827594e-19, 7.826595e-19, 
    7.824399e-19, 7.82198e-19, 7.81855e-19, 7.81606e-19, 7.814402e-19, 
    7.815406e-19, 7.814521e-19, 7.815517e-19, 7.815977e-19, 7.810843e-19, 
    7.813739e-19, 7.809363e-19, 7.809598e-19, 7.811592e-19, 7.809571e-19, 
    7.82917e-19, 7.829727e-19, 7.831722e-19, 7.83016e-19, 7.83298e-19, 
    7.831424e-19, 7.830544e-19, 7.827048e-19, 7.826236e-19, 7.825542e-19, 
    7.824128e-19, 7.822337e-19, 7.819211e-19, 7.816467e-19, 7.813938e-19, 
    7.81412e-19, 7.814058e-19, 7.813512e-19, 7.814889e-19, 7.813285e-19, 
    7.813033e-19, 7.813718e-19, 7.809631e-19, 7.810795e-19, 7.809603e-19, 
    7.810356e-19, 7.829541e-19, 7.828596e-19, 7.82911e-19, 7.828154e-19, 
    7.828842e-19, 7.825838e-19, 7.824938e-19, 7.820684e-19, 7.822382e-19, 
    7.819629e-19, 7.822088e-19, 7.821663e-19, 7.819616e-19, 7.821943e-19, 
    7.816653e-19, 7.820307e-19, 7.813491e-19, 7.817207e-19, 7.813263e-19, 
    7.81395e-19, 7.812794e-19, 7.811779e-19, 7.81047e-19, 7.80811e-19, 
    7.808649e-19, 7.806648e-19, 7.82717e-19, 7.825963e-19, 7.826035e-19, 
    7.824747e-19, 7.823803e-19, 7.821716e-19, 7.818413e-19, 7.819643e-19, 
    7.817348e-19, 7.8169e-19, 7.820367e-19, 7.81827e-19, 7.825128e-19, 
    7.824055e-19, 7.824668e-19, 7.827095e-19, 7.819408e-19, 7.823369e-19, 
    7.816025e-19, 7.81816e-19, 7.811929e-19, 7.81506e-19, 7.808954e-19, 
    7.806438e-19, 7.803915e-19, 7.801155e-19, 7.825267e-19, 7.82609e-19, 
    7.824584e-19, 7.822566e-19, 7.820597e-19, 7.818037e-19, 7.817756e-19, 
    7.817287e-19, 7.81603e-19, 7.81499e-19, 7.817172e-19, 7.814727e-19, 
    7.823874e-19, 7.819048e-19, 7.826433e-19, 7.824254e-19, 7.822669e-19, 
    7.823329e-19, 7.819775e-19, 7.818951e-19, 7.815616e-19, 7.817319e-19, 
    7.807089e-19, 7.811613e-19, 7.798944e-19, 7.802498e-19, 7.826386e-19, 
    7.825253e-19, 7.821362e-19, 7.823206e-19, 7.817847e-19, 7.816546e-19, 
    7.815458e-19, 7.814126e-19, 7.813956e-19, 7.813163e-19, 7.814467e-19, 
    7.813202e-19, 7.818031e-19, 7.815866e-19, 7.821765e-19, 7.820348e-19, 
    7.820988e-19, 7.821715e-19, 7.819474e-19, 7.817147e-19, 7.817041e-19, 
    7.816304e-19, 7.814329e-19, 7.817824e-19, 7.806608e-19, 7.813621e-19, 
    7.82402e-19, 7.821916e-19, 7.821547e-19, 7.822374e-19, 7.816679e-19, 
    7.818747e-19, 7.813175e-19, 7.814667e-19, 7.812208e-19, 7.813434e-19, 
    7.813617e-19, 7.815181e-19, 7.816171e-19, 7.818663e-19, 7.820677e-19, 
    7.822247e-19, 7.821878e-19, 7.820152e-19, 7.816991e-19, 7.813966e-19, 
    7.814635e-19, 7.812394e-19, 7.818237e-19, 7.815813e-19, 7.816768e-19, 
    7.81427e-19, 7.819688e-19, 7.815241e-19, 7.820846e-19, 7.820342e-19, 
    7.818788e-19, 7.815687e-19, 7.814918e-19, 7.814199e-19, 7.814632e-19, 
    7.8169e-19, 7.817248e-19, 7.818812e-19, 7.819272e-19, 7.820448e-19, 
    7.821449e-19, 7.820548e-19, 7.819614e-19, 7.816877e-19, 7.814442e-19, 
    7.811774e-19, 7.811099e-19, 7.808124e-19, 7.810621e-19, 7.806579e-19, 
    7.810129e-19, 7.80393e-19, 7.814901e-19, 7.810124e-19, 7.818698e-19, 
    7.817759e-19, 7.816121e-19, 7.812251e-19, 7.814281e-19, 7.81188e-19, 
    7.817257e-19, 7.82012e-19, 7.820793e-19, 7.822162e-19, 7.820762e-19, 
    7.820873e-19, 7.819537e-19, 7.819963e-19, 7.816785e-19, 7.818489e-19, 
    7.813636e-19, 7.811884e-19, 7.806877e-19, 7.803848e-19, 7.800682e-19, 
    7.799315e-19, 7.798895e-19, 7.798721e-19 ;

 MEG_isoprene =
  6.252617e-19, 6.249928e-19, 6.250438e-19, 6.248299e-19, 6.249466e-19, 
    6.24808e-19, 6.252049e-19, 6.249842e-19, 6.251238e-19, 6.252344e-19, 
    6.24422e-19, 6.248197e-19, 6.239885e-19, 6.242448e-19, 6.235949e-19, 
    6.240313e-19, 6.23506e-19, 6.236023e-19, 6.233003e-19, 6.233865e-19, 
    6.230115e-19, 6.232605e-19, 6.228092e-19, 6.230682e-19, 6.230296e-19, 
    6.232696e-19, 6.247347e-19, 6.244731e-19, 6.247514e-19, 6.247138e-19, 
    6.247296e-19, 6.24946e-19, 6.250586e-19, 6.252789e-19, 6.252379e-19, 
    6.250742e-19, 6.246968e-19, 6.248214e-19, 6.244975e-19, 6.245047e-19, 
    6.241483e-19, 6.24309e-19, 6.237072e-19, 6.238769e-19, 6.233828e-19, 
    6.235077e-19, 6.233895e-19, 6.234247e-19, 6.233891e-19, 6.235719e-19, 
    6.234938e-19, 6.236532e-19, 6.242799e-19, 6.240971e-19, 6.246455e-19, 
    6.249838e-19, 6.251962e-19, 6.253509e-19, 6.253291e-19, 6.252884e-19, 
    6.250733e-19, 6.24867e-19, 6.247114e-19, 6.246082e-19, 6.245058e-19, 
    6.242097e-19, 6.240419e-19, 6.236754e-19, 6.237371e-19, 6.236291e-19, 
    6.235199e-19, 6.233424e-19, 6.23371e-19, 6.232939e-19, 6.236288e-19, 
    6.234077e-19, 6.237734e-19, 6.236739e-19, 6.244953e-19, 6.247869e-19, 
    6.24926e-19, 6.250346e-19, 6.253126e-19, 6.251216e-19, 6.251973e-19, 
    6.250136e-19, 6.248995e-19, 6.249552e-19, 6.246053e-19, 6.247419e-19, 
    6.240321e-19, 6.243373e-19, 6.235326e-19, 6.237241e-19, 6.234861e-19, 
    6.236067e-19, 6.234016e-19, 6.235861e-19, 6.232638e-19, 6.231956e-19, 
    6.232425e-19, 6.230566e-19, 6.235968e-19, 6.233912e-19, 6.249575e-19, 
    6.249486e-19, 6.249048e-19, 6.25098e-19, 6.251088e-19, 6.252808e-19, 
    6.251262e-19, 6.250618e-19, 6.248915e-19, 6.247941e-19, 6.247003e-19, 
    6.244944e-19, 6.242674e-19, 6.239455e-19, 6.237119e-19, 6.235563e-19, 
    6.236505e-19, 6.235675e-19, 6.23661e-19, 6.237041e-19, 6.232223e-19, 
    6.234941e-19, 6.230833e-19, 6.231054e-19, 6.232926e-19, 6.231029e-19, 
    6.24942e-19, 6.249943e-19, 6.251813e-19, 6.250349e-19, 6.252994e-19, 
    6.251535e-19, 6.250708e-19, 6.247429e-19, 6.246667e-19, 6.246015e-19, 
    6.244688e-19, 6.243009e-19, 6.240076e-19, 6.237501e-19, 6.235128e-19, 
    6.235299e-19, 6.23524e-19, 6.234728e-19, 6.23602e-19, 6.234515e-19, 
    6.234278e-19, 6.234921e-19, 6.231085e-19, 6.232178e-19, 6.23106e-19, 
    6.231766e-19, 6.249768e-19, 6.248881e-19, 6.249363e-19, 6.248467e-19, 
    6.249111e-19, 6.246294e-19, 6.245449e-19, 6.241457e-19, 6.243051e-19, 
    6.240468e-19, 6.242775e-19, 6.242376e-19, 6.240456e-19, 6.242639e-19, 
    6.237675e-19, 6.241104e-19, 6.234708e-19, 6.238195e-19, 6.234494e-19, 
    6.235139e-19, 6.234054e-19, 6.233102e-19, 6.231873e-19, 6.229658e-19, 
    6.230164e-19, 6.228285e-19, 6.247543e-19, 6.24641e-19, 6.246478e-19, 
    6.24527e-19, 6.244384e-19, 6.242426e-19, 6.239327e-19, 6.240481e-19, 
    6.238327e-19, 6.237907e-19, 6.24116e-19, 6.239193e-19, 6.245627e-19, 
    6.24462e-19, 6.245196e-19, 6.247473e-19, 6.24026e-19, 6.243978e-19, 
    6.237087e-19, 6.239089e-19, 6.233242e-19, 6.236181e-19, 6.230449e-19, 
    6.228089e-19, 6.22572e-19, 6.223129e-19, 6.245757e-19, 6.24653e-19, 
    6.245116e-19, 6.243223e-19, 6.241376e-19, 6.238974e-19, 6.23871e-19, 
    6.23827e-19, 6.23709e-19, 6.236116e-19, 6.238162e-19, 6.235868e-19, 
    6.244451e-19, 6.239923e-19, 6.246852e-19, 6.244807e-19, 6.24332e-19, 
    6.243939e-19, 6.240605e-19, 6.239832e-19, 6.236702e-19, 6.238301e-19, 
    6.228699e-19, 6.232946e-19, 6.221053e-19, 6.22439e-19, 6.246808e-19, 
    6.245744e-19, 6.242094e-19, 6.243824e-19, 6.238796e-19, 6.237575e-19, 
    6.236554e-19, 6.235304e-19, 6.235145e-19, 6.2344e-19, 6.235625e-19, 
    6.234436e-19, 6.238968e-19, 6.236937e-19, 6.242472e-19, 6.241142e-19, 
    6.241743e-19, 6.242425e-19, 6.240322e-19, 6.238139e-19, 6.238039e-19, 
    6.237348e-19, 6.235495e-19, 6.238774e-19, 6.228248e-19, 6.234831e-19, 
    6.244588e-19, 6.242614e-19, 6.242268e-19, 6.243043e-19, 6.2377e-19, 
    6.23964e-19, 6.234411e-19, 6.235812e-19, 6.233504e-19, 6.234655e-19, 
    6.234827e-19, 6.236294e-19, 6.237223e-19, 6.239561e-19, 6.241452e-19, 
    6.242924e-19, 6.242578e-19, 6.240958e-19, 6.237992e-19, 6.235154e-19, 
    6.235782e-19, 6.233679e-19, 6.239162e-19, 6.236888e-19, 6.237783e-19, 
    6.235439e-19, 6.240523e-19, 6.23635e-19, 6.24161e-19, 6.241137e-19, 
    6.239678e-19, 6.236769e-19, 6.236047e-19, 6.235373e-19, 6.235779e-19, 
    6.237908e-19, 6.238234e-19, 6.239701e-19, 6.240133e-19, 6.241236e-19, 
    6.242175e-19, 6.241331e-19, 6.240454e-19, 6.237886e-19, 6.235601e-19, 
    6.233097e-19, 6.232463e-19, 6.229671e-19, 6.232015e-19, 6.228221e-19, 
    6.231553e-19, 6.225735e-19, 6.236031e-19, 6.231548e-19, 6.239594e-19, 
    6.238714e-19, 6.237175e-19, 6.233544e-19, 6.235449e-19, 6.233196e-19, 
    6.238243e-19, 6.240928e-19, 6.24156e-19, 6.242844e-19, 6.24153e-19, 
    6.241635e-19, 6.240381e-19, 6.240781e-19, 6.2378e-19, 6.239398e-19, 
    6.234845e-19, 6.233201e-19, 6.2285e-19, 6.225658e-19, 6.222685e-19, 
    6.221401e-19, 6.221006e-19, 6.220844e-19 ;

 MEG_methanol =
  8.573229e-17, 8.571757e-17, 8.572036e-17, 8.570866e-17, 8.571504e-17, 
    8.570747e-17, 8.572918e-17, 8.57171e-17, 8.572474e-17, 8.573079e-17, 
    8.568635e-17, 8.57081e-17, 8.566265e-17, 8.567667e-17, 8.564113e-17, 
    8.566498e-17, 8.563628e-17, 8.564153e-17, 8.562505e-17, 8.562975e-17, 
    8.560928e-17, 8.562287e-17, 8.559825e-17, 8.561237e-17, 8.561027e-17, 
    8.562336e-17, 8.570346e-17, 8.568914e-17, 8.570437e-17, 8.570231e-17, 
    8.570318e-17, 8.571501e-17, 8.572116e-17, 8.573322e-17, 8.573098e-17, 
    8.572202e-17, 8.570138e-17, 8.57082e-17, 8.569049e-17, 8.569088e-17, 
    8.567139e-17, 8.568018e-17, 8.564726e-17, 8.565654e-17, 8.562955e-17, 
    8.563636e-17, 8.562992e-17, 8.563183e-17, 8.562989e-17, 8.563987e-17, 
    8.563561e-17, 8.564432e-17, 8.567858e-17, 8.566859e-17, 8.569858e-17, 
    8.571707e-17, 8.57287e-17, 8.573716e-17, 8.573597e-17, 8.573374e-17, 
    8.572197e-17, 8.571069e-17, 8.570218e-17, 8.569654e-17, 8.569094e-17, 
    8.567474e-17, 8.566556e-17, 8.564553e-17, 8.56489e-17, 8.5643e-17, 
    8.563703e-17, 8.562734e-17, 8.56289e-17, 8.562469e-17, 8.564298e-17, 
    8.56309e-17, 8.565089e-17, 8.564544e-17, 8.569036e-17, 8.570631e-17, 
    8.571392e-17, 8.571986e-17, 8.573507e-17, 8.572462e-17, 8.572876e-17, 
    8.571872e-17, 8.571247e-17, 8.571551e-17, 8.569638e-17, 8.570385e-17, 
    8.566503e-17, 8.568172e-17, 8.563773e-17, 8.564819e-17, 8.563519e-17, 
    8.564177e-17, 8.563057e-17, 8.564065e-17, 8.562305e-17, 8.561933e-17, 
    8.562189e-17, 8.561174e-17, 8.564123e-17, 8.563e-17, 8.571564e-17, 
    8.571515e-17, 8.571276e-17, 8.572332e-17, 8.572392e-17, 8.573333e-17, 
    8.572487e-17, 8.572134e-17, 8.571203e-17, 8.57067e-17, 8.570158e-17, 
    8.569031e-17, 8.56779e-17, 8.56603e-17, 8.564752e-17, 8.563902e-17, 
    8.564417e-17, 8.563963e-17, 8.564474e-17, 8.564709e-17, 8.562078e-17, 
    8.563562e-17, 8.561321e-17, 8.561441e-17, 8.562462e-17, 8.561427e-17, 
    8.571479e-17, 8.571765e-17, 8.572789e-17, 8.571987e-17, 8.573435e-17, 
    8.572636e-17, 8.572184e-17, 8.57039e-17, 8.569974e-17, 8.569618e-17, 
    8.568892e-17, 8.567973e-17, 8.566369e-17, 8.56496e-17, 8.563665e-17, 
    8.563758e-17, 8.563725e-17, 8.563446e-17, 8.564152e-17, 8.56333e-17, 
    8.563201e-17, 8.563551e-17, 8.561458e-17, 8.562054e-17, 8.561444e-17, 
    8.56183e-17, 8.57167e-17, 8.571185e-17, 8.571448e-17, 8.570958e-17, 
    8.57131e-17, 8.569769e-17, 8.569307e-17, 8.567124e-17, 8.567996e-17, 
    8.566584e-17, 8.567845e-17, 8.567627e-17, 8.566576e-17, 8.567771e-17, 
    8.565056e-17, 8.566931e-17, 8.563436e-17, 8.565341e-17, 8.563318e-17, 
    8.563671e-17, 8.563078e-17, 8.562558e-17, 8.561888e-17, 8.560679e-17, 
    8.560955e-17, 8.559931e-17, 8.570453e-17, 8.569833e-17, 8.56987e-17, 
    8.56921e-17, 8.568726e-17, 8.567654e-17, 8.56596e-17, 8.566591e-17, 
    8.565414e-17, 8.565183e-17, 8.566962e-17, 8.565886e-17, 8.569405e-17, 
    8.568855e-17, 8.56917e-17, 8.570414e-17, 8.56647e-17, 8.568503e-17, 
    8.564734e-17, 8.56583e-17, 8.562635e-17, 8.564239e-17, 8.561111e-17, 
    8.559823e-17, 8.558533e-17, 8.557122e-17, 8.569476e-17, 8.569899e-17, 
    8.569126e-17, 8.56809e-17, 8.56708e-17, 8.565767e-17, 8.565623e-17, 
    8.565382e-17, 8.564737e-17, 8.564204e-17, 8.565323e-17, 8.564069e-17, 
    8.568761e-17, 8.566286e-17, 8.570075e-17, 8.568957e-17, 8.568143e-17, 
    8.568482e-17, 8.566659e-17, 8.566235e-17, 8.564524e-17, 8.565399e-17, 
    8.560156e-17, 8.562473e-17, 8.555992e-17, 8.557808e-17, 8.570051e-17, 
    8.569469e-17, 8.567472e-17, 8.568419e-17, 8.56567e-17, 8.565001e-17, 
    8.564443e-17, 8.563761e-17, 8.563674e-17, 8.563267e-17, 8.563936e-17, 
    8.563287e-17, 8.565764e-17, 8.564653e-17, 8.567679e-17, 8.566952e-17, 
    8.567281e-17, 8.567654e-17, 8.566504e-17, 8.56531e-17, 8.565256e-17, 
    8.564877e-17, 8.563864e-17, 8.565658e-17, 8.559909e-17, 8.563501e-17, 
    8.568837e-17, 8.567757e-17, 8.567568e-17, 8.567992e-17, 8.56507e-17, 
    8.566131e-17, 8.563273e-17, 8.564038e-17, 8.562778e-17, 8.563406e-17, 
    8.5635e-17, 8.564301e-17, 8.564809e-17, 8.566088e-17, 8.567122e-17, 
    8.567927e-17, 8.567738e-17, 8.566852e-17, 8.56523e-17, 8.563678e-17, 
    8.564022e-17, 8.562873e-17, 8.565869e-17, 8.564625e-17, 8.565116e-17, 
    8.563835e-17, 8.566614e-17, 8.564332e-17, 8.567208e-17, 8.566949e-17, 
    8.566152e-17, 8.564561e-17, 8.564167e-17, 8.563798e-17, 8.56402e-17, 
    8.565184e-17, 8.565362e-17, 8.566165e-17, 8.5664e-17, 8.567004e-17, 
    8.567517e-17, 8.567055e-17, 8.566576e-17, 8.565172e-17, 8.563923e-17, 
    8.562555e-17, 8.56221e-17, 8.560686e-17, 8.561965e-17, 8.559895e-17, 
    8.561712e-17, 8.55854e-17, 8.564157e-17, 8.56171e-17, 8.566106e-17, 
    8.565625e-17, 8.564783e-17, 8.5628e-17, 8.56384e-17, 8.56261e-17, 
    8.565367e-17, 8.566835e-17, 8.56718e-17, 8.567883e-17, 8.567165e-17, 
    8.567222e-17, 8.566537e-17, 8.566755e-17, 8.565125e-17, 8.565999e-17, 
    8.56351e-17, 8.562612e-17, 8.560048e-17, 8.558498e-17, 8.55688e-17, 
    8.556182e-17, 8.555967e-17, 8.555878e-17 ;

 MEG_pinene_a =
  7.460867e-17, 7.459253e-17, 7.459559e-17, 7.458275e-17, 7.458975e-17, 
    7.458144e-17, 7.460526e-17, 7.459201e-17, 7.460039e-17, 7.460703e-17, 
    7.455828e-17, 7.458214e-17, 7.453228e-17, 7.454765e-17, 7.450867e-17, 
    7.453484e-17, 7.450335e-17, 7.450911e-17, 7.449103e-17, 7.449619e-17, 
    7.447373e-17, 7.448865e-17, 7.446163e-17, 7.447713e-17, 7.447482e-17, 
    7.448919e-17, 7.457704e-17, 7.456135e-17, 7.457805e-17, 7.457578e-17, 
    7.457674e-17, 7.458972e-17, 7.459647e-17, 7.46097e-17, 7.460724e-17, 
    7.459741e-17, 7.457477e-17, 7.458224e-17, 7.456282e-17, 7.456324e-17, 
    7.454186e-17, 7.455151e-17, 7.451541e-17, 7.452559e-17, 7.449597e-17, 
    7.450345e-17, 7.449637e-17, 7.449848e-17, 7.449634e-17, 7.45073e-17, 
    7.450262e-17, 7.451217e-17, 7.454976e-17, 7.45388e-17, 7.45717e-17, 
    7.459198e-17, 7.460474e-17, 7.461403e-17, 7.461271e-17, 7.461027e-17, 
    7.459736e-17, 7.458498e-17, 7.457565e-17, 7.456945e-17, 7.456331e-17, 
    7.454554e-17, 7.453548e-17, 7.45135e-17, 7.45172e-17, 7.451073e-17, 
    7.450418e-17, 7.449355e-17, 7.449526e-17, 7.449064e-17, 7.451071e-17, 
    7.449746e-17, 7.451938e-17, 7.451341e-17, 7.456268e-17, 7.458018e-17, 
    7.458852e-17, 7.459504e-17, 7.461172e-17, 7.460026e-17, 7.46048e-17, 
    7.459378e-17, 7.458693e-17, 7.459027e-17, 7.456928e-17, 7.457747e-17, 
    7.45349e-17, 7.45532e-17, 7.450495e-17, 7.451642e-17, 7.450216e-17, 
    7.450938e-17, 7.449709e-17, 7.450815e-17, 7.448884e-17, 7.448476e-17, 
    7.448757e-17, 7.447644e-17, 7.450879e-17, 7.449647e-17, 7.459042e-17, 
    7.458987e-17, 7.458725e-17, 7.459884e-17, 7.45995e-17, 7.460982e-17, 
    7.460053e-17, 7.459667e-17, 7.458645e-17, 7.458061e-17, 7.457498e-17, 
    7.456263e-17, 7.4549e-17, 7.452971e-17, 7.451569e-17, 7.450636e-17, 
    7.451201e-17, 7.450703e-17, 7.451263e-17, 7.451522e-17, 7.448636e-17, 
    7.450264e-17, 7.447804e-17, 7.447936e-17, 7.449057e-17, 7.447921e-17, 
    7.458948e-17, 7.459261e-17, 7.460384e-17, 7.459505e-17, 7.461093e-17, 
    7.460218e-17, 7.459721e-17, 7.457753e-17, 7.457296e-17, 7.456906e-17, 
    7.456109e-17, 7.455102e-17, 7.453343e-17, 7.451797e-17, 7.450376e-17, 
    7.450478e-17, 7.450443e-17, 7.450137e-17, 7.45091e-17, 7.450008e-17, 
    7.449867e-17, 7.450252e-17, 7.447954e-17, 7.448609e-17, 7.447939e-17, 
    7.448362e-17, 7.459157e-17, 7.458625e-17, 7.458914e-17, 7.458376e-17, 
    7.458763e-17, 7.457072e-17, 7.456565e-17, 7.454171e-17, 7.455127e-17, 
    7.453578e-17, 7.454962e-17, 7.454722e-17, 7.45357e-17, 7.45488e-17, 
    7.451902e-17, 7.453959e-17, 7.450125e-17, 7.452214e-17, 7.449996e-17, 
    7.450382e-17, 7.449732e-17, 7.449162e-17, 7.448426e-17, 7.4471e-17, 
    7.447403e-17, 7.446279e-17, 7.457822e-17, 7.457142e-17, 7.457183e-17, 
    7.456458e-17, 7.455927e-17, 7.454752e-17, 7.452893e-17, 7.453586e-17, 
    7.452294e-17, 7.452042e-17, 7.453993e-17, 7.452813e-17, 7.456673e-17, 
    7.456068e-17, 7.456414e-17, 7.45778e-17, 7.453453e-17, 7.455683e-17, 
    7.451549e-17, 7.452751e-17, 7.449246e-17, 7.451006e-17, 7.447574e-17, 
    7.446161e-17, 7.444744e-17, 7.443194e-17, 7.456751e-17, 7.457214e-17, 
    7.456367e-17, 7.455231e-17, 7.454122e-17, 7.452682e-17, 7.452523e-17, 
    7.45226e-17, 7.451552e-17, 7.450968e-17, 7.452195e-17, 7.450819e-17, 
    7.455966e-17, 7.453251e-17, 7.457407e-17, 7.45618e-17, 7.455289e-17, 
    7.45566e-17, 7.45366e-17, 7.453196e-17, 7.451319e-17, 7.452279e-17, 
    7.446526e-17, 7.449068e-17, 7.441953e-17, 7.443948e-17, 7.457381e-17, 
    7.456743e-17, 7.454552e-17, 7.455591e-17, 7.452575e-17, 7.451842e-17, 
    7.45123e-17, 7.450481e-17, 7.450386e-17, 7.44994e-17, 7.450673e-17, 
    7.449961e-17, 7.452678e-17, 7.45146e-17, 7.454779e-17, 7.453982e-17, 
    7.454343e-17, 7.454752e-17, 7.45349e-17, 7.452181e-17, 7.452122e-17, 
    7.451706e-17, 7.450595e-17, 7.452562e-17, 7.446255e-17, 7.450197e-17, 
    7.456049e-17, 7.454865e-17, 7.454658e-17, 7.455123e-17, 7.451918e-17, 
    7.453081e-17, 7.449947e-17, 7.450786e-17, 7.449403e-17, 7.450092e-17, 
    7.450195e-17, 7.451075e-17, 7.451631e-17, 7.453034e-17, 7.454168e-17, 
    7.455051e-17, 7.454844e-17, 7.453872e-17, 7.452093e-17, 7.450391e-17, 
    7.450768e-17, 7.449508e-17, 7.452795e-17, 7.45143e-17, 7.451968e-17, 
    7.450562e-17, 7.453611e-17, 7.451107e-17, 7.454262e-17, 7.453979e-17, 
    7.453104e-17, 7.451359e-17, 7.450927e-17, 7.450522e-17, 7.450766e-17, 
    7.452042e-17, 7.452238e-17, 7.453118e-17, 7.453377e-17, 7.454039e-17, 
    7.454602e-17, 7.454095e-17, 7.45357e-17, 7.452029e-17, 7.450659e-17, 
    7.449159e-17, 7.448779e-17, 7.447108e-17, 7.448511e-17, 7.446239e-17, 
    7.448233e-17, 7.444752e-17, 7.450917e-17, 7.448231e-17, 7.453054e-17, 
    7.452526e-17, 7.451603e-17, 7.449426e-17, 7.450568e-17, 7.449219e-17, 
    7.452244e-17, 7.453854e-17, 7.454233e-17, 7.455003e-17, 7.454215e-17, 
    7.454278e-17, 7.453526e-17, 7.453766e-17, 7.451977e-17, 7.452936e-17, 
    7.450206e-17, 7.449221e-17, 7.446407e-17, 7.444706e-17, 7.442929e-17, 
    7.442162e-17, 7.441926e-17, 7.441829e-17 ;

 MEG_thujene_a =
  1.797621e-18, 1.797262e-18, 1.79733e-18, 1.797045e-18, 1.7972e-18, 
    1.797015e-18, 1.797545e-18, 1.79725e-18, 1.797437e-18, 1.797585e-18, 
    1.7965e-18, 1.797031e-18, 1.795922e-18, 1.796264e-18, 1.795397e-18, 
    1.795979e-18, 1.795279e-18, 1.795407e-18, 1.795005e-18, 1.79512e-18, 
    1.79462e-18, 1.794952e-18, 1.794351e-18, 1.794696e-18, 1.794644e-18, 
    1.794964e-18, 1.796918e-18, 1.796568e-18, 1.79694e-18, 1.79689e-18, 
    1.796911e-18, 1.7972e-18, 1.79735e-18, 1.797644e-18, 1.797589e-18, 
    1.797371e-18, 1.796867e-18, 1.797033e-18, 1.796601e-18, 1.796611e-18, 
    1.796135e-18, 1.79635e-18, 1.795547e-18, 1.795773e-18, 1.795115e-18, 
    1.795281e-18, 1.795124e-18, 1.795171e-18, 1.795123e-18, 1.795367e-18, 
    1.795263e-18, 1.795475e-18, 1.796311e-18, 1.796067e-18, 1.796799e-18, 
    1.79725e-18, 1.797534e-18, 1.79774e-18, 1.797711e-18, 1.797657e-18, 
    1.797369e-18, 1.797094e-18, 1.796887e-18, 1.796749e-18, 1.796612e-18, 
    1.796217e-18, 1.795993e-18, 1.795505e-18, 1.795587e-18, 1.795443e-18, 
    1.795297e-18, 1.795061e-18, 1.795099e-18, 1.794996e-18, 1.795442e-18, 
    1.795148e-18, 1.795635e-18, 1.795502e-18, 1.796598e-18, 1.796987e-18, 
    1.797173e-18, 1.797318e-18, 1.797689e-18, 1.797434e-18, 1.797535e-18, 
    1.79729e-18, 1.797138e-18, 1.797212e-18, 1.796745e-18, 1.796927e-18, 
    1.79598e-18, 1.796387e-18, 1.795314e-18, 1.795569e-18, 1.795252e-18, 
    1.795413e-18, 1.79514e-18, 1.795385e-18, 1.794956e-18, 1.794865e-18, 
    1.794928e-18, 1.79468e-18, 1.7954e-18, 1.795126e-18, 1.797215e-18, 
    1.797203e-18, 1.797145e-18, 1.797402e-18, 1.797417e-18, 1.797646e-18, 
    1.79744e-18, 1.797354e-18, 1.797127e-18, 1.796997e-18, 1.796872e-18, 
    1.796597e-18, 1.796294e-18, 1.795865e-18, 1.795553e-18, 1.795346e-18, 
    1.795471e-18, 1.795361e-18, 1.795485e-18, 1.795543e-18, 1.794901e-18, 
    1.795263e-18, 1.794716e-18, 1.794745e-18, 1.794995e-18, 1.794742e-18, 
    1.797194e-18, 1.797264e-18, 1.797514e-18, 1.797318e-18, 1.797671e-18, 
    1.797476e-18, 1.797366e-18, 1.796928e-18, 1.796827e-18, 1.79674e-18, 
    1.796563e-18, 1.796339e-18, 1.795948e-18, 1.795604e-18, 1.795288e-18, 
    1.795311e-18, 1.795303e-18, 1.795235e-18, 1.795407e-18, 1.795206e-18, 
    1.795175e-18, 1.79526e-18, 1.794749e-18, 1.794895e-18, 1.794746e-18, 
    1.79484e-18, 1.797241e-18, 1.797122e-18, 1.797187e-18, 1.797067e-18, 
    1.797153e-18, 1.796777e-18, 1.796664e-18, 1.796132e-18, 1.796345e-18, 
    1.796e-18, 1.796308e-18, 1.796254e-18, 1.795998e-18, 1.796289e-18, 
    1.795627e-18, 1.796085e-18, 1.795232e-18, 1.795697e-18, 1.795203e-18, 
    1.795289e-18, 1.795145e-18, 1.795018e-18, 1.794854e-18, 1.794559e-18, 
    1.794627e-18, 1.794377e-18, 1.796944e-18, 1.796793e-18, 1.796802e-18, 
    1.796641e-18, 1.796522e-18, 1.796261e-18, 1.795848e-18, 1.796002e-18, 
    1.795714e-18, 1.795658e-18, 1.796092e-18, 1.79583e-18, 1.796688e-18, 
    1.796554e-18, 1.796631e-18, 1.796934e-18, 1.795972e-18, 1.796468e-18, 
    1.795549e-18, 1.795816e-18, 1.795037e-18, 1.795428e-18, 1.794665e-18, 
    1.794351e-18, 1.794036e-18, 1.793691e-18, 1.796706e-18, 1.796809e-18, 
    1.79662e-18, 1.796367e-18, 1.796121e-18, 1.795801e-18, 1.795765e-18, 
    1.795707e-18, 1.795549e-18, 1.79542e-18, 1.795692e-18, 1.795386e-18, 
    1.796531e-18, 1.795927e-18, 1.796852e-18, 1.796579e-18, 1.79638e-18, 
    1.796463e-18, 1.796018e-18, 1.795915e-18, 1.795498e-18, 1.795711e-18, 
    1.794432e-18, 1.794997e-18, 1.793416e-18, 1.793859e-18, 1.796846e-18, 
    1.796704e-18, 1.796217e-18, 1.796448e-18, 1.795777e-18, 1.795614e-18, 
    1.795478e-18, 1.795311e-18, 1.79529e-18, 1.795191e-18, 1.795354e-18, 
    1.795196e-18, 1.7958e-18, 1.795529e-18, 1.796267e-18, 1.79609e-18, 
    1.79617e-18, 1.796261e-18, 1.795981e-18, 1.795689e-18, 1.795676e-18, 
    1.795584e-18, 1.795337e-18, 1.795774e-18, 1.794372e-18, 1.795248e-18, 
    1.79655e-18, 1.796286e-18, 1.79624e-18, 1.796343e-18, 1.795631e-18, 
    1.79589e-18, 1.795192e-18, 1.795379e-18, 1.795071e-18, 1.795225e-18, 
    1.795248e-18, 1.795443e-18, 1.795567e-18, 1.795879e-18, 1.796131e-18, 
    1.796328e-18, 1.796281e-18, 1.796065e-18, 1.79567e-18, 1.795291e-18, 
    1.795375e-18, 1.795095e-18, 1.795826e-18, 1.795522e-18, 1.795642e-18, 
    1.795329e-18, 1.796007e-18, 1.795451e-18, 1.796152e-18, 1.796089e-18, 
    1.795895e-18, 1.795506e-18, 1.79541e-18, 1.79532e-18, 1.795375e-18, 
    1.795659e-18, 1.795702e-18, 1.795898e-18, 1.795955e-18, 1.796102e-18, 
    1.796228e-18, 1.796115e-18, 1.795998e-18, 1.795656e-18, 1.795351e-18, 
    1.795017e-18, 1.794933e-18, 1.794561e-18, 1.794873e-18, 1.794368e-18, 
    1.794811e-18, 1.794037e-18, 1.795408e-18, 1.794811e-18, 1.795883e-18, 
    1.795766e-18, 1.795561e-18, 1.795077e-18, 1.795331e-18, 1.795031e-18, 
    1.795703e-18, 1.796061e-18, 1.796146e-18, 1.796317e-18, 1.796142e-18, 
    1.796155e-18, 1.795988e-18, 1.796042e-18, 1.795644e-18, 1.795857e-18, 
    1.79525e-18, 1.795031e-18, 1.794405e-18, 1.794027e-18, 1.793632e-18, 
    1.793462e-18, 1.793409e-18, 1.793388e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -2.856905e-25, 8.241083e-26, 1.730626e-25, -4.010655e-25, -6.592851e-26, 
    3.159079e-25, -2.747024e-25, 9.889298e-26, 8.515785e-26, -1.785565e-25, 
    -5.494041e-26, 7.142273e-26, -1.098802e-26, -2.472321e-25, 1.977859e-25, 
    -5.219339e-26, -8.240992e-27, 4.422711e-25, 4.752353e-25, 1.346043e-25, 
    5.494058e-26, 7.691677e-26, -1.648214e-25, -2.527262e-25, 1.04387e-25, 
    -5.439108e-25, -4.944636e-26, 5.219355e-26, 2.719555e-25, 1.346043e-25, 
    1.648216e-25, 3.296438e-26, 4.66995e-26, 1.840507e-25, -3.104137e-25, 
    2.554734e-25, 1.181221e-25, 1.730626e-25, -8.241074e-25, 2.032799e-25, 
    6.86757e-26, 2.664615e-25, -1.043869e-25, -1.20869e-25, 4.560062e-25, 
    1.922918e-25, -3.049197e-25, -3.735953e-25, -7.087323e-25, 3.653544e-25, 
    2.225091e-25, -1.620744e-25, -1.071339e-25, 3.955716e-25, 4.31283e-25, 
    -1.813036e-25, -2.3075e-25, -3.323899e-25, -1.23616e-25, -4.202947e-25, 
    2.005329e-25, 1.098818e-26, -1.703155e-25, -3.296421e-26, 3.378841e-25, 
    -3.735953e-25, 8.257462e-32, -2.36244e-25, 6.043463e-26, -6.318148e-26, 
    -1.263631e-25, -3.076667e-25, 1.510864e-25, -1.098809e-25, -2.527262e-25, 
    -4.944636e-26, 4.093068e-25, 4.477651e-25, -1.730625e-25, 2.14268e-25, 
    1.510864e-25, 1.400983e-25, 7.966372e-25, 1.840507e-25, -4.724882e-25, 
    1.703156e-25, -5.493967e-27, 1.840507e-25, 1.428454e-25, 2.197628e-26, 
    -1.098802e-26, -2.774494e-25, -1.785565e-25, -4.395231e-26, 
    -3.021719e-26, 2.527264e-25, 3.296438e-26, -2.472321e-25, -9.339876e-26, 
    2.17015e-25, -8.790471e-26, -1.813036e-25, 1.840507e-25, -2.966786e-25, 
    3.571133e-25, 2.032799e-25, -4.944636e-26, -2.774494e-25, 1.400983e-25, 
    -3.708483e-25, 2.225091e-25, -1.813036e-25, -9.614578e-26, 1.346043e-25, 
    -2.197612e-26, -1.071339e-25, -5.219339e-26, 5.164408e-25, -1.565803e-25, 
    1.373521e-26, 3.845843e-26, 2.856907e-25, -1.648214e-25, 2.747033e-26, 
    -3.021719e-26, -2.28003e-25, -1.098809e-25, -9.339876e-26, -7.142256e-26, 
    -3.021727e-25, -2.747024e-25, -7.691661e-26, 2.856907e-25, 1.620745e-25, 
    1.867978e-25, -3.653542e-25, -7.691661e-26, -1.373504e-26, -3.790893e-25, 
    2.527264e-25, -1.126279e-25, 1.071341e-25, 3.900776e-25, 2.747026e-25, 
    1.428454e-25, -3.131607e-25, -1.483393e-25, -2.582203e-25, -2.33497e-25, 
    4.230419e-25, 1.346043e-25, -6.043446e-26, -4.285358e-25, 1.318573e-25, 
    -2.36244e-25, -3.241488e-25, 1.675686e-25, -2.005327e-25, 2.472331e-26, 
    4.66995e-26, -1.373512e-25, 1.318573e-25, -6.78515e-25, 1.04387e-25, 
    2.197628e-26, -4.038125e-25, -2.609673e-25, 4.065598e-25, -1.922909e-26, 
    1.565805e-25, -1.950387e-25, 1.098811e-25, -5.548989e-25, -4.917174e-25, 
    -2.747016e-26, 5.76876e-26, 2.472323e-25, -1.648207e-26, -3.104137e-25, 
    2.747033e-26, -5.494041e-26, 3.159079e-25, -4.972114e-25, 1.098811e-25, 
    -2.664613e-25, -3.735953e-25, -2.774494e-25, -2.582203e-25, 1.648223e-26, 
    -1.373512e-25, -3.37884e-25, -1.620744e-25, -7.966364e-26, -2.747016e-26, 
    -1.565803e-25, -2.472321e-25, -1.098802e-26, 8.515785e-26, 2.060269e-25, 
    -1.785565e-25, -3.598602e-25, -6.867554e-26, -1.346041e-25, 1.813037e-25, 
    4.999586e-25, -3.626072e-25, 1.263632e-25, -3.131607e-25, -1.538333e-25, 
    2.472323e-25, 3.076668e-25, 5.494132e-27, -1.043869e-25, -1.922909e-26, 
    -1.20869e-25, -2.884375e-25, 2.472323e-25, 2.005329e-25, 1.04387e-25, 
    1.867978e-25, -6.318148e-26, -1.098809e-25, 1.126281e-25, 2.966788e-25, 
    -3.021727e-25, 5.494058e-26, -4.312828e-25, 1.730626e-25, -8.240992e-27, 
    4.395248e-26, 4.395248e-26, -1.648214e-25, 1.098818e-26, 8.515785e-26, 
    -5.054525e-25, 1.922918e-25, -1.510863e-25, -1.082328e-24, 8.241157e-27, 
    -2.527262e-25, -4.669934e-26, 2.362442e-25, -2.747024e-25, 4.395248e-26, 
    4.972116e-25, 4.889705e-25, -2.3075e-25, 4.66995e-26, 1.373513e-25, 
    4.944653e-26, 2.197621e-25, -3.296421e-26, -1.016398e-25, 1.373513e-25, 
    2.472331e-26, 4.779824e-25, 8.790487e-26, 4.889705e-25, -1.813036e-25, 
    -1.922916e-25, -7.416958e-26, -1.15375e-25, 6.86757e-26, -3.873304e-25, 
    7.142273e-26, 1.455924e-25, -3.186548e-25, 1.346043e-25, -1.373512e-25, 
    -3.323899e-25, 1.565805e-25, 3.735955e-25, 2.939317e-25, 2.280031e-25, 
    -5.493967e-27, 3.735955e-25, -3.873304e-25, -2.36244e-25, 4.175478e-25, 
    1.950388e-25, 3.378841e-25, -1.648214e-25, -3.46125e-25, 6.043463e-26, 
    3.26896e-25, 7.142273e-26, 5.219355e-26, -2.499792e-25, -1.703155e-25, 
    5.76876e-26, -4.120529e-26, -4.615001e-25, 5.356699e-25, -1.593274e-25, 
    2.197628e-26, 5.494132e-27, -1.318571e-25, 3.296431e-25, -2.25256e-25, 
    -2.389911e-25, -4.367769e-25, -2.197612e-26, 2.197628e-26, 2.252561e-25, 
    -4.862233e-25, 2.417383e-25, 1.04387e-25, 7.96638e-26, -4.615001e-25, 
    2.664615e-25, -1.867976e-25, -3.021727e-25, -8.515768e-26, -8.515768e-26, 
    2.719555e-25, -3.543661e-25, 7.142273e-26, -6.318156e-25, -3.43378e-25, 
    -5.219339e-26, 1.922926e-26, -5.988513e-25, 8.241157e-27, 1.208692e-25, 
    -2.25256e-25, 2.17015e-25, -6.75768e-25, -2.829435e-25, 1.0164e-25, 
    3.818365e-25, -4.148007e-25, 5.494058e-26, -4.944636e-26, -3.049197e-25, 
    1.620745e-25, -3.681012e-25, -4.395231e-26, 4.3403e-25 ;

 M_LITR2C_TO_LEACHING =
  -1.291101e-25, -4.944639e-26, -5.494044e-26, 2.74703e-26, 1.565805e-25, 
    -1.098805e-26, 1.373518e-26, -1.373507e-26, -2.225089e-25, -3.40631e-25, 
    -3.296424e-26, 4.395245e-26, 8.24108e-26, -1.648209e-26, 5.351427e-32, 
    2.005329e-25, -3.571127e-26, -1.648214e-25, 8.515782e-26, -9.889284e-26, 
    2.087739e-25, 9.889295e-26, 1.09881e-25, -2.966786e-25, -1.483393e-25, 
    -1.373512e-25, -1.730625e-25, -1.922917e-25, -1.648209e-26, 
    -1.648214e-25, 1.64822e-26, -2.170149e-25, 6.592865e-26, -8.515771e-26, 
    2.911847e-25, 5.351457e-32, -4.395234e-26, -6.043449e-26, 1.208691e-25, 
    -3.323899e-25, -4.669937e-26, 1.510864e-25, -2.637143e-25, -2.3075e-25, 
    -8.241069e-26, -7.966367e-26, 9.889295e-26, 1.648215e-25, -1.263631e-25, 
    -1.593274e-25, 3.296435e-26, -1.18122e-25, -1.648209e-26, -1.730625e-25, 
    8.790485e-26, -1.346042e-25, 1.510864e-25, 1.07134e-25, -1.098805e-26, 
    2.472323e-25, -3.818364e-25, 5.351453e-32, 3.021733e-26, -1.648209e-26, 
    -1.373507e-26, -4.395234e-26, -1.648214e-25, 6.592865e-26, -4.120532e-26, 
    -2.032798e-25, -2.115208e-25, 1.09881e-25, 1.565805e-25, -9.339879e-26, 
    5.219352e-26, 1.0164e-25, 3.296435e-26, 2.417382e-25, 9.065187e-26, 
    -1.840506e-25, -1.758095e-25, -3.296424e-26, -3.296424e-26, 
    -2.856905e-25, 3.296435e-26, 1.593275e-25, 5.494103e-27, 3.021728e-25, 
    -2.692084e-25, -1.071339e-25, 1.730626e-25, 9.614592e-26, 2.829436e-25, 
    -4.50512e-25, -1.15375e-25, 5.768757e-26, -1.977857e-25, -1.373512e-25, 
    1.208691e-25, 3.488722e-25, -4.944639e-26, 1.373518e-26, -1.236161e-25, 
    3.845835e-25, -2.032798e-25, -3.40631e-25, -6.867557e-26, -3.708483e-25, 
    -1.922912e-26, -1.291101e-25, 1.428453e-25, -2.747024e-25, -1.400982e-25, 
    -2.197614e-26, 8.241128e-27, 2.747025e-25, 6.318163e-26, 1.07134e-25, 
    -6.867557e-26, -1.098809e-25, 2.417382e-25, 1.373518e-26, -2.142679e-25, 
    -2.582203e-25, 3.84584e-26, 1.455924e-25, -1.18122e-25, 2.197625e-26, 
    -3.296429e-25, 3.84584e-26, 1.977858e-25, 1.0164e-25, -1.346042e-25, 
    -1.373512e-25, 1.758096e-25, -9.614581e-26, -2.142679e-25, 1.181221e-25, 
    4.94465e-26, -3.241489e-25, 4.94465e-26, 1.208691e-25, 5.494055e-26, 
    -8.790474e-26, -6.318152e-26, -3.571127e-26, -3.214019e-25, 1.64822e-26, 
    5.494103e-27, 3.296435e-26, 1.922923e-26, -7.142259e-26, -7.691664e-26, 
    -3.571127e-26, -2.197614e-26, -2.911846e-25, 1.09881e-25, -1.043869e-25, 
    -7.691664e-26, 1.977858e-25, -3.131608e-25, -1.922912e-26, 1.813037e-25, 
    8.24108e-26, 1.291102e-25, -8.241021e-27, 1.593275e-25, 1.04387e-25, 
    9.614592e-26, 6.318163e-26, 7.966377e-26, 3.571138e-26, -6.867557e-26, 
    1.64822e-26, -1.043869e-25, 6.04346e-26, -1.20869e-25, -4.669937e-26, 
    5.351419e-32, 1.09881e-25, 1.648215e-25, -1.098809e-25, -2.005328e-25, 
    -2.060268e-25, -1.373512e-25, 5.494055e-26, -5.493996e-27, -2.170149e-25, 
    -6.867557e-26, -3.021727e-25, -2.389911e-25, -7.691664e-26, 7.966377e-26, 
    -2.115208e-25, 1.09881e-25, 6.592865e-26, -2.142679e-25, -6.592854e-26, 
    4.312829e-25, -7.416961e-26, -8.241069e-26, 4.395245e-26, -2.801965e-25, 
    -1.510863e-25, -8.515771e-26, -1.043869e-25, -2.417381e-25, 1.263632e-25, 
    -5.494044e-26, 1.620745e-25, -2.25256e-25, 9.889295e-26, -4.669937e-26, 
    -1.840506e-25, 1.730626e-25, -7.966367e-26, -9.339879e-26, 7.416973e-26, 
    -3.021722e-26, 8.790485e-26, -1.428452e-25, 2.280031e-25, 1.346043e-25, 
    9.889295e-26, 6.04346e-26, -2.3075e-25, 1.263632e-25, -1.483393e-25, 
    8.515782e-26, 8.241128e-27, -7.966367e-26, -7.142259e-26, 5.494055e-26, 
    9.889295e-26, 5.35145e-32, 5.494103e-27, 1.373513e-25, 1.593275e-25, 
    2.252561e-25, 8.24108e-26, -4.944639e-26, -1.648209e-26, 3.571138e-26, 
    -7.691664e-26, -4.944639e-26, 2.829436e-25, 1.181221e-25, 1.153751e-25, 
    -2.087738e-25, -1.813036e-25, 5.494055e-26, -1.483393e-25, -1.263631e-25, 
    1.565805e-25, 6.592865e-26, 1.813037e-25, 5.494103e-27, 6.592865e-26, 
    2.307501e-25, 2.472328e-26, -1.922917e-25, -7.691664e-26, -2.746971e-27, 
    -3.461251e-25, 6.592865e-26, 8.241128e-27, -1.648209e-26, 2.472323e-25, 
    -2.362441e-25, 4.779824e-25, -3.323899e-25, 3.571138e-26, -1.922912e-26, 
    9.889295e-26, -1.18122e-25, -5.493996e-27, 6.04346e-26, 2.17015e-25, 
    1.922923e-26, -2.197619e-25, 6.04346e-26, -3.873304e-25, -1.758095e-25, 
    3.571138e-26, -7.691664e-26, -2.527262e-25, -9.339879e-26, 2.856906e-25, 
    -2.115208e-25, -2.170149e-25, -1.758095e-25, -3.845829e-26, 
    -1.483393e-25, 1.565805e-25, -1.675685e-25, -1.318571e-25, 7.416973e-26, 
    6.867567e-26, -1.950387e-25, -9.339879e-26, 3.84584e-26, -2.472322e-25, 
    -2.334971e-25, 7.966377e-26, 6.04346e-26, 8.515782e-26, 1.09881e-25, 
    1.0164e-25, 1.483394e-25, -2.911846e-25, 2.856906e-25, -9.614581e-26, 
    -3.296424e-26, -2.389911e-25, -9.889284e-26, 4.395245e-26, -2.472317e-26, 
    -1.263631e-25, -7.142259e-26, -4.944639e-26, -2.417381e-25, 5.494055e-26, 
    1.758096e-25, -6.043449e-26, -1.15375e-25, -9.065177e-26, -4.669937e-26, 
    1.64822e-26, -2.444852e-25, -2.225089e-25, -7.691664e-26, 2.14268e-25, 
    -2.417381e-25, 6.04346e-26, -3.021727e-25, -1.758095e-25, -1.593274e-25, 
    -1.483393e-25 ;

 M_LITR3C_TO_LEACHING =
  -2.197617e-26, 4.944647e-26, 5.494052e-26, 1.373515e-26, -1.607009e-25, 
    3.02173e-26, 6.867565e-26, -5.768749e-26, 5.494076e-27, -1.098807e-26, 
    -4.944642e-26, 1.098813e-26, -5.494023e-27, 1.057605e-25, -5.494023e-27, 
    9.065185e-26, -6.592857e-26, 7.142267e-26, -1.758096e-25, -7.142262e-26, 
    -8.241047e-27, -5.219344e-26, -2.197617e-26, -1.208691e-25, 
    -1.071339e-25, 9.889292e-26, 7.142267e-26, -2.060268e-25, -1.15375e-25, 
    8.241101e-27, 7.416969e-26, 7.416969e-26, 1.373539e-27, -2.609671e-26, 
    -5.219344e-26, 3.845837e-26, -9.889287e-26, -8.927828e-26, -4.532588e-26, 
    3.845837e-26, -1.922915e-26, -1.373512e-25, -3.433778e-26, -3.296427e-26, 
    -6.043452e-26, -4.395237e-26, 4.12054e-26, -5.494047e-26, -5.906101e-26, 
    -1.373512e-25, 9.339887e-26, 2.675714e-32, -1.428453e-25, -5.219344e-26, 
    -4.669939e-26, 4.395242e-26, -1.977858e-25, -6.867559e-26, 1.194956e-25, 
    -1.194956e-25, -7.142262e-26, 3.845837e-26, -3.159076e-26, -9.614584e-26, 
    1.428453e-25, -2.47232e-26, -6.730208e-26, -2.746998e-27, 2.060271e-26, 
    3.02173e-26, 1.181221e-25, 1.373513e-25, 5.494076e-27, -4.944642e-26, 
    -1.098807e-26, 6.867565e-26, -3.708481e-26, -5.768749e-26, -4.944642e-26, 
    1.593275e-25, -3.57113e-26, -3.021725e-26, -4.120535e-26, 4.944647e-26, 
    -1.37351e-26, -1.016399e-25, -9.614584e-26, -9.339881e-26, -1.18122e-25, 
    -8.515774e-26, 6.455511e-26, 1.730626e-25, 2.609676e-26, 1.098813e-26, 
    -1.37351e-26, -8.241071e-26, 5.494076e-27, 3.708486e-26, 3.159081e-26, 
    1.098813e-26, 1.373515e-26, -9.614584e-26, -2.884373e-26, 6.043457e-26, 
    -3.57113e-26, -3.845832e-26, -7.00491e-26, -5.494023e-27, 5.494052e-26, 
    -3.296427e-26, -5.219344e-26, -1.236161e-25, 1.373515e-26, 1.510864e-25, 
    2.747052e-27, -3.57113e-26, -5.494047e-26, -7.279613e-26, 5.21935e-26, 
    3.296432e-26, -1.455923e-25, -9.751935e-26, 6.730214e-26, 1.373515e-26, 
    -1.373486e-27, 1.373539e-27, -5.219344e-26, 8.241077e-26, 1.09881e-25, 
    -9.751935e-26, -5.494023e-27, -1.098807e-26, -7.966369e-26, 
    -8.241071e-26, -1.703155e-25, 4.944647e-26, 2.675728e-32, -1.648212e-26, 
    4.257891e-26, -2.060266e-26, 4.944647e-26, -1.455923e-25, -3.845832e-26, 
    -2.060266e-26, -2.746998e-27, -1.277366e-25, 5.494052e-26, -1.236158e-26, 
    3.983189e-26, -3.296427e-26, -1.854241e-25, 1.648217e-26, 4.395242e-26, 
    -1.648212e-26, -9.61456e-27, -2.334968e-26, 1.92292e-26, -1.002664e-25, 
    -1.593274e-25, 3.571135e-26, 8.927833e-26, -1.332307e-25, 8.515779e-26, 
    -6.318154e-26, -5.494023e-27, -3.983183e-26, 5.21935e-26, -3.57113e-26, 
    -5.768749e-26, -3.159076e-26, -1.085074e-25, -4.669939e-26, 1.153751e-25, 
    6.180808e-26, 1.098813e-26, -3.57113e-26, -1.043869e-25, -2.060266e-26, 
    -5.494047e-26, 8.378428e-26, -1.648212e-26, -5.631398e-26, -8.515774e-26, 
    -8.515774e-26, -9.339881e-26, 3.708486e-26, 5.21935e-26, 3.845837e-26, 
    -6.318154e-26, -1.098807e-26, 5.494052e-26, -3.159076e-26, 2.675718e-32, 
    -9.751935e-26, -1.071339e-25, 6.867589e-27, 6.31816e-26, -7.554316e-26, 
    -7.691667e-26, -1.455923e-25, 2.197622e-26, -1.263631e-25, 4.12054e-26, 
    -3.296427e-26, -1.455923e-25, 6.455511e-26, 6.592862e-26, -7.142262e-26, 
    -1.922915e-26, 1.455923e-25, -8.515774e-26, -1.085074e-25, 7.416969e-26, 
    -1.291101e-25, 7.554321e-26, -9.065179e-26, -1.236161e-25, 1.538334e-25, 
    -6.455506e-26, 5.768755e-26, -1.098807e-26, 3.571135e-26, 2.675724e-32, 
    9.75194e-26, 5.768755e-26, -1.236158e-26, -2.746998e-27, 3.159081e-26, 
    -1.758096e-25, -1.565804e-25, 1.098813e-26, 9.889292e-26, -7.142262e-26, 
    7.279618e-26, -2.609671e-26, 4.12054e-26, -7.691667e-26, -3.57113e-26, 
    -3.296427e-26, -4.669939e-26, -8.241047e-27, 1.57954e-25, -4.669939e-26, 
    3.296432e-26, -4.257886e-26, -6.867559e-26, -4.669939e-26, -4.120535e-26, 
    9.614589e-26, 6.867565e-26, -6.867535e-27, -1.922915e-26, -1.455923e-25, 
    -5.906101e-26, -4.669939e-26, -1.373486e-27, -1.208691e-25, 5.494076e-27, 
    -5.219344e-26, -6.867535e-27, -4.257886e-26, -1.785563e-26, 
    -3.983183e-26, -9.889287e-26, -1.236158e-26, 9.889292e-26, -1.304836e-25, 
    -3.296427e-26, -2.47232e-26, 2.675712e-32, -3.296427e-26, -4.669939e-26, 
    5.494076e-27, -2.47232e-26, -1.030134e-25, 5.494076e-27, -6.592857e-26, 
    -6.043452e-26, -1.455923e-25, -7.142262e-26, -1.15375e-25, -9.61456e-27, 
    -8.241047e-27, -1.071339e-25, -1.09881e-25, -1.208691e-25, -6.318154e-26, 
    -6.180803e-26, -4.120511e-27, -9.61456e-27, 1.648217e-26, 2.884379e-26, 
    7.691672e-26, 9.065185e-26, -2.884373e-26, -1.18122e-25, 3.845837e-26, 
    -1.09881e-25, -4.395237e-26, -8.790477e-26, 6.455511e-26, -1.016399e-25, 
    -1.373512e-25, -1.552069e-25, 2.747028e-26, -1.167485e-25, 1.373515e-26, 
    -9.889287e-26, -9.889287e-26, -1.030134e-25, -7.966369e-26, 
    -2.060266e-26, -2.334968e-26, -1.510863e-25, 9.614589e-26, 2.747028e-26, 
    1.346042e-25, -3.021725e-26, -1.016399e-25, -4.944642e-26, 2.334974e-26, 
    -6.592857e-26, -6.592857e-26, -7.966369e-26, 4.669945e-26, 1.222426e-25, 
    -7.142262e-26, 2.884379e-26, 7.142267e-26, -1.785563e-26, -8.378423e-26, 
    5.494052e-26, 8.241101e-27, -3.57113e-26, -2.47232e-26, 5.768755e-26, 
    1.030135e-25, -2.060266e-26 ;

 M_SOIL1C_TO_LEACHING =
  9.711808e-21, -1.421511e-20, -4.607863e-20, 3.909634e-21, 7.529425e-21, 
    6.995332e-21, 1.302991e-20, 2.963611e-20, 4.223174e-21, -1.623441e-20, 
    -1.356514e-20, 1.981068e-20, 4.890671e-21, -2.297752e-20, 2.283613e-21, 
    3.029855e-20, -2.522834e-20, -1.358238e-20, 3.474082e-20, 4.361404e-20, 
    1.765646e-21, -9.687756e-21, 1.370847e-20, -4.591407e-20, -1.780582e-20, 
    -9.365739e-21, -4.288734e-21, 2.42716e-20, -3.805472e-20, 1.407419e-21, 
    3.938723e-21, -1.703681e-20, -2.77605e-20, 1.525247e-20, 4.613742e-20, 
    1.719397e-20, -1.765172e-20, 4.798932e-20, -1.435718e-21, -2.759168e-21, 
    -2.00866e-20, -1.702944e-20, 1.132702e-20, -1.095695e-20, -7.489819e-21, 
    -3.18649e-20, 3.696707e-21, -3.378626e-21, 5.371329e-21, -5.689671e-21, 
    1.716798e-20, -6.738024e-21, 6.877153e-21, -3.695094e-20, -4.68123e-20, 
    5.458683e-20, 1.326407e-20, 2.271456e-21, 2.321228e-21, -3.872278e-20, 
    -1.696016e-20, -5.580993e-20, 2.470274e-20, 3.233309e-21, -5.511264e-21, 
    -6.325507e-21, -3.252647e-20, 1.298441e-20, -5.019405e-20, -2.521646e-20, 
    1.423069e-20, 1.556944e-20, 3.020721e-20, 2.634768e-21, -4.509045e-20, 
    4.241028e-22, 2.433754e-21, -6.0626e-21, 1.046132e-20, -5.684013e-21, 
    -2.439403e-20, 1.318657e-21, -2.456507e-20, -4.316165e-21, 3.127061e-20, 
    4.613035e-21, -5.505044e-21, 6.206521e-21, -3.180724e-20, -2.791712e-20, 
    -1.563077e-20, 4.48883e-20, -1.912872e-20, 2.206855e-20, -1.03273e-20, 
    -1.82268e-20, 2.576922e-20, 1.94861e-20, 1.818526e-21, 2.845177e-20, 
    2.212794e-20, -1.208929e-20, 2.883231e-20, -2.842604e-20, -3.16931e-22, 
    -5.480446e-21, 1.241216e-20, 3.987635e-21, 7.863882e-21, 2.758972e-20, 
    -9.38072e-21, -1.800628e-20, 6.004634e-21, 1.955536e-20, -1.936931e-20, 
    4.751488e-20, 4.292056e-22, -3.546858e-20, -5.071455e-20, 1.270338e-20, 
    1.601243e-20, 2.339654e-20, -1.884428e-21, -5.470279e-21, 1.277951e-21, 
    -1.513429e-20, 8.351888e-21, 4.518999e-20, 3.951642e-20, 2.675256e-20, 
    1.495982e-20, 9.532829e-21, 2.259642e-20, -1.118623e-20, 4.960766e-20, 
    2.767256e-20, -5.421368e-21, 1.584963e-20, -1.382266e-21, 3.915454e-20, 
    2.688319e-20, -3.892581e-20, -1.572209e-20, -2.279605e-20, -1.133637e-20, 
    -4.267816e-21, 3.39701e-20, -1.998877e-20, 2.893193e-21, -1.909566e-21, 
    -1.279554e-20, -2.751535e-20, -3.042606e-20, 2.05155e-20, -2.879216e-20, 
    1.535792e-20, 3.003729e-21, -1.190568e-21, -1.248534e-21, -1.599888e-20, 
    -5.960253e-21, -3.076083e-20, -1.847353e-21, 1.019754e-20, -9.367445e-21, 
    1.779651e-20, 5.541601e-22, 1.21283e-20, 2.322267e-20, 3.332823e-21, 
    3.971971e-20, 1.186848e-20, -2.308216e-20, -1.662937e-20, -7.851415e-21, 
    2.772317e-20, -1.238502e-20, -5.445334e-22, 8.582292e-21, -1.611274e-21, 
    1.093434e-20, 1.453378e-20, 2.738726e-20, -5.595242e-22, 1.131035e-20, 
    -1.131093e-20, 3.151996e-20, -1.207542e-20, 1.763674e-20, -2.246439e-20, 
    9.065211e-21, 9.30889e-21, -3.95413e-20, 2.206062e-20, 7.235353e-21, 
    1.226712e-20, -1.913691e-20, 1.707072e-20, 3.674512e-20, 5.527441e-20, 
    4.50926e-21, -5.602085e-20, 7.712898e-22, -4.029225e-20, -2.473414e-20, 
    -1.851209e-20, -2.730246e-20, 3.918351e-21, 3.597184e-21, 4.510966e-21, 
    -8.422272e-21, 3.401448e-20, -8.860784e-21, -9.171785e-22, 1.17237e-20, 
    1.067819e-20, 1.317186e-20, 1.57286e-20, -3.840039e-21, 1.387503e-20, 
    -2.24491e-20, 1.127276e-20, 2.66485e-20, 1.987766e-20, -1.139152e-20, 
    2.026444e-20, -4.918381e-21, 3.374392e-20, 1.362225e-20, -3.532147e-21, 
    4.03938e-21, -2.003317e-20, -6.012015e-21, 6.981271e-23, -6.342813e-20, 
    9.278928e-21, 3.674481e-20, 2.099163e-20, -3.379963e-20, -3.112575e-21, 
    2.780117e-21, 2.846166e-20, -1.286678e-20, 4.254542e-21, -2.019885e-20, 
    9.776256e-21, 3.502243e-20, 2.536604e-20, 1.625051e-20, 7.547214e-21, 
    2.198205e-20, -8.379026e-21, 5.555631e-20, 9.171619e-22, -4.342802e-20, 
    4.782929e-20, -2.255543e-20, 1.748634e-20, 4.045312e-20, 2.909864e-21, 
    -2.120339e-20, 1.798253e-20, -3.723846e-20, 4.087382e-20, 3.103819e-20, 
    6.590724e-21, -2.331086e-20, 6.323304e-21, 8.362901e-21, 3.120697e-20, 
    3.948339e-21, 1.171357e-21, 1.402855e-20, -1.337606e-21, -3.304019e-20, 
    2.012872e-20, 1.413146e-20, 5.376676e-21, -7.956613e-21, 9.520111e-21, 
    2.221333e-20, 8.961469e-21, 1.30633e-20, 3.076534e-20, -3.192014e-21, 
    9.344821e-21, -1.925481e-20, 1.126087e-20, 3.528764e-20, 1.463244e-20, 
    1.114919e-20, -1.102538e-20, -8.512169e-21, -2.333378e-20, 4.075792e-20, 
    3.36639e-20, 5.4854e-20, 3.309789e-20, -4.066263e-20, 1.302514e-20, 
    -9.055023e-21, -1.310175e-21, -3.752571e-20, -1.266803e-20, -1.76096e-20, 
    2.680713e-20, 9.43814e-21, 2.75705e-20, 3.921843e-20, -2.607908e-20, 
    -2.21839e-20, 2.601803e-20, 1.530365e-20, -1.350238e-20, 8.149429e-21, 
    -3.605944e-21, -3.172211e-20, -1.345232e-20, 3.458366e-21, 1.079778e-20, 
    3.076762e-20, -1.996702e-20, -2.829291e-21, 4.436582e-20, -1.57467e-20, 
    -2.365268e-20, -7.176562e-21, 1.695168e-20, 1.573511e-20, -2.289412e-20, 
    -2.296707e-20, -5.162383e-20, -1.795256e-20, -1.127134e-20, 1.459994e-20, 
    -7.75955e-21, -1.043151e-22, -9.375356e-21 ;

 M_SOIL2C_TO_LEACHING =
  -1.89913e-20, -2.391054e-20, 1.448487e-20, -1.433303e-20, 1.103101e-20, 
    -1.567658e-20, 1.238616e-20, 4.970689e-21, -1.361631e-20, 3.755796e-20, 
    -5.456197e-20, -4.009603e-20, -1.040958e-20, -1.926048e-20, 
    -2.732029e-21, 1.500649e-20, 5.753564e-21, -3.865466e-20, -1.973205e-20, 
    -2.516296e-21, 4.131545e-20, 2.761489e-20, -6.664244e-21, -4.596354e-20, 
    -2.20301e-20, 1.564547e-20, 5.80531e-21, 4.106652e-21, -2.946027e-20, 
    4.296971e-20, 2.112865e-21, 1.646878e-20, -1.74985e-20, -6.534758e-21, 
    -2.568753e-20, 2.510932e-21, -9.382998e-21, -1.53404e-20, 1.264174e-20, 
    -4.086585e-21, 1.095806e-20, -1.034625e-20, 1.255749e-20, -1.394161e-21, 
    3.722205e-20, -2.213048e-20, 1.896585e-20, -3.51559e-20, 1.286737e-20, 
    -1.972923e-20, -1.25903e-20, -1.008134e-20, -4.628021e-20, 6.941601e-21, 
    1.519116e-21, -8.821767e-21, -2.782634e-20, -7.648442e-21, 4.306833e-21, 
    -2.826262e-20, 4.823048e-20, -1.740688e-20, -1.366891e-20, 1.358551e-20, 
    -2.007121e-21, -2.87065e-20, 1.011883e-21, 3.799675e-20, -1.48151e-20, 
    1.074096e-21, 1.471339e-21, 2.972575e-20, 2.41367e-21, -2.096619e-20, 
    2.563974e-20, -3.234017e-20, 2.196198e-20, -1.193433e-20, -2.307196e-20, 
    -2.56646e-20, 7.128759e-21, -3.501706e-20, 7.826556e-21, -5.10086e-20, 
    1.246333e-20, 2.960492e-21, -4.88033e-20, -6.510444e-21, 1.973376e-20, 
    1.711932e-21, -1.036095e-20, -2.194075e-20, 1.430476e-20, -2.264974e-21, 
    2.682097e-20, -1.744308e-20, -2.697534e-20, 3.224827e-21, -2.589477e-20, 
    -4.375994e-20, 4.463923e-20, -2.14556e-20, -4.21362e-20, -2.526485e-21, 
    2.239598e-20, 2.570899e-20, 1.006749e-20, 2.98479e-20, -7.039141e-21, 
    3.255276e-20, 7.732119e-21, 1.612978e-20, -8.647329e-21, 1.181928e-20, 
    2.062098e-20, 2.559019e-21, 8.467788e-21, 1.186422e-20, -2.3746e-20, 
    -1.561804e-20, -3.476231e-20, -1.922624e-20, -9.311741e-21, 4.477778e-20, 
    2.356589e-20, -2.341266e-20, 2.955779e-20, -5.422409e-20, -3.582748e-21, 
    -1.743713e-20, 3.323795e-21, -7.823159e-21, 3.635917e-21, -1.70563e-20, 
    -5.043523e-20, -1.450975e-20, -1.2251e-20, 3.917495e-21, -2.196677e-20, 
    2.404513e-20, 2.275984e-20, -1.029788e-20, -2.523088e-21, 2.445565e-20, 
    4.626465e-20, -2.463376e-20, -6.981206e-21, -2.247173e-20, -4.826159e-20, 
    -7.927785e-21, 1.980642e-20, -3.113147e-21, 4.855646e-20, -1.010765e-21, 
    -3.277386e-20, -7.997336e-21, 2.341579e-21, 1.400394e-20, 7.018796e-21, 
    8.676157e-21, 2.825441e-20, 1.434859e-20, 8.503409e-21, -1.73919e-20, 
    2.382092e-20, -4.533034e-21, 1.012402e-20, -3.720878e-20, 2.25735e-20, 
    -7.270427e-21, -4.002056e-20, 4.810522e-20, -9.837308e-21, -1.533587e-20, 
    1.645751e-20, 1.848862e-20, 4.548036e-20, 1.339775e-20, -1.223829e-20, 
    1.073616e-20, 2.588458e-20, -3.497099e-21, -6.02698e-21, -1.461237e-20, 
    5.830196e-21, -1.860652e-20, -4.658981e-20, -1.233496e-20, 4.2292e-20, 
    3.978643e-20, 1.282016e-20, -1.958872e-20, 5.179676e-22, 1.788641e-20, 
    -9.99453e-21, 1.99721e-20, 1.488634e-20, 7.246669e-21, -2.035773e-20, 
    -3.529864e-20, 1.436131e-20, -1.877332e-20, -3.345893e-20, 2.092433e-20, 
    4.537826e-21, -1.302174e-20, 2.88355e-21, -2.391308e-20, 1.163805e-20, 
    -1.378624e-20, -6.227984e-21, 7.864455e-21, 5.056366e-21, -4.14002e-21, 
    -2.015051e-20, -3.629073e-20, -3.147584e-20, 2.856686e-20, -6.138911e-21, 
    -1.839476e-20, -1.034709e-20, 4.240482e-20, 3.944095e-20, 3.351941e-20, 
    2.973225e-20, 5.834709e-21, 2.033687e-21, -1.81236e-20, 6.527966e-21, 
    1.135279e-20, 5.135822e-21, 9.859671e-21, 4.927998e-21, 9.000174e-21, 
    -2.686366e-20, -3.876248e-21, -5.33838e-20, -3.378351e-20, 5.269422e-20, 
    1.720048e-20, 3.595477e-21, -1.211982e-20, 3.369866e-21, 1.996813e-20, 
    2.678423e-20, 2.753375e-20, -7.874333e-21, 1.617813e-20, 6.451361e-21, 
    -2.508754e-20, 2.978089e-20, 2.02472e-20, -1.542858e-21, -1.058093e-20, 
    5.975234e-21, 5.268773e-20, 4.467101e-22, -4.468847e-21, 4.210737e-20, 
    9.197521e-21, -1.493782e-20, -4.007426e-20, -4.085752e-21, -2.653372e-20, 
    1.547385e-20, -3.651754e-21, -3.674312e-20, -2.804121e-21, -4.646963e-20, 
    -2.069569e-21, -9.110988e-21, -2.784448e-20, -3.14931e-20, 8.093725e-21, 
    -2.176163e-21, -1.878011e-20, 4.071321e-20, -2.491141e-20, 2.752102e-20, 
    -1.176328e-20, 5.212427e-21, 4.200783e-20, -1.262167e-20, 2.82499e-20, 
    -6.245227e-21, 1.948918e-20, 2.842659e-20, 2.70486e-20, 8.8605e-21, 
    1.789572e-20, 8.058095e-21, 1.343877e-20, -7.099958e-21, -2.660241e-20, 
    -4.418791e-21, 4.074772e-20, 3.561253e-21, 1.483319e-20, 2.440222e-20, 
    -6.976721e-20, -4.574018e-21, 1.460588e-20, -8.330677e-21, 9.25178e-21, 
    -3.229913e-21, -1.706255e-20, -5.929146e-21, 1.302483e-20, 4.385975e-20, 
    1.662344e-20, 2.830729e-20, -9.560523e-21, 1.059138e-20, 9.671941e-21, 
    -1.734016e-20, -4.917649e-20, -1.594488e-20, 1.721265e-21, -2.490586e-21, 
    -2.868616e-20, 8.112412e-21, -2.007502e-20, 2.179298e-21, -5.10951e-20, 
    4.801909e-21, 4.124079e-20, 3.132669e-21, 1.300194e-20, -1.567827e-20, 
    -4.894011e-22, -2.035012e-20, 4.363725e-20, 8.619881e-21, -2.227239e-20, 
    2.798757e-21, 1.202853e-20, -1.915898e-20, 3.756164e-20 ;

 M_SOIL3C_TO_LEACHING =
  5.815942e-20, -1.663446e-20, 3.248291e-21, 1.443426e-20, -2.162864e-20, 
    -1.818214e-20, -8.810444e-21, 1.723077e-20, 1.763957e-20, -2.757587e-20, 
    1.775182e-20, -1.610547e-20, -2.85151e-20, 7.919459e-22, 1.56709e-20, 
    -2.541524e-20, -2.48719e-21, -2.547883e-20, -1.464717e-20, 4.265135e-20, 
    4.202227e-20, -1.756719e-20, 2.371258e-21, -3.163361e-20, 1.130944e-21, 
    -1.802552e-20, 3.589916e-20, -3.591132e-20, 8.773402e-21, 7.489247e-21, 
    8.14093e-21, 3.151261e-20, 3.622261e-20, 8.943915e-21, 1.102961e-20, 
    2.046093e-20, 2.993187e-20, 3.173484e-20, -6.214692e-21, 3.612706e-20, 
    -2.841389e-20, -2.217683e-20, 4.904049e-20, -5.837812e-21, 1.09759e-20, 
    -6.528276e-21, -8.793201e-21, -3.192936e-20, -2.213045e-20, 8.74006e-21, 
    -2.32517e-21, 2.647518e-20, -2.862452e-20, 3.459465e-20, 4.009391e-21, 
    -1.669527e-20, -4.943551e-21, -1.806424e-20, -1.362028e-20, 7.517813e-21, 
    -1.506927e-20, -5.680616e-21, 7.215008e-21, 8.745146e-21, 4.040498e-21, 
    -1.367736e-20, -1.759236e-20, 7.973023e-21, -2.856655e-20, -5.371785e-22, 
    1.809843e-20, -1.118477e-21, 5.369622e-21, 5.051263e-21, 1.271452e-21, 
    7.333186e-21, 1.39635e-20, 1.173278e-20, 4.176386e-20, 1.164935e-20, 
    3.938043e-20, 3.601116e-20, -1.879481e-20, -8.341699e-21, 6.076464e-21, 
    2.546473e-20, -1.718468e-20, 2.159187e-20, 3.031863e-20, -1.630677e-20, 
    -1.247578e-20, 4.387786e-20, 5.580314e-20, -4.474272e-20, -2.036877e-20, 
    6.464357e-21, -7.14206e-22, 5.919268e-21, -1.874081e-20, 2.955952e-21, 
    1.414615e-20, -1.255343e-21, -1.137998e-21, 9.733582e-21, -1.393185e-20, 
    -3.32266e-21, -2.670901e-20, -3.845992e-21, -3.969371e-20, 2.405869e-20, 
    -5.280929e-20, 1.044041e-20, -3.39031e-20, -2.867173e-21, -1.412609e-20, 
    5.934821e-21, 2.933645e-20, -2.004575e-21, -1.713576e-20, 1.021591e-20, 
    6.774528e-21, -8.131051e-21, 3.272155e-20, -1.156948e-21, 1.008839e-20, 
    -2.413106e-20, -1.69644e-20, 2.28325e-20, -1.126908e-20, 2.222574e-20, 
    1.634212e-20, -6.488099e-21, 6.106409e-21, 1.090435e-20, 4.695224e-20, 
    -2.379038e-20, -1.292194e-20, -1.392757e-20, -3.909868e-21, 2.095601e-20, 
    4.116842e-21, -1.337598e-20, -1.566385e-20, -9.777963e-21, -1.114638e-20, 
    1.018029e-20, 2.273042e-20, -5.893526e-21, -1.252497e-20, 1.316735e-20, 
    1.73485e-21, 3.001187e-20, -1.790082e-20, -5.230804e-21, 1.604781e-20, 
    -1.362054e-20, -8.262243e-21, 1.25866e-20, 2.939098e-20, -5.005579e-23, 
    8.67673e-21, 5.884728e-20, -1.702053e-21, 2.219604e-20, -1.061964e-20, 
    -1.119106e-20, -5.252578e-21, -3.795936e-21, -9.201751e-21, 
    -1.107427e-20, -1.365108e-20, 1.75785e-20, 2.279885e-20, -2.84478e-20, 
    -2.077393e-20, 6.435808e-21, 3.639859e-21, 3.614601e-20, -8.544965e-21, 
    -5.278047e-20, -1.541817e-20, -4.569891e-20, 5.871491e-21, -1.144791e-21, 
    -3.099577e-20, 1.254222e-20, 6.10726e-21, 7.779324e-21, -3.892214e-20, 
    1.838626e-20, -1.159818e-20, -1.744562e-20, 4.733251e-20, -9.030709e-21, 
    -2.448873e-20, 7.054694e-21, -3.110152e-20, 2.995333e-20, -1.219218e-20, 
    -2.813879e-20, 1.238673e-20, -1.444471e-20, -2.673275e-20, 9.644803e-21, 
    -9.273842e-21, -3.994949e-22, 4.132084e-21, -1.159818e-20, 1.976881e-20, 
    -1.072426e-20, -2.124989e-21, 1.769328e-20, -1.896983e-20, 3.822351e-20, 
    1.416653e-20, -3.006557e-20, -4.144888e-20, -1.941258e-20, 3.699558e-21, 
    -1.84445e-20, -2.643023e-20, 3.46136e-20, -1.128322e-20, 2.624478e-20, 
    -2.420827e-20, 1.047066e-20, 1.806481e-20, 3.367606e-20, -2.63802e-20, 
    4.56129e-21, 2.229354e-21, 3.085669e-20, 3.664483e-21, 1.958336e-20, 
    -1.888245e-20, -1.011186e-20, 3.332277e-21, -1.662344e-20, -1.611274e-21, 
    -1.882592e-20, 7.866118e-21, -3.866456e-20, -6.423633e-21, -6.291314e-21, 
    -3.060872e-20, -2.47149e-20, -1.391456e-20, -1.455045e-20, 7.372203e-21, 
    -2.92912e-20, 1.720728e-20, 9.7053e-21, -2.181691e-20, -8.065459e-21, 
    -1.99805e-21, 5.166339e-21, -1.27233e-22, -1.792908e-20, 3.234439e-20, 
    3.973809e-20, 1.0059e-20, -2.463659e-20, 3.056234e-20, -2.031701e-20, 
    8.797732e-21, -5.551425e-21, 3.311483e-20, -1.642381e-21, 8.771712e-21, 
    -3.637389e-20, -1.026087e-20, -5.710016e-21, -2.45399e-20, 4.265614e-20, 
    -1.522306e-20, 1.53212e-20, -1.879481e-20, -3.228531e-20, -2.630228e-21, 
    -1.10576e-20, 2.439882e-20, 3.737956e-20, 2.084861e-21, -4.028406e-20, 
    -2.625523e-20, -3.026293e-20, -6.059204e-21, -1.839645e-20, 
    -3.211116e-20, -2.614015e-20, 2.246579e-20, -1.140282e-20, 4.123882e-20, 
    -5.538402e-21, 1.666217e-20, -8.32897e-21, -2.074849e-20, 7.004949e-21, 
    -4.315094e-20, -1.896837e-21, 1.894467e-20, -9.057847e-21, -1.398442e-20, 
    2.001806e-22, 2.875996e-20, 2.510564e-20, 1.464969e-20, 5.430952e-21, 
    -2.113384e-20, -2.823971e-20, 3.267773e-20, -8.74006e-21, 1.666217e-20, 
    -1.76096e-20, 2.014288e-20, 1.613318e-20, 3.631949e-21, -2.534673e-21, 
    2.271544e-20, -3.244322e-21, 1.99277e-20, -2.023392e-20, 2.46202e-21, 
    -1.923472e-20, -1.047801e-20, 2.335467e-20, 1.893441e-21, -1.289816e-20, 
    1.386794e-20, 3.113487e-20, 1.217805e-20, -1.867382e-20, -2.004702e-20, 
    -6.462667e-21, 5.956285e-21, -5.78214e-21, 5.266451e-21, -3.504808e-23 ;

 NBP =
  -6.35757e-08, -6.385525e-08, -6.38009e-08, -6.402639e-08, -6.39013e-08, 
    -6.404895e-08, -6.363237e-08, -6.386636e-08, -6.371698e-08, 
    -6.360087e-08, -6.446398e-08, -6.403645e-08, -6.490803e-08, 
    -6.463537e-08, -6.532027e-08, -6.48656e-08, -6.541195e-08, -6.530715e-08, 
    -6.562256e-08, -6.55322e-08, -6.593564e-08, -6.566426e-08, -6.614476e-08, 
    -6.587083e-08, -6.591368e-08, -6.565531e-08, -6.412248e-08, 
    -6.441075e-08, -6.41054e-08, -6.41465e-08, -6.412806e-08, -6.390389e-08, 
    -6.379093e-08, -6.355432e-08, -6.359728e-08, -6.377105e-08, 
    -6.416499e-08, -6.403126e-08, -6.436827e-08, -6.436066e-08, 
    -6.473585e-08, -6.456669e-08, -6.519728e-08, -6.501806e-08, 
    -6.553597e-08, -6.540572e-08, -6.552985e-08, -6.549221e-08, 
    -6.553034e-08, -6.533932e-08, -6.542116e-08, -6.525307e-08, 
    -6.459837e-08, -6.479079e-08, -6.421691e-08, -6.387185e-08, 
    -6.364264e-08, -6.347999e-08, -6.350298e-08, -6.354682e-08, 
    -6.377207e-08, -6.398385e-08, -6.414524e-08, -6.42532e-08, -6.435957e-08, 
    -6.468156e-08, -6.485197e-08, -6.523353e-08, -6.516466e-08, 
    -6.528133e-08, -6.539276e-08, -6.557987e-08, -6.554907e-08, -6.56315e-08, 
    -6.527824e-08, -6.551303e-08, -6.512544e-08, -6.523145e-08, 
    -6.438852e-08, -6.406734e-08, -6.393085e-08, -6.381136e-08, 
    -6.352067e-08, -6.372141e-08, -6.364228e-08, -6.383054e-08, 
    -6.395017e-08, -6.3891e-08, -6.425615e-08, -6.411419e-08, -6.486207e-08, 
    -6.453993e-08, -6.537977e-08, -6.51788e-08, -6.542793e-08, -6.53008e-08, 
    -6.551863e-08, -6.532259e-08, -6.566219e-08, -6.573613e-08, -6.56856e-08, 
    -6.587971e-08, -6.531172e-08, -6.552985e-08, -6.388935e-08, 
    -6.389899e-08, -6.394394e-08, -6.374634e-08, -6.373425e-08, 
    -6.355315e-08, -6.371429e-08, -6.378291e-08, -6.39571e-08, -6.406013e-08, 
    -6.415808e-08, -6.437342e-08, -6.461393e-08, -6.495023e-08, 
    -6.519183e-08, -6.535377e-08, -6.525447e-08, -6.534214e-08, 
    -6.524414e-08, -6.519819e-08, -6.570843e-08, -6.542193e-08, 
    -6.585179e-08, -6.5828e-08, -6.563347e-08, -6.583068e-08, -6.390577e-08, 
    -6.385024e-08, -6.365745e-08, -6.380832e-08, -6.353343e-08, -6.36873e-08, 
    -6.377579e-08, -6.411717e-08, -6.419216e-08, -6.426171e-08, 
    -6.439907e-08, -6.457535e-08, -6.488458e-08, -6.515364e-08, 
    -6.539925e-08, -6.538125e-08, -6.538759e-08, -6.544246e-08, 
    -6.530654e-08, -6.546477e-08, -6.549133e-08, -6.542189e-08, 
    -6.582482e-08, -6.570971e-08, -6.58275e-08, -6.575254e-08, -6.386828e-08, 
    -6.396172e-08, -6.391124e-08, -6.400618e-08, -6.393929e-08, 
    -6.423671e-08, -6.432588e-08, -6.474312e-08, -6.457188e-08, 
    -6.484441e-08, -6.459956e-08, -6.464295e-08, -6.485331e-08, 
    -6.461279e-08, -6.513881e-08, -6.47822e-08, -6.544459e-08, -6.508849e-08, 
    -6.546691e-08, -6.539818e-08, -6.551196e-08, -6.561386e-08, 
    -6.574206e-08, -6.59786e-08, -6.592382e-08, -6.612164e-08, -6.410102e-08, 
    -6.422221e-08, -6.421153e-08, -6.433836e-08, -6.443215e-08, 
    -6.463544e-08, -6.496149e-08, -6.483888e-08, -6.506396e-08, 
    -6.510916e-08, -6.476719e-08, -6.497716e-08, -6.430331e-08, 
    -6.441219e-08, -6.434736e-08, -6.411058e-08, -6.486714e-08, 
    -6.447888e-08, -6.519582e-08, -6.498549e-08, -6.559934e-08, 
    -6.529406e-08, -6.589367e-08, -6.615002e-08, -6.639124e-08, 
    -6.667317e-08, -6.428834e-08, -6.4206e-08, -6.435344e-08, -6.455743e-08, 
    -6.47467e-08, -6.499832e-08, -6.502406e-08, -6.507121e-08, -6.51933e-08, 
    -6.529596e-08, -6.508611e-08, -6.532169e-08, -6.443745e-08, 
    -6.490084e-08, -6.417487e-08, -6.439348e-08, -6.454541e-08, 
    -6.447876e-08, -6.482487e-08, -6.490644e-08, -6.523793e-08, 
    -6.506657e-08, -6.608675e-08, -6.56354e-08, -6.688783e-08, -6.653783e-08, 
    -6.417723e-08, -6.428806e-08, -6.467379e-08, -6.449026e-08, 
    -6.501512e-08, -6.514431e-08, -6.524932e-08, -6.538358e-08, 
    -6.539807e-08, -6.547761e-08, -6.534727e-08, -6.547246e-08, 
    -6.499886e-08, -6.52105e-08, -6.46297e-08, -6.477106e-08, -6.470603e-08, 
    -6.463469e-08, -6.485485e-08, -6.508942e-08, -6.509442e-08, 
    -6.516963e-08, -6.53816e-08, -6.501724e-08, -6.614502e-08, -6.544855e-08, 
    -6.440892e-08, -6.46224e-08, -6.465288e-08, -6.457019e-08, -6.513136e-08, 
    -6.492802e-08, -6.547567e-08, -6.532766e-08, -6.557018e-08, 
    -6.544967e-08, -6.543194e-08, -6.527716e-08, -6.51808e-08, -6.493735e-08, 
    -6.473926e-08, -6.458218e-08, -6.46187e-08, -6.479126e-08, -6.510376e-08, 
    -6.539939e-08, -6.533463e-08, -6.555175e-08, -6.497706e-08, 
    -6.521804e-08, -6.512491e-08, -6.536776e-08, -6.483562e-08, 
    -6.528879e-08, -6.471979e-08, -6.476968e-08, -6.492399e-08, -6.52344e-08, 
    -6.530306e-08, -6.537638e-08, -6.533113e-08, -6.51117e-08, -6.507574e-08, 
    -6.492024e-08, -6.487731e-08, -6.475882e-08, -6.466072e-08, 
    -6.475035e-08, -6.484448e-08, -6.511178e-08, -6.535268e-08, 
    -6.561532e-08, -6.567959e-08, -6.598647e-08, -6.573666e-08, -6.61489e-08, 
    -6.579844e-08, -6.64051e-08, -6.531504e-08, -6.578811e-08, -6.493101e-08, 
    -6.502334e-08, -6.519036e-08, -6.557342e-08, -6.536661e-08, 
    -6.560847e-08, -6.507433e-08, -6.479721e-08, -6.47255e-08, -6.459173e-08, 
    -6.472856e-08, -6.471743e-08, -6.484837e-08, -6.480629e-08, 
    -6.512066e-08, -6.49518e-08, -6.54315e-08, -6.560656e-08, -6.610091e-08, 
    -6.640397e-08, -6.671245e-08, -6.684864e-08, -6.689009e-08, -6.690742e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371698e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441075e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379093e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377207e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523353e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.56315e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529406e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.532169e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547246e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.46224e-08, 6.465288e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532766e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472856e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.35757e-08, -6.385525e-08, -6.38009e-08, -6.402639e-08, -6.39013e-08, 
    -6.404895e-08, -6.363237e-08, -6.386636e-08, -6.371698e-08, 
    -6.360087e-08, -6.446398e-08, -6.403645e-08, -6.490803e-08, 
    -6.463537e-08, -6.532027e-08, -6.48656e-08, -6.541195e-08, -6.530715e-08, 
    -6.562256e-08, -6.55322e-08, -6.593564e-08, -6.566426e-08, -6.614476e-08, 
    -6.587083e-08, -6.591368e-08, -6.565531e-08, -6.412248e-08, 
    -6.441075e-08, -6.41054e-08, -6.41465e-08, -6.412806e-08, -6.390389e-08, 
    -6.379093e-08, -6.355432e-08, -6.359728e-08, -6.377105e-08, 
    -6.416499e-08, -6.403126e-08, -6.436827e-08, -6.436066e-08, 
    -6.473585e-08, -6.456669e-08, -6.519728e-08, -6.501806e-08, 
    -6.553597e-08, -6.540572e-08, -6.552985e-08, -6.549221e-08, 
    -6.553034e-08, -6.533932e-08, -6.542116e-08, -6.525307e-08, 
    -6.459837e-08, -6.479079e-08, -6.421691e-08, -6.387185e-08, 
    -6.364264e-08, -6.347999e-08, -6.350298e-08, -6.354682e-08, 
    -6.377207e-08, -6.398385e-08, -6.414524e-08, -6.42532e-08, -6.435957e-08, 
    -6.468156e-08, -6.485197e-08, -6.523353e-08, -6.516466e-08, 
    -6.528133e-08, -6.539276e-08, -6.557987e-08, -6.554907e-08, -6.56315e-08, 
    -6.527824e-08, -6.551303e-08, -6.512544e-08, -6.523145e-08, 
    -6.438852e-08, -6.406734e-08, -6.393085e-08, -6.381136e-08, 
    -6.352067e-08, -6.372141e-08, -6.364228e-08, -6.383054e-08, 
    -6.395017e-08, -6.3891e-08, -6.425615e-08, -6.411419e-08, -6.486207e-08, 
    -6.453993e-08, -6.537977e-08, -6.51788e-08, -6.542793e-08, -6.53008e-08, 
    -6.551863e-08, -6.532259e-08, -6.566219e-08, -6.573613e-08, -6.56856e-08, 
    -6.587971e-08, -6.531172e-08, -6.552985e-08, -6.388935e-08, 
    -6.389899e-08, -6.394394e-08, -6.374634e-08, -6.373425e-08, 
    -6.355315e-08, -6.371429e-08, -6.378291e-08, -6.39571e-08, -6.406013e-08, 
    -6.415808e-08, -6.437342e-08, -6.461393e-08, -6.495023e-08, 
    -6.519183e-08, -6.535377e-08, -6.525447e-08, -6.534214e-08, 
    -6.524414e-08, -6.519819e-08, -6.570843e-08, -6.542193e-08, 
    -6.585179e-08, -6.5828e-08, -6.563347e-08, -6.583068e-08, -6.390577e-08, 
    -6.385024e-08, -6.365745e-08, -6.380832e-08, -6.353343e-08, -6.36873e-08, 
    -6.377579e-08, -6.411717e-08, -6.419216e-08, -6.426171e-08, 
    -6.439907e-08, -6.457535e-08, -6.488458e-08, -6.515364e-08, 
    -6.539925e-08, -6.538125e-08, -6.538759e-08, -6.544246e-08, 
    -6.530654e-08, -6.546477e-08, -6.549133e-08, -6.542189e-08, 
    -6.582482e-08, -6.570971e-08, -6.58275e-08, -6.575254e-08, -6.386828e-08, 
    -6.396172e-08, -6.391124e-08, -6.400618e-08, -6.393929e-08, 
    -6.423671e-08, -6.432588e-08, -6.474312e-08, -6.457188e-08, 
    -6.484441e-08, -6.459956e-08, -6.464295e-08, -6.485331e-08, 
    -6.461279e-08, -6.513881e-08, -6.47822e-08, -6.544459e-08, -6.508849e-08, 
    -6.546691e-08, -6.539818e-08, -6.551196e-08, -6.561386e-08, 
    -6.574206e-08, -6.59786e-08, -6.592382e-08, -6.612164e-08, -6.410102e-08, 
    -6.422221e-08, -6.421153e-08, -6.433836e-08, -6.443215e-08, 
    -6.463544e-08, -6.496149e-08, -6.483888e-08, -6.506396e-08, 
    -6.510916e-08, -6.476719e-08, -6.497716e-08, -6.430331e-08, 
    -6.441219e-08, -6.434736e-08, -6.411058e-08, -6.486714e-08, 
    -6.447888e-08, -6.519582e-08, -6.498549e-08, -6.559934e-08, 
    -6.529406e-08, -6.589367e-08, -6.615002e-08, -6.639124e-08, 
    -6.667317e-08, -6.428834e-08, -6.4206e-08, -6.435344e-08, -6.455743e-08, 
    -6.47467e-08, -6.499832e-08, -6.502406e-08, -6.507121e-08, -6.51933e-08, 
    -6.529596e-08, -6.508611e-08, -6.532169e-08, -6.443745e-08, 
    -6.490084e-08, -6.417487e-08, -6.439348e-08, -6.454541e-08, 
    -6.447876e-08, -6.482487e-08, -6.490644e-08, -6.523793e-08, 
    -6.506657e-08, -6.608675e-08, -6.56354e-08, -6.688783e-08, -6.653783e-08, 
    -6.417723e-08, -6.428806e-08, -6.467379e-08, -6.449026e-08, 
    -6.501512e-08, -6.514431e-08, -6.524932e-08, -6.538358e-08, 
    -6.539807e-08, -6.547761e-08, -6.534727e-08, -6.547246e-08, 
    -6.499886e-08, -6.52105e-08, -6.46297e-08, -6.477106e-08, -6.470603e-08, 
    -6.463469e-08, -6.485485e-08, -6.508942e-08, -6.509442e-08, 
    -6.516963e-08, -6.53816e-08, -6.501724e-08, -6.614502e-08, -6.544855e-08, 
    -6.440892e-08, -6.46224e-08, -6.465288e-08, -6.457019e-08, -6.513136e-08, 
    -6.492802e-08, -6.547567e-08, -6.532766e-08, -6.557018e-08, 
    -6.544967e-08, -6.543194e-08, -6.527716e-08, -6.51808e-08, -6.493735e-08, 
    -6.473926e-08, -6.458218e-08, -6.46187e-08, -6.479126e-08, -6.510376e-08, 
    -6.539939e-08, -6.533463e-08, -6.555175e-08, -6.497706e-08, 
    -6.521804e-08, -6.512491e-08, -6.536776e-08, -6.483562e-08, 
    -6.528879e-08, -6.471979e-08, -6.476968e-08, -6.492399e-08, -6.52344e-08, 
    -6.530306e-08, -6.537638e-08, -6.533113e-08, -6.51117e-08, -6.507574e-08, 
    -6.492024e-08, -6.487731e-08, -6.475882e-08, -6.466072e-08, 
    -6.475035e-08, -6.484448e-08, -6.511178e-08, -6.535268e-08, 
    -6.561532e-08, -6.567959e-08, -6.598647e-08, -6.573666e-08, -6.61489e-08, 
    -6.579844e-08, -6.64051e-08, -6.531504e-08, -6.578811e-08, -6.493101e-08, 
    -6.502334e-08, -6.519036e-08, -6.557342e-08, -6.536661e-08, 
    -6.560847e-08, -6.507433e-08, -6.479721e-08, -6.47255e-08, -6.459173e-08, 
    -6.472856e-08, -6.471743e-08, -6.484837e-08, -6.480629e-08, 
    -6.512066e-08, -6.49518e-08, -6.54315e-08, -6.560656e-08, -6.610091e-08, 
    -6.640397e-08, -6.671245e-08, -6.684864e-08, -6.689009e-08, -6.690742e-08 ;

 NET_NMIN =
  8.956404e-09, 8.995784e-09, 8.988128e-09, 9.019892e-09, 9.002271e-09, 
    9.02307e-09, 8.964387e-09, 8.997348e-09, 8.976306e-09, 8.959948e-09, 
    9.081533e-09, 9.021308e-09, 9.144085e-09, 9.105677e-09, 9.202157e-09, 
    9.138109e-09, 9.215071e-09, 9.200308e-09, 9.244739e-09, 9.23201e-09, 
    9.288842e-09, 9.250614e-09, 9.3183e-09, 9.279711e-09, 9.285748e-09, 
    9.249352e-09, 9.033427e-09, 9.074036e-09, 9.031021e-09, 9.036812e-09, 
    9.034213e-09, 9.002636e-09, 8.986722e-09, 8.953393e-09, 8.959444e-09, 
    8.983923e-09, 9.039416e-09, 9.020578e-09, 9.068052e-09, 9.06698e-09, 
    9.119832e-09, 9.096002e-09, 9.184832e-09, 9.159585e-09, 9.232542e-09, 
    9.214194e-09, 9.231679e-09, 9.226378e-09, 9.231749e-09, 9.20484e-09, 
    9.216369e-09, 9.192691e-09, 9.100465e-09, 9.127571e-09, 9.04673e-09, 
    8.998122e-09, 8.965833e-09, 8.942921e-09, 8.94616e-09, 8.952335e-09, 
    8.984067e-09, 9.013899e-09, 9.036634e-09, 9.051842e-09, 9.066826e-09, 
    9.112184e-09, 9.136189e-09, 9.189939e-09, 9.180237e-09, 9.196671e-09, 
    9.212369e-09, 9.238725e-09, 9.234387e-09, 9.246e-09, 9.196237e-09, 
    9.22931e-09, 9.174712e-09, 9.189645e-09, 9.070903e-09, 9.02566e-09, 
    9.006433e-09, 8.9896e-09, 8.948651e-09, 8.976929e-09, 8.965782e-09, 
    8.992302e-09, 9.009154e-09, 9.000819e-09, 9.052258e-09, 9.032259e-09, 
    9.137612e-09, 9.092234e-09, 9.210538e-09, 9.182228e-09, 9.217323e-09, 
    9.199415e-09, 9.2301e-09, 9.202483e-09, 9.250321e-09, 9.260738e-09, 
    9.253619e-09, 9.280963e-09, 9.200953e-09, 9.23168e-09, 9.000586e-09, 
    9.001945e-09, 9.008278e-09, 8.980441e-09, 8.978739e-09, 8.953227e-09, 
    8.975927e-09, 8.985593e-09, 9.01013e-09, 9.024645e-09, 9.038442e-09, 
    9.068778e-09, 9.102657e-09, 9.15003e-09, 9.184063e-09, 9.206877e-09, 
    9.192887e-09, 9.205238e-09, 9.191432e-09, 9.18496e-09, 9.256835e-09, 
    9.216477e-09, 9.27703e-09, 9.27368e-09, 9.246276e-09, 9.274057e-09, 
    9.0029e-09, 8.995078e-09, 8.967919e-09, 8.989173e-09, 8.950449e-09, 
    8.972125e-09, 8.984589e-09, 9.032679e-09, 9.043243e-09, 9.053041e-09, 
    9.07239e-09, 9.097222e-09, 9.140783e-09, 9.178684e-09, 9.213282e-09, 
    9.210747e-09, 9.211639e-09, 9.219368e-09, 9.200223e-09, 9.222512e-09, 
    9.226253e-09, 9.216472e-09, 9.27323e-09, 9.257015e-09, 9.273608e-09, 
    9.26305e-09, 8.99762e-09, 9.010782e-09, 9.00367e-09, 9.017044e-09, 
    9.007622e-09, 9.049519e-09, 9.06208e-09, 9.120856e-09, 9.096733e-09, 
    9.135123e-09, 9.100632e-09, 9.106745e-09, 9.136377e-09, 9.102497e-09, 
    9.176595e-09, 9.12636e-09, 9.219669e-09, 9.169507e-09, 9.222813e-09, 
    9.213132e-09, 9.22916e-09, 9.243514e-09, 9.261572e-09, 9.294893e-09, 
    9.287177e-09, 9.315042e-09, 9.030404e-09, 9.047476e-09, 9.045972e-09, 
    9.063838e-09, 9.07705e-09, 9.105687e-09, 9.151616e-09, 9.134345e-09, 
    9.166052e-09, 9.172417e-09, 9.124246e-09, 9.153823e-09, 9.058901e-09, 
    9.074238e-09, 9.065106e-09, 9.03175e-09, 9.138326e-09, 9.083633e-09, 
    9.184626e-09, 9.154998e-09, 9.241467e-09, 9.198465e-09, 9.28293e-09, 
    9.31904e-09, 9.35302e-09, 9.392735e-09, 9.056793e-09, 9.045192e-09, 
    9.065962e-09, 9.094698e-09, 9.12136e-09, 9.156805e-09, 9.160431e-09, 
    9.167072e-09, 9.184271e-09, 9.198732e-09, 9.169172e-09, 9.202358e-09, 
    9.077796e-09, 9.143073e-09, 9.040807e-09, 9.071603e-09, 9.093005e-09, 
    9.083616e-09, 9.13237e-09, 9.143862e-09, 9.190557e-09, 9.166418e-09, 
    9.310128e-09, 9.246548e-09, 9.422972e-09, 9.37367e-09, 9.041139e-09, 
    9.056752e-09, 9.11109e-09, 9.085236e-09, 9.15917e-09, 9.177369e-09, 
    9.192163e-09, 9.211075e-09, 9.213116e-09, 9.224322e-09, 9.20596e-09, 
    9.223596e-09, 9.156881e-09, 9.186694e-09, 9.104878e-09, 9.124792e-09, 
    9.11563e-09, 9.105581e-09, 9.136595e-09, 9.169637e-09, 9.170342e-09, 
    9.180937e-09, 9.210796e-09, 9.15947e-09, 9.318336e-09, 9.220227e-09, 
    9.073776e-09, 9.10385e-09, 9.108144e-09, 9.096495e-09, 9.175545e-09, 
    9.146903e-09, 9.224048e-09, 9.203198e-09, 9.23736e-09, 9.220384e-09, 
    9.217888e-09, 9.196084e-09, 9.18251e-09, 9.148216e-09, 9.120313e-09, 
    9.098184e-09, 9.10333e-09, 9.127636e-09, 9.171658e-09, 9.213302e-09, 
    9.20418e-09, 9.234764e-09, 9.15381e-09, 9.187756e-09, 9.174636e-09, 
    9.208845e-09, 9.133886e-09, 9.197723e-09, 9.117569e-09, 9.124596e-09, 
    9.146334e-09, 9.190059e-09, 9.199732e-09, 9.210061e-09, 9.203687e-09, 
    9.172775e-09, 9.167711e-09, 9.145806e-09, 9.139758e-09, 9.123067e-09, 
    9.109248e-09, 9.121874e-09, 9.135134e-09, 9.172788e-09, 9.206722e-09, 
    9.243719e-09, 9.252772e-09, 9.296001e-09, 9.260813e-09, 9.318883e-09, 
    9.269515e-09, 9.354972e-09, 9.201419e-09, 9.268061e-09, 9.147323e-09, 
    9.16033e-09, 9.183857e-09, 9.237817e-09, 9.208684e-09, 9.242754e-09, 
    9.167512e-09, 9.128476e-09, 9.118374e-09, 9.09953e-09, 9.118805e-09, 
    9.117237e-09, 9.135682e-09, 9.129755e-09, 9.174038e-09, 9.150251e-09, 
    9.217825e-09, 9.242485e-09, 9.312123e-09, 9.354813e-09, 9.398266e-09, 
    9.417451e-09, 9.42329e-09, 9.425731e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14 ;

 O_SCALAR =
  0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8 ;

 PCH4 =
  0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993 ;

 PCO2 =
  29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  4.490659e-14, 4.502776e-14, 4.500422e-14, 4.510186e-14, 4.504772e-14, 
    4.511163e-14, 4.493118e-14, 4.503255e-14, 4.496786e-14, 4.491752e-14, 
    4.529107e-14, 4.510622e-14, 4.548291e-14, 4.536523e-14, 4.566065e-14, 
    4.546458e-14, 4.570015e-14, 4.565504e-14, 4.579087e-14, 4.575198e-14, 
    4.592545e-14, 4.580882e-14, 4.601533e-14, 4.589763e-14, 4.591603e-14, 
    4.580496e-14, 4.514348e-14, 4.526806e-14, 4.513609e-14, 4.515386e-14, 
    4.51459e-14, 4.504883e-14, 4.499986e-14, 4.489735e-14, 4.491597e-14, 
    4.499127e-14, 4.516186e-14, 4.510401e-14, 4.524983e-14, 4.524654e-14, 
    4.540864e-14, 4.533558e-14, 4.560769e-14, 4.553044e-14, 4.57536e-14, 
    4.569751e-14, 4.575096e-14, 4.573476e-14, 4.575117e-14, 4.56689e-14, 
    4.570415e-14, 4.563174e-14, 4.534926e-14, 4.543234e-14, 4.518434e-14, 
    4.503489e-14, 4.493562e-14, 4.48651e-14, 4.487507e-14, 4.489407e-14, 
    4.499171e-14, 4.508348e-14, 4.515334e-14, 4.520005e-14, 4.524606e-14, 
    4.538511e-14, 4.545872e-14, 4.562329e-14, 4.559364e-14, 4.564389e-14, 
    4.569193e-14, 4.577248e-14, 4.575923e-14, 4.57947e-14, 4.564259e-14, 
    4.57437e-14, 4.557676e-14, 4.562242e-14, 4.525843e-14, 4.511962e-14, 
    4.506046e-14, 4.500874e-14, 4.488274e-14, 4.496976e-14, 4.493546e-14, 
    4.501708e-14, 4.506889e-14, 4.504327e-14, 4.520133e-14, 4.51399e-14, 
    4.546308e-14, 4.532399e-14, 4.568633e-14, 4.559973e-14, 4.570708e-14, 
    4.565232e-14, 4.574612e-14, 4.56617e-14, 4.580791e-14, 4.583971e-14, 
    4.581798e-14, 4.590147e-14, 4.565702e-14, 4.575095e-14, 4.504255e-14, 
    4.504672e-14, 4.50662e-14, 4.498056e-14, 4.497533e-14, 4.489683e-14, 
    4.496669e-14, 4.499642e-14, 4.50719e-14, 4.51165e-14, 4.515889e-14, 
    4.525204e-14, 4.535595e-14, 4.550115e-14, 4.560534e-14, 4.567514e-14, 
    4.563236e-14, 4.567013e-14, 4.56279e-14, 4.56081e-14, 4.582779e-14, 
    4.570447e-14, 4.588947e-14, 4.587924e-14, 4.579554e-14, 4.58804e-14, 
    4.504966e-14, 4.502562e-14, 4.494205e-14, 4.500745e-14, 4.488828e-14, 
    4.495499e-14, 4.499331e-14, 4.514116e-14, 4.517365e-14, 4.520372e-14, 
    4.526313e-14, 4.533932e-14, 4.547282e-14, 4.558886e-14, 4.569473e-14, 
    4.568698e-14, 4.56897e-14, 4.571333e-14, 4.565478e-14, 4.572294e-14, 
    4.573436e-14, 4.570447e-14, 4.587787e-14, 4.582837e-14, 4.587902e-14, 
    4.58468e-14, 4.503343e-14, 4.50739e-14, 4.505203e-14, 4.509313e-14, 
    4.506417e-14, 4.519288e-14, 4.523144e-14, 4.541174e-14, 4.533781e-14, 
    4.545548e-14, 4.534978e-14, 4.536851e-14, 4.545926e-14, 4.53555e-14, 
    4.558244e-14, 4.542859e-14, 4.571425e-14, 4.556073e-14, 4.572385e-14, 
    4.569427e-14, 4.574327e-14, 4.578711e-14, 4.584228e-14, 4.594395e-14, 
    4.592042e-14, 4.600542e-14, 4.51342e-14, 4.518662e-14, 4.518203e-14, 
    4.523688e-14, 4.527743e-14, 4.536528e-14, 4.550603e-14, 4.545313e-14, 
    4.555025e-14, 4.556973e-14, 4.542219e-14, 4.551277e-14, 4.522171e-14, 
    4.526876e-14, 4.524076e-14, 4.513832e-14, 4.546528e-14, 4.529759e-14, 
    4.560706e-14, 4.551639e-14, 4.578086e-14, 4.564937e-14, 4.590746e-14, 
    4.601754e-14, 4.612116e-14, 4.624198e-14, 4.521525e-14, 4.517964e-14, 
    4.524341e-14, 4.533154e-14, 4.541332e-14, 4.552192e-14, 4.553304e-14, 
    4.555336e-14, 4.560599e-14, 4.565023e-14, 4.555976e-14, 4.566132e-14, 
    4.527962e-14, 4.547984e-14, 4.516615e-14, 4.526067e-14, 4.532636e-14, 
    4.529757e-14, 4.544709e-14, 4.548229e-14, 4.562519e-14, 4.555137e-14, 
    4.599036e-14, 4.579634e-14, 4.633398e-14, 4.618398e-14, 4.516718e-14, 
    4.521514e-14, 4.538182e-14, 4.530255e-14, 4.552917e-14, 4.558485e-14, 
    4.563014e-14, 4.568796e-14, 4.569422e-14, 4.572846e-14, 4.567234e-14, 
    4.572626e-14, 4.552215e-14, 4.56134e-14, 4.536281e-14, 4.542384e-14, 
    4.539578e-14, 4.536497e-14, 4.546003e-14, 4.556118e-14, 4.556338e-14, 
    4.559576e-14, 4.568695e-14, 4.553009e-14, 4.60153e-14, 4.571581e-14, 
    4.52674e-14, 4.53596e-14, 4.537281e-14, 4.53371e-14, 4.557929e-14, 
    4.549159e-14, 4.572763e-14, 4.566389e-14, 4.576832e-14, 4.571644e-14, 
    4.57088e-14, 4.564213e-14, 4.560059e-14, 4.549561e-14, 4.541011e-14, 
    4.534228e-14, 4.535806e-14, 4.543255e-14, 4.556737e-14, 4.569476e-14, 
    4.566686e-14, 4.576039e-14, 4.551275e-14, 4.561662e-14, 4.557649e-14, 
    4.568115e-14, 4.545171e-14, 4.5647e-14, 4.540172e-14, 4.542326e-14, 
    4.548985e-14, 4.562364e-14, 4.565328e-14, 4.568485e-14, 4.566539e-14, 
    4.55708e-14, 4.555531e-14, 4.548824e-14, 4.54697e-14, 4.541857e-14, 
    4.537621e-14, 4.54149e-14, 4.545552e-14, 4.557085e-14, 4.567464e-14, 
    4.578773e-14, 4.581541e-14, 4.594725e-14, 4.583988e-14, 4.601695e-14, 
    4.586634e-14, 4.612697e-14, 4.565836e-14, 4.586199e-14, 4.549289e-14, 
    4.553273e-14, 4.560467e-14, 4.576966e-14, 4.568066e-14, 4.578475e-14, 
    4.555471e-14, 4.54351e-14, 4.540418e-14, 4.53464e-14, 4.540551e-14, 
    4.54007e-14, 4.545723e-14, 4.543907e-14, 4.557468e-14, 4.550186e-14, 
    4.570859e-14, 4.578394e-14, 4.59965e-14, 4.612657e-14, 4.625888e-14, 
    4.631722e-14, 4.633497e-14, 4.634239e-14 ;

 POT_F_DENIT =
  1.021992e-12, 1.024837e-12, 1.024282e-12, 1.026577e-12, 1.025303e-12, 
    1.026805e-12, 1.022566e-12, 1.024947e-12, 1.023426e-12, 1.022243e-12, 
    1.031025e-12, 1.026675e-12, 1.035534e-12, 1.032762e-12, 1.039719e-12, 
    1.035103e-12, 1.040649e-12, 1.039584e-12, 1.042784e-12, 1.041867e-12, 
    1.045961e-12, 1.043206e-12, 1.04808e-12, 1.045302e-12, 1.045736e-12, 
    1.043113e-12, 1.027553e-12, 1.030487e-12, 1.027378e-12, 1.027797e-12, 
    1.027608e-12, 1.025328e-12, 1.024179e-12, 1.021769e-12, 1.022206e-12, 
    1.023975e-12, 1.027981e-12, 1.02662e-12, 1.030046e-12, 1.029968e-12, 
    1.033781e-12, 1.032062e-12, 1.038468e-12, 1.036646e-12, 1.041904e-12, 
    1.040582e-12, 1.041842e-12, 1.041458e-12, 1.041845e-12, 1.039906e-12, 
    1.040736e-12, 1.03903e-12, 1.03239e-12, 1.034345e-12, 1.028512e-12, 
    1.025003e-12, 1.022668e-12, 1.021013e-12, 1.021246e-12, 1.021693e-12, 
    1.023984e-12, 1.026137e-12, 1.027778e-12, 1.028875e-12, 1.029956e-12, 
    1.033231e-12, 1.034961e-12, 1.038835e-12, 1.038135e-12, 1.039319e-12, 
    1.04045e-12, 1.042348e-12, 1.042035e-12, 1.042871e-12, 1.039284e-12, 
    1.041668e-12, 1.037732e-12, 1.038809e-12, 1.030259e-12, 1.026989e-12, 
    1.025602e-12, 1.024385e-12, 1.021426e-12, 1.023469e-12, 1.022663e-12, 
    1.024577e-12, 1.025794e-12, 1.025191e-12, 1.028905e-12, 1.02746e-12, 
    1.035063e-12, 1.031789e-12, 1.040318e-12, 1.038277e-12, 1.040806e-12, 
    1.039515e-12, 1.041726e-12, 1.039735e-12, 1.043181e-12, 1.043932e-12, 
    1.043418e-12, 1.045387e-12, 1.039622e-12, 1.041837e-12, 1.025177e-12, 
    1.025276e-12, 1.025732e-12, 1.023722e-12, 1.023599e-12, 1.021755e-12, 
    1.023394e-12, 1.024092e-12, 1.025863e-12, 1.02691e-12, 1.027906e-12, 
    1.030095e-12, 1.03254e-12, 1.035956e-12, 1.038409e-12, 1.040052e-12, 
    1.039044e-12, 1.039933e-12, 1.038938e-12, 1.03847e-12, 1.04365e-12, 
    1.040742e-12, 1.045102e-12, 1.044861e-12, 1.042887e-12, 1.044887e-12, 
    1.025344e-12, 1.024778e-12, 1.022816e-12, 1.02435e-12, 1.021553e-12, 
    1.023119e-12, 1.024019e-12, 1.027491e-12, 1.028252e-12, 1.028959e-12, 
    1.030355e-12, 1.032146e-12, 1.035289e-12, 1.03802e-12, 1.040513e-12, 
    1.04033e-12, 1.040394e-12, 1.04095e-12, 1.03957e-12, 1.041176e-12, 
    1.041445e-12, 1.04074e-12, 1.044827e-12, 1.04366e-12, 1.044854e-12, 
    1.044093e-12, 1.024961e-12, 1.025911e-12, 1.025396e-12, 1.026362e-12, 
    1.025681e-12, 1.028707e-12, 1.029613e-12, 1.033853e-12, 1.032111e-12, 
    1.034881e-12, 1.032391e-12, 1.032832e-12, 1.034971e-12, 1.032524e-12, 
    1.037869e-12, 1.034246e-12, 1.040971e-12, 1.037357e-12, 1.041197e-12, 
    1.040498e-12, 1.041652e-12, 1.042687e-12, 1.043986e-12, 1.046387e-12, 
    1.04583e-12, 1.047836e-12, 1.027327e-12, 1.028559e-12, 1.028449e-12, 
    1.029738e-12, 1.030691e-12, 1.032757e-12, 1.03607e-12, 1.034823e-12, 
    1.037109e-12, 1.037568e-12, 1.034093e-12, 1.036227e-12, 1.029378e-12, 
    1.030485e-12, 1.029825e-12, 1.027417e-12, 1.035107e-12, 1.031161e-12, 
    1.038444e-12, 1.036307e-12, 1.042538e-12, 1.03944e-12, 1.045523e-12, 
    1.048125e-12, 1.050567e-12, 1.053425e-12, 1.02923e-12, 1.028392e-12, 
    1.02989e-12, 1.031965e-12, 1.033887e-12, 1.036443e-12, 1.036703e-12, 
    1.037182e-12, 1.038421e-12, 1.039463e-12, 1.037333e-12, 1.039723e-12, 
    1.030743e-12, 1.035449e-12, 1.028069e-12, 1.030293e-12, 1.031836e-12, 
    1.031158e-12, 1.034674e-12, 1.035502e-12, 1.038869e-12, 1.037128e-12, 
    1.047482e-12, 1.042903e-12, 1.055596e-12, 1.052052e-12, 1.028099e-12, 
    1.029225e-12, 1.033146e-12, 1.03128e-12, 1.036612e-12, 1.037924e-12, 
    1.038989e-12, 1.040353e-12, 1.040498e-12, 1.041306e-12, 1.039982e-12, 
    1.041253e-12, 1.036443e-12, 1.038592e-12, 1.032691e-12, 1.034128e-12, 
    1.033466e-12, 1.03274e-12, 1.034977e-12, 1.037361e-12, 1.03741e-12, 
    1.038173e-12, 1.040329e-12, 1.036624e-12, 1.048073e-12, 1.041006e-12, 
    1.030453e-12, 1.032624e-12, 1.032932e-12, 1.032091e-12, 1.037791e-12, 
    1.035726e-12, 1.041286e-12, 1.039783e-12, 1.042244e-12, 1.041021e-12, 
    1.04084e-12, 1.039269e-12, 1.038289e-12, 1.035817e-12, 1.033803e-12, 
    1.032207e-12, 1.032577e-12, 1.034331e-12, 1.037505e-12, 1.040506e-12, 
    1.039848e-12, 1.04205e-12, 1.036215e-12, 1.038663e-12, 1.037716e-12, 
    1.040182e-12, 1.034788e-12, 1.039394e-12, 1.03361e-12, 1.034116e-12, 
    1.035684e-12, 1.038838e-12, 1.039532e-12, 1.040277e-12, 1.039816e-12, 
    1.037589e-12, 1.037223e-12, 1.035642e-12, 1.035206e-12, 1.034001e-12, 
    1.033003e-12, 1.033915e-12, 1.03487e-12, 1.037585e-12, 1.040031e-12, 
    1.042696e-12, 1.043347e-12, 1.046462e-12, 1.043927e-12, 1.04811e-12, 
    1.044556e-12, 1.050705e-12, 1.039658e-12, 1.044459e-12, 1.035755e-12, 
    1.036692e-12, 1.038389e-12, 1.042277e-12, 1.040176e-12, 1.042632e-12, 
    1.037208e-12, 1.034393e-12, 1.033663e-12, 1.032303e-12, 1.033693e-12, 
    1.03358e-12, 1.034909e-12, 1.034481e-12, 1.037674e-12, 1.035959e-12, 
    1.040829e-12, 1.042606e-12, 1.04762e-12, 1.050692e-12, 1.053816e-12, 
    1.055194e-12, 1.055614e-12, 1.055789e-12 ;

 POT_F_NIT =
  4.014551e-11, 4.049193e-11, 4.042445e-11, 4.070474e-11, 4.054912e-11, 
    4.073283e-11, 4.021559e-11, 4.050569e-11, 4.032037e-11, 4.017659e-11, 
    4.125151e-11, 4.071723e-11, 4.181026e-11, 4.146671e-11, 4.233246e-11, 
    4.17567e-11, 4.244905e-11, 4.231578e-11, 4.27175e-11, 4.260221e-11, 
    4.31182e-11, 4.277076e-11, 4.338693e-11, 4.303508e-11, 4.309002e-11, 
    4.27593e-11, 4.082448e-11, 4.118483e-11, 4.080318e-11, 4.085445e-11, 
    4.083144e-11, 4.055232e-11, 4.041205e-11, 4.011905e-11, 4.017215e-11, 
    4.038738e-11, 4.087749e-11, 4.071076e-11, 4.113158e-11, 4.112206e-11, 
    4.159313e-11, 4.138039e-11, 4.21763e-11, 4.194928e-11, 4.260701e-11, 
    4.24411e-11, 4.25992e-11, 4.255122e-11, 4.259982e-11, 4.235663e-11, 
    4.246073e-11, 4.224705e-11, 4.142024e-11, 4.166238e-11, 4.094233e-11, 
    4.05125e-11, 4.022828e-11, 4.002723e-11, 4.005561e-11, 4.010976e-11, 
    4.038864e-11, 4.065173e-11, 4.085283e-11, 4.098763e-11, 4.112067e-11, 
    4.152479e-11, 4.173948e-11, 4.222228e-11, 4.213492e-11, 4.228295e-11, 
    4.24246e-11, 4.266299e-11, 4.26237e-11, 4.272889e-11, 4.227901e-11, 
    4.257773e-11, 4.208518e-11, 4.22196e-11, 4.115696e-11, 4.075572e-11, 
    4.058582e-11, 4.043738e-11, 4.007744e-11, 4.032583e-11, 4.022781e-11, 
    4.046117e-11, 4.060982e-11, 4.053626e-11, 4.099131e-11, 4.081408e-11, 
    4.175221e-11, 4.134678e-11, 4.240807e-11, 4.215283e-11, 4.246935e-11, 
    4.230769e-11, 4.258488e-11, 4.233536e-11, 4.276807e-11, 4.28626e-11, 
    4.279798e-11, 4.304643e-11, 4.232152e-11, 4.259916e-11, 4.053422e-11, 
    4.054622e-11, 4.06021e-11, 4.035672e-11, 4.034173e-11, 4.011757e-11, 
    4.031698e-11, 4.040206e-11, 4.061843e-11, 4.07467e-11, 4.086882e-11, 
    4.113801e-11, 4.143972e-11, 4.186351e-11, 4.216935e-11, 4.2375e-11, 
    4.224883e-11, 4.236021e-11, 4.22357e-11, 4.217741e-11, 4.282716e-11, 
    4.246168e-11, 4.301064e-11, 4.298017e-11, 4.273137e-11, 4.298359e-11, 
    4.055463e-11, 4.048563e-11, 4.024659e-11, 4.043359e-11, 4.009319e-11, 
    4.028355e-11, 4.039321e-11, 4.081778e-11, 4.091136e-11, 4.099825e-11, 
    4.117012e-11, 4.139123e-11, 4.178061e-11, 4.212092e-11, 4.243283e-11, 
    4.240993e-11, 4.241799e-11, 4.248782e-11, 4.231495e-11, 4.251622e-11, 
    4.255005e-11, 4.246162e-11, 4.297608e-11, 4.282877e-11, 4.297951e-11, 
    4.288355e-11, 4.050804e-11, 4.062419e-11, 4.05614e-11, 4.06795e-11, 
    4.059628e-11, 4.096701e-11, 4.10785e-11, 4.160226e-11, 4.138687e-11, 
    4.172991e-11, 4.142164e-11, 4.147618e-11, 4.174113e-11, 4.143826e-11, 
    4.210211e-11, 4.165145e-11, 4.249052e-11, 4.203836e-11, 4.251894e-11, 
    4.243145e-11, 4.257633e-11, 4.270632e-11, 4.287013e-11, 4.317326e-11, 
    4.310296e-11, 4.33571e-11, 4.079765e-11, 4.094889e-11, 4.093556e-11, 
    4.10941e-11, 4.121157e-11, 4.146675e-11, 4.187774e-11, 4.172293e-11, 
    4.200734e-11, 4.206455e-11, 4.163255e-11, 4.189752e-11, 4.105023e-11, 
    4.118651e-11, 4.110533e-11, 4.080952e-11, 4.175855e-11, 4.127009e-11, 
    4.217436e-11, 4.190802e-11, 4.268777e-11, 4.229906e-11, 4.306429e-11, 
    4.339361e-11, 4.370469e-11, 4.406973e-11, 4.103155e-11, 4.092864e-11, 
    4.111297e-11, 4.136873e-11, 4.160675e-11, 4.192429e-11, 4.195684e-11, 
    4.201649e-11, 4.217119e-11, 4.230151e-11, 4.203536e-11, 4.23342e-11, 
    4.121816e-11, 4.180109e-11, 4.088972e-11, 4.116307e-11, 4.135357e-11, 
    4.126994e-11, 4.170521e-11, 4.180813e-11, 4.222776e-11, 4.201057e-11, 
    4.33122e-11, 4.273379e-11, 4.434871e-11, 4.389429e-11, 4.089271e-11, 
    4.103117e-11, 4.151497e-11, 4.128441e-11, 4.194552e-11, 4.210908e-11, 
    4.224228e-11, 4.241289e-11, 4.243132e-11, 4.253259e-11, 4.236669e-11, 
    4.252602e-11, 4.192493e-11, 4.219299e-11, 4.145947e-11, 4.163739e-11, 
    4.155548e-11, 4.146574e-11, 4.174302e-11, 4.20395e-11, 4.204583e-11, 
    4.214112e-11, 4.24103e-11, 4.194813e-11, 4.338715e-11, 4.24955e-11, 
    4.118243e-11, 4.145034e-11, 4.148866e-11, 4.138473e-11, 4.209266e-11, 
    4.183543e-11, 4.253012e-11, 4.234177e-11, 4.265058e-11, 4.249698e-11, 
    4.24744e-11, 4.22776e-11, 4.215531e-11, 4.184718e-11, 4.159732e-11, 
    4.139974e-11, 4.144563e-11, 4.166282e-11, 4.205765e-11, 4.243294e-11, 
    4.235058e-11, 4.262701e-11, 4.189732e-11, 4.22025e-11, 4.208441e-11, 
    4.239267e-11, 4.171881e-11, 4.22924e-11, 4.157284e-11, 4.163567e-11, 
    4.183032e-11, 4.222332e-11, 4.231049e-11, 4.240371e-11, 4.234616e-11, 
    4.206773e-11, 4.202219e-11, 4.182556e-11, 4.177135e-11, 4.162195e-11, 
    4.149846e-11, 4.161127e-11, 4.172991e-11, 4.206781e-11, 4.237352e-11, 
    4.270813e-11, 4.279021e-11, 4.318331e-11, 4.286318e-11, 4.339213e-11, 
    4.294223e-11, 4.372255e-11, 4.232573e-11, 4.29291e-11, 4.183919e-11, 
    4.19559e-11, 4.216745e-11, 4.26547e-11, 4.239127e-11, 4.269943e-11, 
    4.20204e-11, 4.167033e-11, 4.157999e-11, 4.141174e-11, 4.158383e-11, 
    4.156982e-11, 4.173482e-11, 4.168175e-11, 4.207904e-11, 4.186539e-11, 
    4.247378e-11, 4.269693e-11, 4.333038e-11, 4.372109e-11, 4.412066e-11, 
    4.429766e-11, 4.435161e-11, 4.437416e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.001208389, 0.001208317, 0.001208331, 0.001208274, 0.001208305, 
    0.001208268, 0.001208373, 0.001208315, 0.001208352, 0.001208381, 
    0.001208166, 0.001208271, 0.00120805, 0.001208118, 0.001207944, 
    0.001208062, 0.00120792, 0.001207946, 0.001207866, 0.001207888, 
    0.001207789, 0.001207855, 0.001207735, 0.001207804, 0.001207793, 
    0.001207857, 0.001208249, 0.001208179, 0.001208253, 0.001208243, 
    0.001208247, 0.001208305, 0.001208335, 0.001208393, 0.001208382, 
    0.001208339, 0.001208239, 0.001208272, 0.001208186, 0.001208187, 
    0.001208093, 0.001208135, 0.001207974, 0.001208021, 0.001207887, 
    0.001207921, 0.001207889, 0.001207899, 0.001207889, 0.001207938, 
    0.001207917, 0.001207959, 0.001208128, 0.001208079, 0.001208225, 
    0.001208315, 0.001208371, 0.001208412, 0.001208406, 0.001208396, 
    0.001208339, 0.001208284, 0.001208242, 0.001208215, 0.001208188, 
    0.001208109, 0.001208064, 0.001207965, 0.001207982, 0.001207953, 
    0.001207924, 0.001207877, 0.001207884, 0.001207864, 0.001207953, 
    0.001207894, 0.001207993, 0.001207965, 0.001208185, 0.001208263, 
    0.001208299, 0.001208328, 0.001208402, 0.001208351, 0.001208371, 
    0.001208323, 0.001208292, 0.001208307, 0.001208214, 0.001208251, 
    0.001208062, 0.001208143, 0.001207927, 0.001207978, 0.001207915, 
    0.001207947, 0.001207892, 0.001207942, 0.001207856, 0.001207838, 
    0.00120785, 0.001207801, 0.001207944, 0.00120789, 0.001208308, 
    0.001208305, 0.001208294, 0.001208345, 0.001208348, 0.001208394, 
    0.001208353, 0.001208336, 0.00120829, 0.001208264, 0.001208239, 
    0.001208185, 0.001208124, 0.001208039, 0.001207975, 0.001207934, 
    0.001207959, 0.001207937, 0.001207961, 0.001207973, 0.001207845, 
    0.001207917, 0.001207808, 0.001207814, 0.001207863, 0.001207813, 
    0.001208304, 0.001208318, 0.001208367, 0.001208328, 0.001208399, 
    0.00120836, 0.001208338, 0.001208251, 0.001208231, 0.001208213, 
    0.001208178, 0.001208133, 0.001208055, 0.001207985, 0.001207922, 
    0.001207927, 0.001207925, 0.001207911, 0.001207946, 0.001207906, 
    0.001207899, 0.001207917, 0.001207814, 0.001207844, 0.001207814, 
    0.001207833, 0.001208313, 0.001208289, 0.001208302, 0.001208278, 
    0.001208295, 0.001208221, 0.001208198, 0.001208092, 0.001208134, 
    0.001208066, 0.001208127, 0.001208117, 0.001208065, 0.001208124, 
    0.00120799, 0.001208083, 0.001207911, 0.001208005, 0.001207905, 
    0.001207922, 0.001207893, 0.001207868, 0.001207835, 0.001207776, 
    0.00120779, 0.00120774, 0.001208254, 0.001208224, 0.001208225, 
    0.001208193, 0.00120817, 0.001208118, 0.001208035, 0.001208066, 
    0.001208009, 0.001207998, 0.001208084, 0.001208032, 0.001208203, 
    0.001208176, 0.001208191, 0.001208252, 0.00120806, 0.001208159, 
    0.001207974, 0.001208029, 0.001207872, 0.00120795, 0.001207797, 
    0.001207735, 0.001207671, 0.001207602, 0.001208206, 0.001208227, 
    0.001208189, 0.001208139, 0.00120809, 0.001208026, 0.001208019, 
    0.001208007, 0.001207974, 0.001207948, 0.001208004, 0.001207942, 
    0.001208172, 0.001208051, 0.001208235, 0.001208181, 0.001208142, 
    0.001208158, 0.001208069, 0.001208049, 0.001207964, 0.001208008, 
    0.001207751, 0.001207864, 0.001207547, 0.001207636, 0.001208234, 
    0.001208206, 0.001208109, 0.001208155, 0.001208021, 0.001207987, 
    0.00120796, 0.001207927, 0.001207922, 0.001207903, 0.001207935, 
    0.001207904, 0.001208026, 0.00120797, 0.001208119, 0.001208084, 
    0.0012081, 0.001208118, 0.001208062, 0.001208004, 0.001208001, 
    0.001207981, 0.001207932, 0.001208021, 0.001207739, 0.001207914, 
    0.001208175, 0.001208123, 0.001208114, 0.001208134, 0.001207992, 
    0.001208044, 0.001207903, 0.00120794, 0.001207879, 0.001207909, 
    0.001207914, 0.001207953, 0.001207978, 0.001208042, 0.001208092, 
    0.001208131, 0.001208122, 0.001208079, 0.001208, 0.001207923, 
    0.001207939, 0.001207883, 0.001208031, 0.001207969, 0.001207994, 
    0.00120793, 0.001208067, 0.001207955, 0.001208096, 0.001208084, 
    0.001208045, 0.001207966, 0.001207947, 0.001207929, 0.001207939, 
    0.001207998, 0.001208006, 0.001208045, 0.001208057, 0.001208086, 
    0.001208111, 0.001208089, 0.001208065, 0.001207997, 0.001207935, 
    0.001207868, 0.001207851, 0.001207777, 0.001207839, 0.001207738, 
    0.001207827, 0.001207672, 0.001207946, 0.001207827, 0.001208042, 
    0.001208019, 0.001207977, 0.00120788, 0.001207931, 0.001207871, 
    0.001208007, 0.001208078, 0.001208095, 0.001208129, 0.001208094, 
    0.001208097, 0.001208063, 0.001208074, 0.001207995, 0.001208037, 
    0.001207915, 0.001207871, 0.001207746, 0.00120767, 0.00120759, 
    0.001207556, 0.001207546, 0.001207541 ;

 QBOT =
  0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_NODYNLNDUSE =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_R =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  3.259637e-06, 3.265722e-06, 3.264538e-06, 3.269444e-06, 3.266726e-06, 
    3.269934e-06, 3.26087e-06, 3.265963e-06, 3.262711e-06, 3.260185e-06, 
    3.278961e-06, 3.269663e-06, 3.288659e-06, 3.282704e-06, 3.298332e-06, 
    3.28773e-06, 3.300348e-06, 3.298046e-06, 3.304988e-06, 3.302998e-06, 
    3.311891e-06, 3.305907e-06, 3.316518e-06, 3.310462e-06, 3.311408e-06, 
    3.30571e-06, 3.271533e-06, 3.277802e-06, 3.271162e-06, 3.272055e-06, 
    3.271655e-06, 3.266782e-06, 3.264319e-06, 3.259174e-06, 3.260107e-06, 
    3.263887e-06, 3.272457e-06, 3.269551e-06, 3.276884e-06, 3.276718e-06, 
    3.284898e-06, 3.281206e-06, 3.295633e-06, 3.29107e-06, 3.303081e-06, 
    3.300214e-06, 3.302946e-06, 3.302117e-06, 3.302956e-06, 3.298753e-06, 
    3.300553e-06, 3.296858e-06, 3.281897e-06, 3.286098e-06, 3.273587e-06, 
    3.26608e-06, 3.261093e-06, 3.257558e-06, 3.258058e-06, 3.25901e-06, 
    3.263909e-06, 3.268522e-06, 3.272029e-06, 3.274378e-06, 3.276694e-06, 
    3.283708e-06, 3.287433e-06, 3.296428e-06, 3.294918e-06, 3.297477e-06, 
    3.299928e-06, 3.304047e-06, 3.303369e-06, 3.305184e-06, 3.297411e-06, 
    3.302574e-06, 3.293422e-06, 3.296384e-06, 3.277318e-06, 3.270335e-06, 
    3.267367e-06, 3.264765e-06, 3.258442e-06, 3.262807e-06, 3.261085e-06, 
    3.265185e-06, 3.26779e-06, 3.266502e-06, 3.274442e-06, 3.271354e-06, 
    3.287654e-06, 3.280622e-06, 3.299643e-06, 3.295228e-06, 3.300702e-06, 
    3.297907e-06, 3.302698e-06, 3.298386e-06, 3.305861e-06, 3.30749e-06, 
    3.306376e-06, 3.310661e-06, 3.298147e-06, 3.302945e-06, 3.266466e-06, 
    3.266676e-06, 3.267656e-06, 3.263349e-06, 3.263086e-06, 3.259148e-06, 
    3.262652e-06, 3.264146e-06, 3.267941e-06, 3.270178e-06, 3.272308e-06, 
    3.276995e-06, 3.282235e-06, 3.289583e-06, 3.295514e-06, 3.299072e-06, 
    3.29689e-06, 3.298816e-06, 3.296663e-06, 3.295654e-06, 3.306879e-06, 
    3.300569e-06, 3.310044e-06, 3.309519e-06, 3.305227e-06, 3.309578e-06, 
    3.266824e-06, 3.265614e-06, 3.261415e-06, 3.264701e-06, 3.258719e-06, 
    3.262065e-06, 3.26399e-06, 3.271417e-06, 3.273049e-06, 3.274562e-06, 
    3.277554e-06, 3.281395e-06, 3.288148e-06, 3.294675e-06, 3.300072e-06, 
    3.299676e-06, 3.299815e-06, 3.301022e-06, 3.298033e-06, 3.301513e-06, 
    3.302096e-06, 3.300569e-06, 3.309449e-06, 3.306909e-06, 3.309508e-06, 
    3.307854e-06, 3.266007e-06, 3.268041e-06, 3.266943e-06, 3.269006e-06, 
    3.267554e-06, 3.274017e-06, 3.275957e-06, 3.285055e-06, 3.281319e-06, 
    3.287269e-06, 3.281923e-06, 3.282869e-06, 3.28746e-06, 3.282212e-06, 
    3.294347e-06, 3.285907e-06, 3.301069e-06, 3.292607e-06, 3.30156e-06, 
    3.300048e-06, 3.302552e-06, 3.304796e-06, 3.307622e-06, 3.312844e-06, 
    3.311634e-06, 3.316008e-06, 3.271067e-06, 3.273702e-06, 3.273471e-06, 
    3.276232e-06, 3.278274e-06, 3.282706e-06, 3.289831e-06, 3.28715e-06, 
    3.292075e-06, 3.293065e-06, 3.285583e-06, 3.290173e-06, 3.275467e-06, 
    3.277837e-06, 3.276427e-06, 3.271274e-06, 3.287766e-06, 3.27929e-06, 
    3.295601e-06, 3.290356e-06, 3.304476e-06, 3.297757e-06, 3.310968e-06, 
    3.316631e-06, 3.321982e-06, 3.328237e-06, 3.275142e-06, 3.27335e-06, 
    3.27656e-06, 3.281002e-06, 3.285135e-06, 3.290637e-06, 3.291201e-06, 
    3.292233e-06, 3.295547e-06, 3.297801e-06, 3.292558e-06, 3.298367e-06, 
    3.278384e-06, 3.288503e-06, 3.272672e-06, 3.27743e-06, 3.280741e-06, 
    3.279289e-06, 3.286844e-06, 3.288627e-06, 3.296524e-06, 3.292132e-06, 
    3.315231e-06, 3.305267e-06, 3.333016e-06, 3.325231e-06, 3.272724e-06, 
    3.275137e-06, 3.283542e-06, 3.27954e-06, 3.291005e-06, 3.294471e-06, 
    3.296777e-06, 3.299726e-06, 3.300046e-06, 3.301795e-06, 3.298929e-06, 
    3.301682e-06, 3.290648e-06, 3.295924e-06, 3.282581e-06, 3.285667e-06, 
    3.284247e-06, 3.28269e-06, 3.287499e-06, 3.29263e-06, 3.292742e-06, 
    3.295026e-06, 3.299672e-06, 3.291052e-06, 3.316513e-06, 3.301146e-06, 
    3.277768e-06, 3.282419e-06, 3.283086e-06, 3.281283e-06, 3.293551e-06, 
    3.289099e-06, 3.301753e-06, 3.298498e-06, 3.303834e-06, 3.301181e-06, 
    3.30079e-06, 3.297388e-06, 3.295272e-06, 3.289302e-06, 3.284972e-06, 
    3.281544e-06, 3.282341e-06, 3.286108e-06, 3.292945e-06, 3.300073e-06, 
    3.298649e-06, 3.303428e-06, 3.290172e-06, 3.296088e-06, 3.293408e-06, 
    3.299378e-06, 3.287078e-06, 3.297635e-06, 3.284548e-06, 3.285638e-06, 
    3.28901e-06, 3.296445e-06, 3.297957e-06, 3.299567e-06, 3.298574e-06, 
    3.293119e-06, 3.292332e-06, 3.288929e-06, 3.287989e-06, 3.2854e-06, 
    3.283258e-06, 3.285215e-06, 3.287271e-06, 3.293122e-06, 3.299046e-06, 
    3.304827e-06, 3.306245e-06, 3.313012e-06, 3.307498e-06, 3.316598e-06, 
    3.308853e-06, 3.322279e-06, 3.298215e-06, 3.308632e-06, 3.289165e-06, 
    3.291186e-06, 3.295479e-06, 3.303901e-06, 3.299353e-06, 3.304674e-06, 
    3.292302e-06, 3.286237e-06, 3.284673e-06, 3.281752e-06, 3.284739e-06, 
    3.284496e-06, 3.287358e-06, 3.286438e-06, 3.293317e-06, 3.28962e-06, 
    3.30078e-06, 3.304633e-06, 3.315548e-06, 3.32226e-06, 3.329115e-06, 
    3.332145e-06, 3.333068e-06, 3.333454e-06 ;

 QVEGE =
  -6.4823e-07, -6.477904e-07, -6.478738e-07, -6.475231e-07, -6.477144e-07, 
    -6.474871e-07, -6.481369e-07, -6.477765e-07, -6.480044e-07, 
    -6.481849e-07, -6.468516e-07, -6.475064e-07, -6.461358e-07, 
    -6.465586e-07, -6.454831e-07, -6.462071e-07, -6.453341e-07, 
    -6.454948e-07, -6.449875e-07, -6.451326e-07, -6.444997e-07, 
    -6.449203e-07, -6.441542e-07, -6.445953e-07, -6.4453e-07, -6.449357e-07, 
    -6.47366e-07, -6.469356e-07, -6.473935e-07, -6.473317e-07, -6.473574e-07, 
    -6.477136e-07, -6.478986e-07, -6.482572e-07, -6.481906e-07, 
    -6.479237e-07, -6.473037e-07, -6.475086e-07, -6.469734e-07, 
    -6.469853e-07, -6.463993e-07, -6.466638e-07, -6.456701e-07, -6.4595e-07, 
    -6.451264e-07, -6.453363e-07, -6.451378e-07, -6.451968e-07, -6.45137e-07, 
    -6.454441e-07, -6.453132e-07, -6.455799e-07, -6.466161e-07, 
    -6.463148e-07, -6.472188e-07, -6.477767e-07, -6.481228e-07, 
    -6.483744e-07, -6.483389e-07, -6.48273e-07, -6.479223e-07, -6.475835e-07, 
    -6.473272e-07, -6.471567e-07, -6.469871e-07, -6.465019e-07, 
    -6.462242e-07, -6.456174e-07, -6.457199e-07, -6.455401e-07, 
    -6.453567e-07, -6.450586e-07, -6.451066e-07, -6.449768e-07, 
    -6.455392e-07, -6.451687e-07, -6.45778e-07, -6.456143e-07, -6.469723e-07, 
    -6.474519e-07, -6.476817e-07, -6.478589e-07, -6.483123e-07, 
    -6.480012e-07, -6.481246e-07, -6.47824e-07, -6.47637e-07, -6.477282e-07, 
    -6.47152e-07, -6.473777e-07, -6.462078e-07, -6.467108e-07, -6.453781e-07, 
    -6.456982e-07, -6.453e-07, -6.455019e-07, -6.451583e-07, -6.454675e-07, 
    -6.449259e-07, -6.448111e-07, -6.448903e-07, -6.44575e-07, -6.454855e-07, 
    -6.451408e-07, -6.477322e-07, -6.477176e-07, -6.476454e-07, 
    -6.479626e-07, -6.479802e-07, -6.482606e-07, -6.480083e-07, 
    -6.479033e-07, -6.476236e-07, -6.474637e-07, -6.473093e-07, 
    -6.469684e-07, -6.465959e-07, -6.460643e-07, -6.456779e-07, 
    -6.454176e-07, -6.455752e-07, -6.454363e-07, -6.455928e-07, 
    -6.456646e-07, -6.448562e-07, -6.453139e-07, -6.446205e-07, -6.44658e-07, 
    -6.449749e-07, -6.446537e-07, -6.477067e-07, -6.477923e-07, 
    -6.480985e-07, -6.478588e-07, -6.482906e-07, -6.480531e-07, 
    -6.479186e-07, -6.473797e-07, -6.472534e-07, -6.47146e-07, -6.469264e-07, 
    -6.466505e-07, -6.46167e-07, -6.457416e-07, -6.453447e-07, -6.453732e-07, 
    -6.453635e-07, -6.452779e-07, -6.454943e-07, -6.452419e-07, 
    -6.452025e-07, -6.453103e-07, -6.446631e-07, -6.448482e-07, 
    -6.446588e-07, -6.447785e-07, -6.477637e-07, -6.476182e-07, 
    -6.476973e-07, -6.475503e-07, -6.476563e-07, -6.471925e-07, -6.47053e-07, 
    -6.463956e-07, -6.466577e-07, -6.462317e-07, -6.46612e-07, -6.465465e-07, 
    -6.46231e-07, -6.465895e-07, -6.457713e-07, -6.463377e-07, -6.452744e-07, 
    -6.458563e-07, -6.452385e-07, -6.453465e-07, -6.451644e-07, 
    -6.450043e-07, -6.447967e-07, -6.444213e-07, -6.445071e-07, -6.44187e-07, 
    -6.473982e-07, -6.472116e-07, -6.472222e-07, -6.470223e-07, 
    -6.468766e-07, -6.465544e-07, -6.460428e-07, -6.462334e-07, 
    -6.458766e-07, -6.458068e-07, -6.463455e-07, -6.460207e-07, 
    -6.470819e-07, -6.469161e-07, -6.470103e-07, -6.473869e-07, 
    -6.461976e-07, -6.468104e-07, -6.456725e-07, -6.460034e-07, -6.45028e-07, 
    -6.455218e-07, -6.445557e-07, -6.441545e-07, -6.437471e-07, -6.43301e-07, 
    -6.471031e-07, -6.472308e-07, -6.469969e-07, -6.466864e-07, 
    -6.463815e-07, -6.459842e-07, -6.459402e-07, -6.458674e-07, 
    -6.456729e-07, -6.455101e-07, -6.458499e-07, -6.454687e-07, 
    -6.468895e-07, -6.461416e-07, -6.472844e-07, -6.469468e-07, 
    -6.467021e-07, -6.468035e-07, -6.462537e-07, -6.46126e-07, -6.456087e-07, 
    -6.458723e-07, -6.442589e-07, -6.449788e-07, -6.429395e-07, 
    -6.435187e-07, -6.472768e-07, -6.471008e-07, -6.465002e-07, 
    -6.467845e-07, -6.459545e-07, -6.457538e-07, -6.455834e-07, 
    -6.453746e-07, -6.453477e-07, -6.452228e-07, -6.454279e-07, 
    -6.452287e-07, -6.459834e-07, -6.456474e-07, -6.465618e-07, 
    -6.463429e-07, -6.464417e-07, -6.465543e-07, -6.462072e-07, 
    -6.458461e-07, -6.458288e-07, -6.457163e-07, -6.454092e-07, -6.45951e-07, 
    -6.441831e-07, -6.452977e-07, -6.469098e-07, -6.465863e-07, 
    -6.465286e-07, -6.46656e-07, -6.457724e-07, -6.460947e-07, -6.452245e-07, 
    -6.454593e-07, -6.450718e-07, -6.452655e-07, -6.452943e-07, -6.4554e-07, 
    -6.456951e-07, -6.460817e-07, -6.46394e-07, -6.466364e-07, -6.465794e-07, 
    -6.463127e-07, -6.458217e-07, -6.453495e-07, -6.454549e-07, 
    -6.451012e-07, -6.460153e-07, -6.456395e-07, -6.457868e-07, -6.45397e-07, 
    -6.462407e-07, -6.455518e-07, -6.464198e-07, -6.463418e-07, -6.46101e-07, 
    -6.456202e-07, -6.454988e-07, -6.453861e-07, -6.454537e-07, 
    -6.458075e-07, -6.458613e-07, -6.461045e-07, -6.461762e-07, 
    -6.463581e-07, -6.465131e-07, -6.463738e-07, -6.462295e-07, 
    -6.458034e-07, -6.454245e-07, -6.450035e-07, -6.448964e-07, 
    -6.444248e-07, -6.448221e-07, -6.441788e-07, -6.447459e-07, 
    -6.437515e-07, -6.454976e-07, -6.447431e-07, -6.460868e-07, 
    -6.459408e-07, -6.45688e-07, -6.450796e-07, -6.453988e-07, -6.450208e-07, 
    -6.458627e-07, -6.463083e-07, -6.464116e-07, -6.466234e-07, 
    -6.464068e-07, -6.46424e-07, -6.462168e-07, -6.462828e-07, -6.45789e-07, 
    -6.460543e-07, -6.452976e-07, -6.450214e-07, -6.44224e-07, -6.437371e-07, 
    -6.432229e-07, -6.43e-07, -6.429311e-07, -6.429029e-07 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  84.71109, 84.71065, 84.71073, 84.71039, 84.71057, 84.71035, 84.711, 
    84.71063, 84.71086, 84.71104, 84.70977, 84.71037, 84.70921, 84.70954, 
    84.70829, 84.70927, 84.70818, 84.70831, 84.70795, 84.70805, 84.70761, 
    84.7079, 84.70739, 84.70768, 84.70763, 84.70791, 84.71024, 84.70984, 
    84.71027, 84.71021, 84.71024, 84.71057, 84.71075, 84.71112, 84.71105, 
    84.71078, 84.71018, 84.71037, 84.70988, 84.70989, 84.70942, 84.70963, 
    84.70843, 84.70908, 84.70804, 84.70819, 84.70805, 84.70809, 84.70805, 
    84.70827, 84.70818, 84.70837, 84.70959, 84.70935, 84.71011, 84.71062, 
    84.71098, 84.71124, 84.7112, 84.71114, 84.71078, 84.71045, 84.71021, 
    84.71005, 84.7099, 84.70949, 84.70928, 84.70839, 84.70847, 84.70834, 
    84.70821, 84.70799, 84.70803, 84.70794, 84.70834, 84.70807, 84.70895, 
    84.70839, 84.70987, 84.71032, 84.71053, 84.71072, 84.71118, 84.71085, 
    84.71098, 84.71068, 84.71049, 84.71059, 84.71004, 84.71025, 84.70927, 
    84.70966, 84.70822, 84.70845, 84.70816, 84.70831, 84.70806, 84.70828, 
    84.7079, 84.70782, 84.70788, 84.70766, 84.7083, 84.70805, 84.71059, 
    84.71057, 84.7105, 84.71082, 84.71084, 84.71113, 84.71087, 84.71076, 
    84.71049, 84.71033, 84.71019, 84.70988, 84.70957, 84.70916, 84.70844, 
    84.70824, 84.70836, 84.70826, 84.70837, 84.70843, 84.70786, 84.70818, 
    84.7077, 84.70772, 84.70794, 84.70772, 84.71056, 84.71065, 84.71096, 
    84.71072, 84.71116, 84.71091, 84.71077, 84.71025, 84.71014, 84.71004, 
    84.70985, 84.70962, 84.70924, 84.70848, 84.7082, 84.70821, 84.70821, 
    84.70815, 84.70831, 84.70812, 84.70809, 84.70817, 84.70773, 84.70785, 
    84.70773, 84.7078, 84.71062, 84.71048, 84.71056, 84.71041, 84.71051, 
    84.71008, 84.70995, 84.70941, 84.70963, 84.70929, 84.70959, 84.70953, 
    84.70928, 84.70957, 84.7085, 84.70937, 84.70815, 84.709, 84.70812, 
    84.7082, 84.70807, 84.70795, 84.70782, 84.70756, 84.70762, 84.70741, 
    84.71027, 84.7101, 84.71011, 84.70993, 84.7098, 84.70954, 84.70914, 
    84.70929, 84.70902, 84.70897, 84.70938, 84.70913, 84.70998, 84.70983, 
    84.70992, 84.71026, 84.70926, 84.70975, 84.70843, 84.70911, 84.70797, 
    84.70832, 84.70765, 84.70738, 84.70713, 84.70686, 84.71, 84.71012, 
    84.70991, 84.70964, 84.7094, 84.7091, 84.70907, 84.70901, 84.70844, 
    84.70831, 84.709, 84.70828, 84.7098, 84.70922, 84.71017, 84.70985, 
    84.70966, 84.70974, 84.7093, 84.70921, 84.70838, 84.70902, 84.70745, 
    84.70793, 84.70664, 84.70699, 84.71016, 84.71, 84.7095, 84.70972, 
    84.70908, 84.70849, 84.70837, 84.70821, 84.7082, 84.70811, 84.70825, 
    84.70811, 84.7091, 84.70841, 84.70955, 84.70937, 84.70945, 84.70954, 
    84.70927, 84.709, 84.70899, 84.70846, 84.70823, 84.70908, 84.70739, 
    84.70815, 84.70983, 84.70956, 84.70952, 84.70963, 84.70895, 84.70918, 
    84.70811, 84.70827, 84.708, 84.70814, 84.70816, 84.70834, 84.70845, 
    84.70918, 84.70941, 84.70961, 84.70956, 84.70935, 84.70898, 84.7082, 
    84.70827, 84.70802, 84.70913, 84.7084, 84.70895, 84.70823, 84.7093, 
    84.70833, 84.70943, 84.70937, 84.70919, 84.70839, 84.70831, 84.70822, 
    84.70827, 84.70897, 84.70901, 84.70919, 84.70924, 84.70939, 84.70951, 
    84.7094, 84.70928, 84.70897, 84.70825, 84.70795, 84.70789, 84.70756, 
    84.70782, 84.70739, 84.70776, 84.70712, 84.7083, 84.70777, 84.70918, 
    84.70907, 84.70844, 84.708, 84.70824, 84.70796, 84.70901, 84.70934, 
    84.70943, 84.70959, 84.70943, 84.70944, 84.70928, 84.70933, 84.70896, 
    84.70916, 84.70816, 84.70797, 84.70744, 84.70712, 84.70681, 84.70668, 
    84.70664, 84.70663 ;

 RH2M_R =
  84.71109, 84.71065, 84.71073, 84.71039, 84.71057, 84.71035, 84.711, 
    84.71063, 84.71086, 84.71104, 84.70977, 84.71037, 84.70921, 84.70954, 
    84.70829, 84.70927, 84.70818, 84.70831, 84.70795, 84.70805, 84.70761, 
    84.7079, 84.70739, 84.70768, 84.70763, 84.70791, 84.71024, 84.70984, 
    84.71027, 84.71021, 84.71024, 84.71057, 84.71075, 84.71112, 84.71105, 
    84.71078, 84.71018, 84.71037, 84.70988, 84.70989, 84.70942, 84.70963, 
    84.70843, 84.70908, 84.70804, 84.70819, 84.70805, 84.70809, 84.70805, 
    84.70827, 84.70818, 84.70837, 84.70959, 84.70935, 84.71011, 84.71062, 
    84.71098, 84.71124, 84.7112, 84.71114, 84.71078, 84.71045, 84.71021, 
    84.71005, 84.7099, 84.70949, 84.70928, 84.70839, 84.70847, 84.70834, 
    84.70821, 84.70799, 84.70803, 84.70794, 84.70834, 84.70807, 84.70895, 
    84.70839, 84.70987, 84.71032, 84.71053, 84.71072, 84.71118, 84.71085, 
    84.71098, 84.71068, 84.71049, 84.71059, 84.71004, 84.71025, 84.70927, 
    84.70966, 84.70822, 84.70845, 84.70816, 84.70831, 84.70806, 84.70828, 
    84.7079, 84.70782, 84.70788, 84.70766, 84.7083, 84.70805, 84.71059, 
    84.71057, 84.7105, 84.71082, 84.71084, 84.71113, 84.71087, 84.71076, 
    84.71049, 84.71033, 84.71019, 84.70988, 84.70957, 84.70916, 84.70844, 
    84.70824, 84.70836, 84.70826, 84.70837, 84.70843, 84.70786, 84.70818, 
    84.7077, 84.70772, 84.70794, 84.70772, 84.71056, 84.71065, 84.71096, 
    84.71072, 84.71116, 84.71091, 84.71077, 84.71025, 84.71014, 84.71004, 
    84.70985, 84.70962, 84.70924, 84.70848, 84.7082, 84.70821, 84.70821, 
    84.70815, 84.70831, 84.70812, 84.70809, 84.70817, 84.70773, 84.70785, 
    84.70773, 84.7078, 84.71062, 84.71048, 84.71056, 84.71041, 84.71051, 
    84.71008, 84.70995, 84.70941, 84.70963, 84.70929, 84.70959, 84.70953, 
    84.70928, 84.70957, 84.7085, 84.70937, 84.70815, 84.709, 84.70812, 
    84.7082, 84.70807, 84.70795, 84.70782, 84.70756, 84.70762, 84.70741, 
    84.71027, 84.7101, 84.71011, 84.70993, 84.7098, 84.70954, 84.70914, 
    84.70929, 84.70902, 84.70897, 84.70938, 84.70913, 84.70998, 84.70983, 
    84.70992, 84.71026, 84.70926, 84.70975, 84.70843, 84.70911, 84.70797, 
    84.70832, 84.70765, 84.70738, 84.70713, 84.70686, 84.71, 84.71012, 
    84.70991, 84.70964, 84.7094, 84.7091, 84.70907, 84.70901, 84.70844, 
    84.70831, 84.709, 84.70828, 84.7098, 84.70922, 84.71017, 84.70985, 
    84.70966, 84.70974, 84.7093, 84.70921, 84.70838, 84.70902, 84.70745, 
    84.70793, 84.70664, 84.70699, 84.71016, 84.71, 84.7095, 84.70972, 
    84.70908, 84.70849, 84.70837, 84.70821, 84.7082, 84.70811, 84.70825, 
    84.70811, 84.7091, 84.70841, 84.70955, 84.70937, 84.70945, 84.70954, 
    84.70927, 84.709, 84.70899, 84.70846, 84.70823, 84.70908, 84.70739, 
    84.70815, 84.70983, 84.70956, 84.70952, 84.70963, 84.70895, 84.70918, 
    84.70811, 84.70827, 84.708, 84.70814, 84.70816, 84.70834, 84.70845, 
    84.70918, 84.70941, 84.70961, 84.70956, 84.70935, 84.70898, 84.7082, 
    84.70827, 84.70802, 84.70913, 84.7084, 84.70895, 84.70823, 84.7093, 
    84.70833, 84.70943, 84.70937, 84.70919, 84.70839, 84.70831, 84.70822, 
    84.70827, 84.70897, 84.70901, 84.70919, 84.70924, 84.70939, 84.70951, 
    84.7094, 84.70928, 84.70897, 84.70825, 84.70795, 84.70789, 84.70756, 
    84.70782, 84.70739, 84.70776, 84.70712, 84.7083, 84.70777, 84.70918, 
    84.70907, 84.70844, 84.708, 84.70824, 84.70796, 84.70901, 84.70934, 
    84.70943, 84.70959, 84.70943, 84.70944, 84.70928, 84.70933, 84.70896, 
    84.70916, 84.70816, 84.70797, 84.70744, 84.70712, 84.70681, 84.70668, 
    84.70664, 84.70663 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004631664, 0.0004651067, 0.0004647294, 0.0004662944, 0.0004654261, 
    0.0004664508, 0.0004635594, 0.0004651835, 0.0004641466, 0.0004633405, 
    0.000469331, 0.0004663637, 0.0004724115, 0.0004705196, 0.0004752712, 
    0.0004721171, 0.000475907, 0.0004751798, 0.0004773675, 0.0004767407, 
    0.000479539, 0.0004776566, 0.000480989, 0.0004790893, 0.0004793865, 
    0.0004775943, 0.0004669611, 0.000468962, 0.0004668424, 0.0004671278, 
    0.0004669997, 0.0004654439, 0.00046466, 0.0004630174, 0.0004633155, 
    0.0004645218, 0.0004672557, 0.0004663274, 0.0004686661, 0.0004686132, 
    0.0004712165, 0.0004700428, 0.0004744177, 0.0004731742, 0.0004767668, 
    0.0004758633, 0.0004767243, 0.0004764631, 0.0004767276, 0.0004754026, 
    0.0004759702, 0.0004748042, 0.0004702633, 0.0004715983, 0.0004676162, 
    0.0004652217, 0.0004636305, 0.0004625015, 0.0004626609, 0.0004629653, 
    0.0004645287, 0.0004659984, 0.0004671183, 0.0004678674, 0.0004686055, 
    0.0004708402, 0.0004720222, 0.0004746691, 0.0004741912, 0.0004750005, 
    0.0004757734, 0.0004770711, 0.0004768574, 0.0004774292, 0.0004749787, 
    0.0004766074, 0.0004739186, 0.0004746541, 0.0004688075, 0.0004665781, 
    0.0004656311, 0.0004648014, 0.0004627836, 0.0004641771, 0.0004636278, 
    0.0004649343, 0.0004657645, 0.0004653537, 0.0004678879, 0.0004669027, 
    0.0004720922, 0.000469857, 0.0004756833, 0.0004742891, 0.0004760172, 
    0.0004751354, 0.0004766463, 0.0004752864, 0.0004776418, 0.0004781548, 
    0.0004778041, 0.0004791503, 0.0004752107, 0.0004767238, 0.0004653426, 
    0.0004654096, 0.0004657215, 0.0004643501, 0.0004642661, 0.0004630089, 
    0.0004641273, 0.0004646037, 0.0004658124, 0.0004665275, 0.0004672071, 
    0.0004687015, 0.0004703704, 0.0004727036, 0.0004743795, 0.0004755027, 
    0.0004748139, 0.000475422, 0.0004747421, 0.0004744233, 0.0004779625, 
    0.0004759753, 0.0004789566, 0.0004787916, 0.0004774424, 0.00047881, 
    0.0004654565, 0.000465071, 0.000463733, 0.00046478, 0.0004628719, 
    0.0004639401, 0.0004645542, 0.0004669233, 0.0004674436, 0.0004679263, 
    0.0004688793, 0.0004701024, 0.000472248, 0.0004741145, 0.0004758181, 
    0.0004756932, 0.0004757371, 0.0004761177, 0.0004751749, 0.0004762723, 
    0.0004764565, 0.0004759748, 0.0004787693, 0.000477971, 0.0004787878, 
    0.0004782679, 0.0004651962, 0.0004658446, 0.0004654941, 0.0004661531, 
    0.0004656888, 0.000467753, 0.0004683718, 0.0004712668, 0.0004700784, 
    0.0004719694, 0.0004702703, 0.0004705714, 0.0004720312, 0.0004703619, 
    0.0004740116, 0.0004715375, 0.0004761324, 0.0004736624, 0.0004762871, 
    0.0004758103, 0.0004765994, 0.0004773063, 0.0004781952, 0.0004798358, 
    0.0004794557, 0.0004808276, 0.0004668112, 0.0004676523, 0.0004675781, 
    0.0004684581, 0.0004691089, 0.0004705194, 0.0004727816, 0.0004719308, 
    0.0004734923, 0.0004738058, 0.0004714332, 0.0004728901, 0.0004682145, 
    0.0004689701, 0.00046852, 0.0004668768, 0.0004721266, 0.0004694326, 
    0.0004744066, 0.0004729473, 0.0004772053, 0.000475088, 0.0004792466, 
    0.0004810246, 0.0004826968, 0.0004846518, 0.0004681111, 0.0004675395, 
    0.0004685626, 0.0004699783, 0.0004712913, 0.000473037, 0.0004732154, 
    0.0004735424, 0.0004743893, 0.0004751015, 0.0004736459, 0.0004752799, 
    0.0004691456, 0.0004723603, 0.0004673229, 0.0004688401, 0.0004698941, 
    0.0004694315, 0.0004718328, 0.0004723987, 0.0004746984, 0.0004735095, 
    0.0004805857, 0.0004774554, 0.0004861396, 0.0004837133, 0.0004673398, 
    0.0004681088, 0.0004707855, 0.0004695119, 0.0004731533, 0.0004740496, 
    0.0004747779, 0.0004757093, 0.0004758096, 0.0004763615, 0.0004754571, 
    0.0004763256, 0.0004730401, 0.0004745084, 0.0004704788, 0.0004714596, 
    0.0004710083, 0.0004705132, 0.0004720407, 0.0004736682, 0.0004737026, 
    0.0004742244, 0.0004756954, 0.000473167, 0.00048099, 0.0004761595, 
    0.0004689474, 0.0004704289, 0.0004706402, 0.0004700663, 0.0004739596, 
    0.000472549, 0.000476348, 0.0004753212, 0.0004770033, 0.0004761674, 
    0.0004760443, 0.0004749707, 0.0004743022, 0.0004726133, 0.0004712389, 
    0.0004701489, 0.0004704022, 0.0004715995, 0.0004737675, 0.0004758182, 
    0.000475369, 0.0004768747, 0.0004728882, 0.00047456, 0.0004739139, 
    0.0004755984, 0.000471908, 0.0004750524, 0.0004711042, 0.0004714503, 
    0.0004725209, 0.0004746745, 0.0004751504, 0.0004756591, 0.000475345, 
    0.0004738229, 0.0004735734, 0.0004724944, 0.0004721966, 0.0004713744, 
    0.0004706937, 0.0004713156, 0.0004719686, 0.000473823, 0.0004754941, 
    0.0004773157, 0.0004777613, 0.00047989, 0.0004781575, 0.0004810167, 
    0.0004785863, 0.0004827928, 0.000475234, 0.0004785154, 0.0004725695, 
    0.00047321, 0.0004743689, 0.0004770259, 0.0004755911, 0.0004772689, 
    0.0004735635, 0.000471641, 0.0004711433, 0.0004702151, 0.0004711644, 
    0.0004710871, 0.0004719955, 0.0004717035, 0.0004738844, 0.0004727129, 
    0.0004760406, 0.0004772549, 0.0004806833, 0.0004827847, 0.0004849232, 
    0.0004858673, 0.0004861546, 0.0004862747 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.117403e-14, 3.125812e-14, 3.124178e-14, 3.130955e-14, 3.127198e-14, 
    3.131633e-14, 3.11911e-14, 3.126144e-14, 3.121655e-14, 3.118162e-14, 
    3.144085e-14, 3.131257e-14, 3.157399e-14, 3.149233e-14, 3.169734e-14, 
    3.156127e-14, 3.172475e-14, 3.169344e-14, 3.178771e-14, 3.176072e-14, 
    3.18811e-14, 3.180016e-14, 3.194348e-14, 3.186179e-14, 3.187457e-14, 
    3.179749e-14, 3.133843e-14, 3.142488e-14, 3.13333e-14, 3.134563e-14, 
    3.134011e-14, 3.127274e-14, 3.123875e-14, 3.116761e-14, 3.118054e-14, 
    3.12328e-14, 3.135118e-14, 3.131103e-14, 3.141223e-14, 3.140995e-14, 
    3.152244e-14, 3.147174e-14, 3.166058e-14, 3.160698e-14, 3.176184e-14, 
    3.172292e-14, 3.176001e-14, 3.174877e-14, 3.176016e-14, 3.170306e-14, 
    3.172753e-14, 3.167727e-14, 3.148123e-14, 3.15389e-14, 3.136678e-14, 
    3.126307e-14, 3.119418e-14, 3.114524e-14, 3.115216e-14, 3.116534e-14, 
    3.12331e-14, 3.129679e-14, 3.134527e-14, 3.137769e-14, 3.140962e-14, 
    3.150612e-14, 3.155721e-14, 3.167141e-14, 3.165083e-14, 3.168571e-14, 
    3.171904e-14, 3.177495e-14, 3.176575e-14, 3.179037e-14, 3.168481e-14, 
    3.175497e-14, 3.163912e-14, 3.167081e-14, 3.141821e-14, 3.132187e-14, 
    3.128081e-14, 3.124492e-14, 3.115748e-14, 3.121787e-14, 3.119407e-14, 
    3.12507e-14, 3.128666e-14, 3.126889e-14, 3.137858e-14, 3.133595e-14, 
    3.156023e-14, 3.14637e-14, 3.171516e-14, 3.165506e-14, 3.172956e-14, 
    3.169155e-14, 3.175665e-14, 3.169807e-14, 3.179953e-14, 3.18216e-14, 
    3.180652e-14, 3.186446e-14, 3.169482e-14, 3.176e-14, 3.126838e-14, 
    3.127128e-14, 3.12848e-14, 3.122536e-14, 3.122173e-14, 3.116725e-14, 
    3.121574e-14, 3.123637e-14, 3.128875e-14, 3.13197e-14, 3.134912e-14, 
    3.141377e-14, 3.148588e-14, 3.158665e-14, 3.165895e-14, 3.170739e-14, 
    3.16777e-14, 3.170391e-14, 3.167461e-14, 3.166087e-14, 3.181333e-14, 
    3.172775e-14, 3.185613e-14, 3.184904e-14, 3.179095e-14, 3.184984e-14, 
    3.127332e-14, 3.125663e-14, 3.119864e-14, 3.124403e-14, 3.116132e-14, 
    3.120761e-14, 3.123421e-14, 3.133682e-14, 3.135937e-14, 3.138024e-14, 
    3.142147e-14, 3.147434e-14, 3.156699e-14, 3.164752e-14, 3.172099e-14, 
    3.171561e-14, 3.17175e-14, 3.17339e-14, 3.169327e-14, 3.174056e-14, 
    3.174849e-14, 3.172775e-14, 3.184809e-14, 3.181373e-14, 3.184889e-14, 
    3.182652e-14, 3.126206e-14, 3.129014e-14, 3.127496e-14, 3.130349e-14, 
    3.128339e-14, 3.137271e-14, 3.139947e-14, 3.152459e-14, 3.147329e-14, 
    3.155495e-14, 3.14816e-14, 3.14946e-14, 3.155757e-14, 3.148557e-14, 
    3.164306e-14, 3.153629e-14, 3.173453e-14, 3.1628e-14, 3.17412e-14, 
    3.172067e-14, 3.175467e-14, 3.17851e-14, 3.182338e-14, 3.189394e-14, 
    3.187761e-14, 3.19366e-14, 3.133199e-14, 3.136837e-14, 3.136518e-14, 
    3.140325e-14, 3.143139e-14, 3.149236e-14, 3.159003e-14, 3.155332e-14, 
    3.162072e-14, 3.163424e-14, 3.153185e-14, 3.159471e-14, 3.139272e-14, 
    3.142537e-14, 3.140595e-14, 3.133485e-14, 3.156176e-14, 3.144538e-14, 
    3.166015e-14, 3.159722e-14, 3.178076e-14, 3.168951e-14, 3.186862e-14, 
    3.194501e-14, 3.201693e-14, 3.210078e-14, 3.138824e-14, 3.136352e-14, 
    3.140778e-14, 3.146894e-14, 3.15257e-14, 3.160106e-14, 3.160878e-14, 
    3.162288e-14, 3.16594e-14, 3.16901e-14, 3.162732e-14, 3.16978e-14, 
    3.14329e-14, 3.157186e-14, 3.135416e-14, 3.141976e-14, 3.146534e-14, 
    3.144537e-14, 3.154913e-14, 3.157356e-14, 3.167273e-14, 3.16215e-14, 
    3.192615e-14, 3.17915e-14, 3.216462e-14, 3.206052e-14, 3.135488e-14, 
    3.138816e-14, 3.150384e-14, 3.144882e-14, 3.16061e-14, 3.164474e-14, 
    3.167616e-14, 3.171629e-14, 3.172063e-14, 3.17444e-14, 3.170545e-14, 
    3.174287e-14, 3.160122e-14, 3.166454e-14, 3.149064e-14, 3.1533e-14, 
    3.151352e-14, 3.149214e-14, 3.155811e-14, 3.162831e-14, 3.162983e-14, 
    3.16523e-14, 3.171559e-14, 3.160673e-14, 3.194346e-14, 3.173562e-14, 
    3.142442e-14, 3.148841e-14, 3.149758e-14, 3.14728e-14, 3.164088e-14, 
    3.158001e-14, 3.174382e-14, 3.169959e-14, 3.177206e-14, 3.173605e-14, 
    3.173075e-14, 3.168448e-14, 3.165566e-14, 3.15828e-14, 3.152347e-14, 
    3.147639e-14, 3.148735e-14, 3.153904e-14, 3.16326e-14, 3.172101e-14, 
    3.170165e-14, 3.176656e-14, 3.15947e-14, 3.166678e-14, 3.163893e-14, 
    3.171157e-14, 3.155234e-14, 3.168786e-14, 3.151765e-14, 3.153259e-14, 
    3.15788e-14, 3.167165e-14, 3.169223e-14, 3.171414e-14, 3.170062e-14, 
    3.163498e-14, 3.162423e-14, 3.157769e-14, 3.156482e-14, 3.152934e-14, 
    3.149994e-14, 3.15268e-14, 3.155498e-14, 3.163502e-14, 3.170705e-14, 
    3.178553e-14, 3.180474e-14, 3.189624e-14, 3.182172e-14, 3.194461e-14, 
    3.184008e-14, 3.202096e-14, 3.169575e-14, 3.183706e-14, 3.158092e-14, 
    3.160856e-14, 3.165849e-14, 3.177299e-14, 3.171123e-14, 3.178346e-14, 
    3.162381e-14, 3.154081e-14, 3.151936e-14, 3.147925e-14, 3.152027e-14, 
    3.151694e-14, 3.155617e-14, 3.154356e-14, 3.163768e-14, 3.158714e-14, 
    3.173061e-14, 3.17829e-14, 3.193041e-14, 3.202068e-14, 3.21125e-14, 
    3.215298e-14, 3.216531e-14, 3.217045e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.036534e-14, 1.039333e-14, 1.038789e-14, 1.041044e-14, 1.039794e-14, 
    1.04127e-14, 1.037102e-14, 1.039443e-14, 1.037949e-14, 1.036786e-14, 
    1.045414e-14, 1.041145e-14, 1.049846e-14, 1.047128e-14, 1.053951e-14, 
    1.049422e-14, 1.054863e-14, 1.053821e-14, 1.056959e-14, 1.05606e-14, 
    1.060067e-14, 1.057373e-14, 1.062143e-14, 1.059425e-14, 1.05985e-14, 
    1.057284e-14, 1.042006e-14, 1.044883e-14, 1.041835e-14, 1.042245e-14, 
    1.042061e-14, 1.039819e-14, 1.038688e-14, 1.03632e-14, 1.036751e-14, 
    1.03849e-14, 1.04243e-14, 1.041094e-14, 1.044462e-14, 1.044386e-14, 
    1.04813e-14, 1.046442e-14, 1.052728e-14, 1.050944e-14, 1.056098e-14, 
    1.054802e-14, 1.056037e-14, 1.055663e-14, 1.056042e-14, 1.054141e-14, 
    1.054956e-14, 1.053283e-14, 1.046758e-14, 1.048678e-14, 1.042949e-14, 
    1.039497e-14, 1.037204e-14, 1.035576e-14, 1.035806e-14, 1.036245e-14, 
    1.0385e-14, 1.04062e-14, 1.042233e-14, 1.043312e-14, 1.044375e-14, 
    1.047587e-14, 1.049287e-14, 1.053088e-14, 1.052403e-14, 1.053564e-14, 
    1.054673e-14, 1.056534e-14, 1.056228e-14, 1.057047e-14, 1.053534e-14, 
    1.055869e-14, 1.052013e-14, 1.053068e-14, 1.044661e-14, 1.041454e-14, 
    1.040088e-14, 1.038893e-14, 1.035983e-14, 1.037993e-14, 1.037201e-14, 
    1.039086e-14, 1.040283e-14, 1.039691e-14, 1.043342e-14, 1.041923e-14, 
    1.049388e-14, 1.046175e-14, 1.054544e-14, 1.052544e-14, 1.055023e-14, 
    1.053759e-14, 1.055925e-14, 1.053975e-14, 1.057352e-14, 1.058087e-14, 
    1.057585e-14, 1.059514e-14, 1.053867e-14, 1.056037e-14, 1.039674e-14, 
    1.039771e-14, 1.04022e-14, 1.038243e-14, 1.038122e-14, 1.036308e-14, 
    1.037922e-14, 1.038609e-14, 1.040352e-14, 1.041382e-14, 1.042361e-14, 
    1.044513e-14, 1.046913e-14, 1.050267e-14, 1.052673e-14, 1.054286e-14, 
    1.053297e-14, 1.05417e-14, 1.053194e-14, 1.052737e-14, 1.057812e-14, 
    1.054963e-14, 1.059236e-14, 1.059e-14, 1.057067e-14, 1.059027e-14, 
    1.039838e-14, 1.039283e-14, 1.037353e-14, 1.038864e-14, 1.036111e-14, 
    1.037652e-14, 1.038537e-14, 1.041952e-14, 1.042702e-14, 1.043397e-14, 
    1.044769e-14, 1.046529e-14, 1.049613e-14, 1.052293e-14, 1.054738e-14, 
    1.054559e-14, 1.054622e-14, 1.055168e-14, 1.053815e-14, 1.05539e-14, 
    1.055654e-14, 1.054963e-14, 1.058968e-14, 1.057825e-14, 1.058995e-14, 
    1.058251e-14, 1.039464e-14, 1.040398e-14, 1.039893e-14, 1.040843e-14, 
    1.040174e-14, 1.043146e-14, 1.044037e-14, 1.048202e-14, 1.046494e-14, 
    1.049212e-14, 1.046771e-14, 1.047203e-14, 1.049299e-14, 1.046903e-14, 
    1.052145e-14, 1.048591e-14, 1.055189e-14, 1.051643e-14, 1.055411e-14, 
    1.054728e-14, 1.055859e-14, 1.056872e-14, 1.058146e-14, 1.060495e-14, 
    1.059951e-14, 1.061914e-14, 1.041791e-14, 1.043002e-14, 1.042896e-14, 
    1.044163e-14, 1.045099e-14, 1.047129e-14, 1.050379e-14, 1.049158e-14, 
    1.051401e-14, 1.051851e-14, 1.048443e-14, 1.050535e-14, 1.043812e-14, 
    1.044899e-14, 1.044253e-14, 1.041886e-14, 1.049438e-14, 1.045565e-14, 
    1.052713e-14, 1.050619e-14, 1.056728e-14, 1.05369e-14, 1.059652e-14, 
    1.062194e-14, 1.064588e-14, 1.067379e-14, 1.043663e-14, 1.042841e-14, 
    1.044314e-14, 1.046349e-14, 1.048238e-14, 1.050746e-14, 1.051003e-14, 
    1.051473e-14, 1.052688e-14, 1.05371e-14, 1.051621e-14, 1.053966e-14, 
    1.04515e-14, 1.049775e-14, 1.042529e-14, 1.044712e-14, 1.04623e-14, 
    1.045565e-14, 1.049018e-14, 1.049831e-14, 1.053132e-14, 1.051427e-14, 
    1.061567e-14, 1.057085e-14, 1.069504e-14, 1.066039e-14, 1.042553e-14, 
    1.043661e-14, 1.047511e-14, 1.04568e-14, 1.050914e-14, 1.0522e-14, 
    1.053246e-14, 1.054582e-14, 1.054726e-14, 1.055517e-14, 1.054221e-14, 
    1.055466e-14, 1.050752e-14, 1.052859e-14, 1.047071e-14, 1.048481e-14, 
    1.047833e-14, 1.047121e-14, 1.049317e-14, 1.051653e-14, 1.051704e-14, 
    1.052452e-14, 1.054558e-14, 1.050935e-14, 1.062143e-14, 1.055225e-14, 
    1.044868e-14, 1.046997e-14, 1.047303e-14, 1.046478e-14, 1.052072e-14, 
    1.050046e-14, 1.055498e-14, 1.054026e-14, 1.056438e-14, 1.05524e-14, 
    1.055063e-14, 1.053523e-14, 1.052564e-14, 1.050139e-14, 1.048164e-14, 
    1.046597e-14, 1.046962e-14, 1.048682e-14, 1.051796e-14, 1.054739e-14, 
    1.054094e-14, 1.056255e-14, 1.050535e-14, 1.052934e-14, 1.052007e-14, 
    1.054425e-14, 1.049125e-14, 1.053636e-14, 1.04797e-14, 1.048468e-14, 
    1.050006e-14, 1.053096e-14, 1.053781e-14, 1.05451e-14, 1.05406e-14, 
    1.051876e-14, 1.051518e-14, 1.049969e-14, 1.04954e-14, 1.04836e-14, 
    1.047381e-14, 1.048275e-14, 1.049213e-14, 1.051877e-14, 1.054274e-14, 
    1.056886e-14, 1.057526e-14, 1.060571e-14, 1.058091e-14, 1.062181e-14, 
    1.058702e-14, 1.064722e-14, 1.053898e-14, 1.058602e-14, 1.050076e-14, 
    1.050996e-14, 1.052658e-14, 1.056469e-14, 1.054413e-14, 1.056818e-14, 
    1.051504e-14, 1.048741e-14, 1.048027e-14, 1.046693e-14, 1.048058e-14, 
    1.047947e-14, 1.049252e-14, 1.048833e-14, 1.051965e-14, 1.050283e-14, 
    1.055058e-14, 1.056799e-14, 1.061708e-14, 1.064713e-14, 1.067769e-14, 
    1.069117e-14, 1.069527e-14, 1.069698e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.365502e-11, -8.402314e-11, -8.395157e-11, -8.424849e-11, -8.408378e-11, 
    -8.427821e-11, -8.372965e-11, -8.403776e-11, -8.384107e-11, 
    -8.368815e-11, -8.482471e-11, -8.426174e-11, -8.540944e-11, 
    -8.505041e-11, -8.595229e-11, -8.535358e-11, -8.607302e-11, 
    -8.593501e-11, -8.635035e-11, -8.623136e-11, -8.676262e-11, 
    -8.640526e-11, -8.7038e-11, -8.667728e-11, -8.673371e-11, -8.639348e-11, 
    -8.437502e-11, -8.475463e-11, -8.435253e-11, -8.440666e-11, 
    -8.438238e-11, -8.408719e-11, -8.393844e-11, -8.362688e-11, 
    -8.368344e-11, -8.391227e-11, -8.4431e-11, -8.425491e-11, -8.469869e-11, 
    -8.468867e-11, -8.518272e-11, -8.495996e-11, -8.579034e-11, 
    -8.555433e-11, -8.623633e-11, -8.606481e-11, -8.622827e-11, 
    -8.617871e-11, -8.622892e-11, -8.597738e-11, -8.608515e-11, -8.58638e-11, 
    -8.500169e-11, -8.525506e-11, -8.449937e-11, -8.404499e-11, 
    -8.374317e-11, -8.352899e-11, -8.355927e-11, -8.3617e-11, -8.391361e-11, 
    -8.419248e-11, -8.4405e-11, -8.454715e-11, -8.468723e-11, -8.511123e-11, 
    -8.533562e-11, -8.583807e-11, -8.574739e-11, -8.590101e-11, 
    -8.604775e-11, -8.629414e-11, -8.625358e-11, -8.636213e-11, 
    -8.589695e-11, -8.620612e-11, -8.569574e-11, -8.583533e-11, 
    -8.472534e-11, -8.430242e-11, -8.412268e-11, -8.396533e-11, 
    -8.358255e-11, -8.384689e-11, -8.374269e-11, -8.399059e-11, 
    -8.414812e-11, -8.407021e-11, -8.455105e-11, -8.436411e-11, 
    -8.534892e-11, -8.492473e-11, -8.603063e-11, -8.5766e-11, -8.609406e-11, 
    -8.592666e-11, -8.62135e-11, -8.595535e-11, -8.640253e-11, -8.649991e-11, 
    -8.643337e-11, -8.668898e-11, -8.594103e-11, -8.622827e-11, 
    -8.406803e-11, -8.408074e-11, -8.413993e-11, -8.387972e-11, -8.38638e-11, 
    -8.362533e-11, -8.383752e-11, -8.392788e-11, -8.415725e-11, 
    -8.429293e-11, -8.44219e-11, -8.470547e-11, -8.502217e-11, -8.546502e-11, 
    -8.578315e-11, -8.599641e-11, -8.586564e-11, -8.59811e-11, -8.585203e-11, 
    -8.579154e-11, -8.646343e-11, -8.608616e-11, -8.665221e-11, 
    -8.662088e-11, -8.636471e-11, -8.662442e-11, -8.408966e-11, 
    -8.401654e-11, -8.376267e-11, -8.396134e-11, -8.359936e-11, 
    -8.380199e-11, -8.39185e-11, -8.436803e-11, -8.446678e-11, -8.455837e-11, 
    -8.473924e-11, -8.497136e-11, -8.537857e-11, -8.573287e-11, 
    -8.605629e-11, -8.603259e-11, -8.604093e-11, -8.611319e-11, 
    -8.593421e-11, -8.614257e-11, -8.617754e-11, -8.608611e-11, 
    -8.661669e-11, -8.646511e-11, -8.662022e-11, -8.652152e-11, -8.40403e-11, 
    -8.416334e-11, -8.409685e-11, -8.422188e-11, -8.41338e-11, -8.452544e-11, 
    -8.464287e-11, -8.519229e-11, -8.49668e-11, -8.532566e-11, -8.500325e-11, 
    -8.506038e-11, -8.533738e-11, -8.502067e-11, -8.571334e-11, 
    -8.524374e-11, -8.6116e-11, -8.564708e-11, -8.614538e-11, -8.605489e-11, 
    -8.620471e-11, -8.63389e-11, -8.650771e-11, -8.68192e-11, -8.674706e-11, 
    -8.700755e-11, -8.434676e-11, -8.450635e-11, -8.449229e-11, 
    -8.465929e-11, -8.478281e-11, -8.505049e-11, -8.547984e-11, 
    -8.531838e-11, -8.561479e-11, -8.567429e-11, -8.522398e-11, 
    -8.550047e-11, -8.461314e-11, -8.475651e-11, -8.467115e-11, 
    -8.435935e-11, -8.53556e-11, -8.484433e-11, -8.578841e-11, -8.551145e-11, 
    -8.631977e-11, -8.591778e-11, -8.670736e-11, -8.704491e-11, 
    -8.736258e-11, -8.773383e-11, -8.459344e-11, -8.4485e-11, -8.467915e-11, 
    -8.494778e-11, -8.5197e-11, -8.552834e-11, -8.556224e-11, -8.562431e-11, 
    -8.578509e-11, -8.592028e-11, -8.564395e-11, -8.595417e-11, 
    -8.478978e-11, -8.539998e-11, -8.444401e-11, -8.473189e-11, 
    -8.493194e-11, -8.484417e-11, -8.529993e-11, -8.540735e-11, 
    -8.584385e-11, -8.561821e-11, -8.696161e-11, -8.636725e-11, 
    -8.801649e-11, -8.755561e-11, -8.444712e-11, -8.459306e-11, -8.5101e-11, 
    -8.485932e-11, -8.555046e-11, -8.572058e-11, -8.585887e-11, 
    -8.603566e-11, -8.605474e-11, -8.615949e-11, -8.598784e-11, -8.61527e-11, 
    -8.552905e-11, -8.580774e-11, -8.504293e-11, -8.522909e-11, 
    -8.514345e-11, -8.504951e-11, -8.533942e-11, -8.56483e-11, -8.565489e-11, 
    -8.575393e-11, -8.603305e-11, -8.555326e-11, -8.703834e-11, 
    -8.612121e-11, -8.475221e-11, -8.503333e-11, -8.507346e-11, 
    -8.496457e-11, -8.570353e-11, -8.543578e-11, -8.615694e-11, 
    -8.596203e-11, -8.628138e-11, -8.612269e-11, -8.609934e-11, 
    -8.589553e-11, -8.576864e-11, -8.544806e-11, -8.518721e-11, 
    -8.498036e-11, -8.502846e-11, -8.525568e-11, -8.566719e-11, 
    -8.605647e-11, -8.59712e-11, -8.625711e-11, -8.550034e-11, -8.581767e-11, 
    -8.569503e-11, -8.601482e-11, -8.53141e-11, -8.591083e-11, -8.516157e-11, 
    -8.522726e-11, -8.543046e-11, -8.58392e-11, -8.592962e-11, -8.602618e-11, 
    -8.596659e-11, -8.567764e-11, -8.563029e-11, -8.542552e-11, 
    -8.536899e-11, -8.521295e-11, -8.508379e-11, -8.520181e-11, 
    -8.532576e-11, -8.567776e-11, -8.599497e-11, -8.634081e-11, 
    -8.642544e-11, -8.682956e-11, -8.650061e-11, -8.704346e-11, 
    -8.658196e-11, -8.738082e-11, -8.59454e-11, -8.656836e-11, -8.54397e-11, 
    -8.556129e-11, -8.578123e-11, -8.628565e-11, -8.601331e-11, -8.63318e-11, 
    -8.562843e-11, -8.526353e-11, -8.516909e-11, -8.499294e-11, 
    -8.517312e-11, -8.515846e-11, -8.533088e-11, -8.527547e-11, 
    -8.568944e-11, -8.546708e-11, -8.609876e-11, -8.632928e-11, 
    -8.698026e-11, -8.737933e-11, -8.778554e-11, -8.796489e-11, 
    -8.801947e-11, -8.804229e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -2.016235e-12, -2.025105e-12, -2.023381e-12, -2.030535e-12, -2.026566e-12, 
    -2.031251e-12, -2.018033e-12, -2.025457e-12, -2.020718e-12, 
    -2.017033e-12, -2.04442e-12, -2.030854e-12, -2.05851e-12, -2.049858e-12, 
    -2.071591e-12, -2.057164e-12, -2.074499e-12, -2.071174e-12, 
    -2.081182e-12, -2.078315e-12, -2.091116e-12, -2.082505e-12, 
    -2.097752e-12, -2.08906e-12, -2.09042e-12, -2.082221e-12, -2.033584e-12, 
    -2.042731e-12, -2.033042e-12, -2.034346e-12, -2.033761e-12, 
    -2.026648e-12, -2.023064e-12, -2.015556e-12, -2.016919e-12, 
    -2.022433e-12, -2.034933e-12, -2.03069e-12, -2.041383e-12, -2.041142e-12, 
    -2.053047e-12, -2.047679e-12, -2.067688e-12, -2.062001e-12, 
    -2.078435e-12, -2.074302e-12, -2.078241e-12, -2.077046e-12, 
    -2.078256e-12, -2.072195e-12, -2.074792e-12, -2.069458e-12, 
    -2.048684e-12, -2.05479e-12, -2.036581e-12, -2.025632e-12, -2.018359e-12, 
    -2.013198e-12, -2.013927e-12, -2.015318e-12, -2.022466e-12, 
    -2.029185e-12, -2.034306e-12, -2.037732e-12, -2.041107e-12, 
    -2.051324e-12, -2.056731e-12, -2.068838e-12, -2.066653e-12, 
    -2.070355e-12, -2.073891e-12, -2.079828e-12, -2.07885e-12, -2.081466e-12, 
    -2.070257e-12, -2.077707e-12, -2.065408e-12, -2.068772e-12, 
    -2.042026e-12, -2.031835e-12, -2.027504e-12, -2.023712e-12, 
    -2.014488e-12, -2.020858e-12, -2.018347e-12, -2.024321e-12, 
    -2.028117e-12, -2.026239e-12, -2.037825e-12, -2.033321e-12, 
    -2.057052e-12, -2.04683e-12, -2.073478e-12, -2.067101e-12, -2.075007e-12, 
    -2.070973e-12, -2.077885e-12, -2.071664e-12, -2.082439e-12, 
    -2.084786e-12, -2.083183e-12, -2.089342e-12, -2.071319e-12, 
    -2.078241e-12, -2.026187e-12, -2.026493e-12, -2.027919e-12, 
    -2.021649e-12, -2.021266e-12, -2.015519e-12, -2.020632e-12, 
    -2.022809e-12, -2.028336e-12, -2.031606e-12, -2.034714e-12, 
    -2.041547e-12, -2.049178e-12, -2.059849e-12, -2.067515e-12, 
    -2.072654e-12, -2.069503e-12, -2.072284e-12, -2.069175e-12, 
    -2.067717e-12, -2.083907e-12, -2.074816e-12, -2.088456e-12, 
    -2.087701e-12, -2.081528e-12, -2.087786e-12, -2.026708e-12, 
    -2.024946e-12, -2.018828e-12, -2.023616e-12, -2.014893e-12, 
    -2.019776e-12, -2.022583e-12, -2.033415e-12, -2.035795e-12, 
    -2.038002e-12, -2.04236e-12, -2.047954e-12, -2.057766e-12, -2.066303e-12, 
    -2.074096e-12, -2.073525e-12, -2.073726e-12, -2.075467e-12, 
    -2.071155e-12, -2.076175e-12, -2.077018e-12, -2.074815e-12, -2.0876e-12, 
    -2.083947e-12, -2.087685e-12, -2.085307e-12, -2.025518e-12, 
    -2.028483e-12, -2.026881e-12, -2.029894e-12, -2.027771e-12, 
    -2.037209e-12, -2.040038e-12, -2.053277e-12, -2.047844e-12, 
    -2.056491e-12, -2.048722e-12, -2.050099e-12, -2.056774e-12, 
    -2.049142e-12, -2.065833e-12, -2.054517e-12, -2.075535e-12, 
    -2.064236e-12, -2.076243e-12, -2.074063e-12, -2.077673e-12, 
    -2.080906e-12, -2.084974e-12, -2.092479e-12, -2.090741e-12, 
    -2.097018e-12, -2.032903e-12, -2.036748e-12, -2.03641e-12, -2.040434e-12, 
    -2.04341e-12, -2.04986e-12, -2.060206e-12, -2.056316e-12, -2.063458e-12, 
    -2.064892e-12, -2.054041e-12, -2.060703e-12, -2.039322e-12, 
    -2.042777e-12, -2.04072e-12, -2.033207e-12, -2.057212e-12, -2.044893e-12, 
    -2.067642e-12, -2.060968e-12, -2.080445e-12, -2.070759e-12, 
    -2.089785e-12, -2.097918e-12, -2.105573e-12, -2.114519e-12, 
    -2.038847e-12, -2.036234e-12, -2.040913e-12, -2.047385e-12, 
    -2.053391e-12, -2.061375e-12, -2.062192e-12, -2.063687e-12, 
    -2.067562e-12, -2.070819e-12, -2.06416e-12, -2.071636e-12, -2.043578e-12, 
    -2.058282e-12, -2.035246e-12, -2.042183e-12, -2.047004e-12, 
    -2.044889e-12, -2.055871e-12, -2.058459e-12, -2.068978e-12, -2.06354e-12, 
    -2.095911e-12, -2.081589e-12, -2.12133e-12, -2.110224e-12, -2.035321e-12, 
    -2.038838e-12, -2.051077e-12, -2.045254e-12, -2.061908e-12, 
    -2.066007e-12, -2.069339e-12, -2.073599e-12, -2.074059e-12, 
    -2.076583e-12, -2.072447e-12, -2.07642e-12, -2.061392e-12, -2.068107e-12, 
    -2.049678e-12, -2.054164e-12, -2.0521e-12, -2.049837e-12, -2.056823e-12, 
    -2.064265e-12, -2.064424e-12, -2.066811e-12, -2.073536e-12, 
    -2.061975e-12, -2.09776e-12, -2.075661e-12, -2.042673e-12, -2.049447e-12, 
    -2.050414e-12, -2.04779e-12, -2.065596e-12, -2.059144e-12, -2.076521e-12, 
    -2.071825e-12, -2.07952e-12, -2.075696e-12, -2.075134e-12, -2.070223e-12, 
    -2.067165e-12, -2.05944e-12, -2.053155e-12, -2.04817e-12, -2.049329e-12, 
    -2.054805e-12, -2.064721e-12, -2.074101e-12, -2.072046e-12, 
    -2.078935e-12, -2.0607e-12, -2.068347e-12, -2.065391e-12, -2.073097e-12, 
    -2.056212e-12, -2.070592e-12, -2.052537e-12, -2.05412e-12, -2.059016e-12, 
    -2.068865e-12, -2.071044e-12, -2.073371e-12, -2.071935e-12, 
    -2.064972e-12, -2.063831e-12, -2.058897e-12, -2.057535e-12, 
    -2.053775e-12, -2.050663e-12, -2.053507e-12, -2.056493e-12, 
    -2.064975e-12, -2.072619e-12, -2.080952e-12, -2.082992e-12, 
    -2.092729e-12, -2.084803e-12, -2.097883e-12, -2.086763e-12, 
    -2.106012e-12, -2.071424e-12, -2.086435e-12, -2.059239e-12, 
    -2.062169e-12, -2.067468e-12, -2.079623e-12, -2.073061e-12, 
    -2.080735e-12, -2.063787e-12, -2.054994e-12, -2.052718e-12, 
    -2.048474e-12, -2.052815e-12, -2.052462e-12, -2.056617e-12, 
    -2.055282e-12, -2.065257e-12, -2.059898e-12, -2.07512e-12, -2.080674e-12, 
    -2.09636e-12, -2.105977e-12, -2.115765e-12, -2.120086e-12, -2.121401e-12, 
    -2.121951e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.367222e-15, 3.376314e-15, 3.374547e-15, 3.381874e-15, 3.377812e-15, 
    3.382607e-15, 3.369067e-15, 3.376673e-15, 3.371819e-15, 3.368042e-15, 
    3.39607e-15, 3.382201e-15, 3.410466e-15, 3.401636e-15, 3.423802e-15, 
    3.40909e-15, 3.426766e-15, 3.423381e-15, 3.433573e-15, 3.430655e-15, 
    3.443671e-15, 3.43492e-15, 3.450415e-15, 3.441583e-15, 3.442964e-15, 
    3.43463e-15, 3.384996e-15, 3.394344e-15, 3.384442e-15, 3.385776e-15, 
    3.385178e-15, 3.377895e-15, 3.37422e-15, 3.366528e-15, 3.367926e-15, 
    3.373576e-15, 3.386375e-15, 3.382034e-15, 3.392976e-15, 3.392729e-15, 
    3.404892e-15, 3.39941e-15, 3.419828e-15, 3.414032e-15, 3.430776e-15, 
    3.426567e-15, 3.430578e-15, 3.429363e-15, 3.430594e-15, 3.424421e-15, 
    3.427066e-15, 3.421633e-15, 3.400437e-15, 3.406671e-15, 3.388062e-15, 
    3.376849e-15, 3.3694e-15, 3.364109e-15, 3.364857e-15, 3.366283e-15, 
    3.373609e-15, 3.380494e-15, 3.385737e-15, 3.389241e-15, 3.392694e-15, 
    3.403127e-15, 3.40865e-15, 3.420999e-15, 3.418774e-15, 3.422544e-15, 
    3.426149e-15, 3.432193e-15, 3.431199e-15, 3.433861e-15, 3.422447e-15, 
    3.430033e-15, 3.417507e-15, 3.420933e-15, 3.393622e-15, 3.383206e-15, 
    3.378767e-15, 3.374887e-15, 3.365432e-15, 3.371962e-15, 3.369388e-15, 
    3.375512e-15, 3.3794e-15, 3.377477e-15, 3.389337e-15, 3.384728e-15, 
    3.408978e-15, 3.398541e-15, 3.425728e-15, 3.41923e-15, 3.427286e-15, 
    3.423177e-15, 3.430215e-15, 3.423881e-15, 3.434852e-15, 3.437237e-15, 
    3.435607e-15, 3.441872e-15, 3.423529e-15, 3.430577e-15, 3.377423e-15, 
    3.377737e-15, 3.379198e-15, 3.372772e-15, 3.37238e-15, 3.366489e-15, 
    3.371732e-15, 3.373962e-15, 3.379626e-15, 3.382972e-15, 3.386153e-15, 
    3.393142e-15, 3.400939e-15, 3.411834e-15, 3.419652e-15, 3.424889e-15, 
    3.421679e-15, 3.424513e-15, 3.421344e-15, 3.419859e-15, 3.436343e-15, 
    3.42709e-15, 3.440971e-15, 3.440204e-15, 3.433923e-15, 3.440291e-15, 
    3.377957e-15, 3.376153e-15, 3.369882e-15, 3.37479e-15, 3.365848e-15, 
    3.370853e-15, 3.373729e-15, 3.384822e-15, 3.38726e-15, 3.389517e-15, 
    3.393975e-15, 3.399691e-15, 3.409709e-15, 3.418415e-15, 3.426359e-15, 
    3.425777e-15, 3.425982e-15, 3.427755e-15, 3.423362e-15, 3.428476e-15, 
    3.429333e-15, 3.42709e-15, 3.440101e-15, 3.436386e-15, 3.440188e-15, 
    3.437769e-15, 3.376739e-15, 3.379775e-15, 3.378135e-15, 3.381219e-15, 
    3.379045e-15, 3.388703e-15, 3.391596e-15, 3.405125e-15, 3.399578e-15, 
    3.408407e-15, 3.400476e-15, 3.401881e-15, 3.408691e-15, 3.400905e-15, 
    3.417933e-15, 3.406389e-15, 3.427823e-15, 3.416305e-15, 3.428545e-15, 
    3.426325e-15, 3.430001e-15, 3.433291e-15, 3.43743e-15, 3.445059e-15, 
    3.443294e-15, 3.449672e-15, 3.3843e-15, 3.388233e-15, 3.387889e-15, 
    3.392005e-15, 3.395047e-15, 3.401639e-15, 3.4122e-15, 3.408231e-15, 
    3.415518e-15, 3.416979e-15, 3.405909e-15, 3.412706e-15, 3.390866e-15, 
    3.394396e-15, 3.392296e-15, 3.384609e-15, 3.409143e-15, 3.39656e-15, 
    3.419781e-15, 3.412977e-15, 3.432822e-15, 3.422955e-15, 3.442321e-15, 
    3.450581e-15, 3.458357e-15, 3.467423e-15, 3.390381e-15, 3.387709e-15, 
    3.392495e-15, 3.399107e-15, 3.405244e-15, 3.413392e-15, 3.414226e-15, 
    3.415751e-15, 3.4197e-15, 3.42302e-15, 3.416231e-15, 3.423852e-15, 
    3.395211e-15, 3.410235e-15, 3.386697e-15, 3.393789e-15, 3.398718e-15, 
    3.396558e-15, 3.407777e-15, 3.410419e-15, 3.421141e-15, 3.415602e-15, 
    3.448542e-15, 3.433983e-15, 3.474326e-15, 3.46307e-15, 3.386775e-15, 
    3.390373e-15, 3.40288e-15, 3.396932e-15, 3.413937e-15, 3.418114e-15, 
    3.421512e-15, 3.425851e-15, 3.42632e-15, 3.42889e-15, 3.424679e-15, 
    3.428725e-15, 3.413409e-15, 3.420256e-15, 3.401453e-15, 3.406033e-15, 
    3.403927e-15, 3.401615e-15, 3.408748e-15, 3.416338e-15, 3.416503e-15, 
    3.418933e-15, 3.425775e-15, 3.414005e-15, 3.450413e-15, 3.427941e-15, 
    3.394294e-15, 3.401213e-15, 3.402204e-15, 3.399524e-15, 3.417697e-15, 
    3.411117e-15, 3.428828e-15, 3.424045e-15, 3.431881e-15, 3.427988e-15, 
    3.427415e-15, 3.422412e-15, 3.419295e-15, 3.411418e-15, 3.405003e-15, 
    3.399913e-15, 3.401097e-15, 3.406687e-15, 3.416803e-15, 3.426362e-15, 
    3.424268e-15, 3.431286e-15, 3.412705e-15, 3.420498e-15, 3.417487e-15, 
    3.42534e-15, 3.408124e-15, 3.422777e-15, 3.404373e-15, 3.405989e-15, 
    3.410986e-15, 3.421025e-15, 3.423249e-15, 3.425618e-15, 3.424157e-15, 
    3.41706e-15, 3.415898e-15, 3.410865e-15, 3.409474e-15, 3.405638e-15, 
    3.402459e-15, 3.405363e-15, 3.40841e-15, 3.417064e-15, 3.424852e-15, 
    3.433338e-15, 3.435414e-15, 3.445307e-15, 3.43725e-15, 3.450537e-15, 
    3.439235e-15, 3.458793e-15, 3.42363e-15, 3.43891e-15, 3.411214e-15, 
    3.414203e-15, 3.419602e-15, 3.431981e-15, 3.425303e-15, 3.433114e-15, 
    3.415852e-15, 3.406878e-15, 3.404558e-15, 3.400222e-15, 3.404657e-15, 
    3.404297e-15, 3.408539e-15, 3.407176e-15, 3.417351e-15, 3.411887e-15, 
    3.4274e-15, 3.433053e-15, 3.449002e-15, 3.458762e-15, 3.46869e-15, 
    3.473068e-15, 3.4744e-15, 3.474956e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.758231e-09, -8.796739e-09, -8.789253e-09, -8.820313e-09, -8.803083e-09, 
    -8.823421e-09, -8.766038e-09, -8.798269e-09, -8.777693e-09, 
    -8.761697e-09, -8.88059e-09, -8.821698e-09, -8.941757e-09, -8.9042e-09, 
    -8.998543e-09, -8.935913e-09, -9.011171e-09, -8.996735e-09, 
    -9.040182e-09, -9.027735e-09, -9.083308e-09, -9.045927e-09, 
    -9.112114e-09, -9.07438e-09, -9.080283e-09, -9.044694e-09, -8.833549e-09, 
    -8.873259e-09, -8.831196e-09, -8.836859e-09, -8.834318e-09, 
    -8.803439e-09, -8.787879e-09, -8.755287e-09, -8.761203e-09, 
    -8.785142e-09, -8.839406e-09, -8.820985e-09, -8.867407e-09, 
    -8.866359e-09, -8.918041e-09, -8.894738e-09, -8.981602e-09, 
    -8.956914e-09, -9.028255e-09, -9.010313e-09, -9.027412e-09, 
    -9.022227e-09, -9.027479e-09, -9.001167e-09, -9.012441e-09, 
    -8.989287e-09, -8.899103e-09, -8.925608e-09, -8.846557e-09, 
    -8.799026e-09, -8.767452e-09, -8.745046e-09, -8.748215e-09, 
    -8.754252e-09, -8.785281e-09, -8.814453e-09, -8.836684e-09, 
    -8.851556e-09, -8.866208e-09, -8.910562e-09, -8.934035e-09, 
    -8.986595e-09, -8.977109e-09, -8.993178e-09, -9.008528e-09, 
    -9.034302e-09, -9.030059e-09, -9.041415e-09, -8.992753e-09, 
    -9.025094e-09, -8.971705e-09, -8.986308e-09, -8.870195e-09, 
    -8.825954e-09, -8.807152e-09, -8.790693e-09, -8.750649e-09, 
    -8.778303e-09, -8.767402e-09, -8.793335e-09, -8.809813e-09, 
    -8.801663e-09, -8.851963e-09, -8.832408e-09, -8.935427e-09, 
    -8.891053e-09, -9.006738e-09, -8.979056e-09, -9.013373e-09, 
    -8.995862e-09, -9.025867e-09, -8.998862e-09, -9.045641e-09, 
    -9.055827e-09, -9.048866e-09, -9.075604e-09, -8.997366e-09, 
    -9.027413e-09, -8.801435e-09, -8.802764e-09, -8.808956e-09, 
    -8.781736e-09, -8.780071e-09, -8.755125e-09, -8.777322e-09, 
    -8.786774e-09, -8.810768e-09, -8.824961e-09, -8.838453e-09, 
    -8.868117e-09, -8.901246e-09, -8.947571e-09, -8.98085e-09, -9.003158e-09, 
    -8.989478e-09, -9.001556e-09, -8.988056e-09, -8.981727e-09, 
    -9.052011e-09, -9.012546e-09, -9.071758e-09, -9.068482e-09, 
    -9.041685e-09, -9.068851e-09, -8.803697e-09, -8.796048e-09, 
    -8.769491e-09, -8.790274e-09, -8.752408e-09, -8.773604e-09, 
    -8.785793e-09, -8.832817e-09, -8.843148e-09, -8.852728e-09, 
    -8.871649e-09, -8.895931e-09, -8.938528e-09, -8.975589e-09, 
    -9.009422e-09, -9.006943e-09, -9.007815e-09, -9.015373e-09, 
    -8.996651e-09, -9.018447e-09, -9.022106e-09, -9.012541e-09, 
    -9.068043e-09, -9.052187e-09, -9.068412e-09, -9.058088e-09, 
    -8.798534e-09, -8.811405e-09, -8.804451e-09, -8.817529e-09, 
    -8.808315e-09, -8.849285e-09, -8.861567e-09, -8.919042e-09, 
    -8.895453e-09, -8.932994e-09, -8.899266e-09, -8.905243e-09, -8.93422e-09, 
    -8.901089e-09, -8.973546e-09, -8.924424e-09, -9.015667e-09, 
    -8.966615e-09, -9.018741e-09, -9.009275e-09, -9.024948e-09, 
    -9.038985e-09, -9.056643e-09, -9.089225e-09, -9.08168e-09, -9.108929e-09, 
    -8.830592e-09, -8.847286e-09, -8.845817e-09, -8.863286e-09, 
    -8.876206e-09, -8.904209e-09, -8.949121e-09, -8.932232e-09, 
    -8.963237e-09, -8.969462e-09, -8.922357e-09, -8.95128e-09, -8.858459e-09, 
    -8.873457e-09, -8.864526e-09, -8.831909e-09, -8.936125e-09, 
    -8.882642e-09, -8.981401e-09, -8.952427e-09, -9.036983e-09, 
    -8.994933e-09, -9.077527e-09, -9.112838e-09, -9.146065e-09, 
    -9.184901e-09, -8.856397e-09, -8.845054e-09, -8.865364e-09, 
    -8.893464e-09, -8.919534e-09, -8.954195e-09, -8.95774e-09, -8.964235e-09, 
    -8.981052e-09, -8.995194e-09, -8.966288e-09, -8.99874e-09, -8.876936e-09, 
    -8.940767e-09, -8.840765e-09, -8.87088e-09, -8.891807e-09, -8.882626e-09, 
    -8.930302e-09, -8.941538e-09, -8.987199e-09, -8.963595e-09, 
    -9.104123e-09, -9.04195e-09, -9.214468e-09, -9.166258e-09, -8.841091e-09, 
    -8.856357e-09, -8.909492e-09, -8.884211e-09, -8.956508e-09, 
    -8.974304e-09, -8.988771e-09, -9.007263e-09, -9.00926e-09, -9.020217e-09, 
    -9.002262e-09, -9.019508e-09, -8.954268e-09, -8.983422e-09, 
    -8.903418e-09, -8.922891e-09, -8.913932e-09, -8.904106e-09, 
    -8.934433e-09, -8.966744e-09, -8.967432e-09, -8.977793e-09, 
    -9.006991e-09, -8.956802e-09, -9.11215e-09, -9.016213e-09, -8.873005e-09, 
    -8.902413e-09, -8.906611e-09, -8.895221e-09, -8.972521e-09, 
    -8.944512e-09, -9.01995e-09, -8.999561e-09, -9.032967e-09, -9.016367e-09, 
    -9.013925e-09, -8.992605e-09, -8.979331e-09, -8.945796e-09, -8.91851e-09, 
    -8.896873e-09, -8.901903e-09, -8.925673e-09, -8.968719e-09, 
    -9.009441e-09, -9.000521e-09, -9.030428e-09, -8.951266e-09, 
    -8.984461e-09, -8.971631e-09, -9.005084e-09, -8.931783e-09, 
    -8.994206e-09, -8.915828e-09, -8.9227e-09, -8.943956e-09, -8.986714e-09, 
    -8.996171e-09, -9.006271e-09, -9.000039e-09, -8.969812e-09, 
    -8.964859e-09, -8.943439e-09, -8.937525e-09, -8.921203e-09, 
    -8.907691e-09, -8.920037e-09, -8.933003e-09, -8.969824e-09, 
    -9.003007e-09, -9.039185e-09, -9.048037e-09, -9.09031e-09, -9.0559e-09, 
    -9.112684e-09, -9.06441e-09, -9.147975e-09, -8.997822e-09, -9.062988e-09, 
    -8.944923e-09, -8.957642e-09, -8.980648e-09, -9.033413e-09, 
    -9.004927e-09, -9.038241e-09, -8.964665e-09, -8.926493e-09, 
    -8.916615e-09, -8.898188e-09, -8.917036e-09, -8.915503e-09, 
    -8.933539e-09, -8.927743e-09, -8.971047e-09, -8.947787e-09, 
    -9.013864e-09, -9.037977e-09, -9.106073e-09, -9.147819e-09, -9.19031e-09, 
    -9.20907e-09, -9.21478e-09, -9.217167e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.039262e-10, -1.043833e-10, -1.042944e-10, -1.046631e-10, -1.044586e-10, 
    -1.047e-10, -1.040189e-10, -1.044015e-10, -1.041572e-10, -1.039673e-10, 
    -1.053787e-10, -1.046796e-10, -1.061048e-10, -1.05659e-10, -1.067789e-10, 
    -1.060354e-10, -1.069288e-10, -1.067575e-10, -1.072732e-10, 
    -1.071255e-10, -1.077852e-10, -1.073414e-10, -1.081272e-10, 
    -1.076792e-10, -1.077493e-10, -1.073268e-10, -1.048203e-10, 
    -1.052917e-10, -1.047923e-10, -1.048596e-10, -1.048294e-10, 
    -1.044628e-10, -1.042781e-10, -1.038912e-10, -1.039615e-10, 
    -1.042456e-10, -1.048898e-10, -1.046711e-10, -1.052222e-10, 
    -1.052098e-10, -1.058233e-10, -1.055466e-10, -1.065778e-10, 
    -1.062847e-10, -1.071316e-10, -1.069187e-10, -1.071216e-10, 
    -1.070601e-10, -1.071224e-10, -1.068101e-10, -1.069439e-10, -1.06669e-10, 
    -1.055985e-10, -1.059131e-10, -1.049747e-10, -1.044104e-10, 
    -1.040356e-10, -1.037697e-10, -1.038073e-10, -1.03879e-10, -1.042473e-10, 
    -1.045936e-10, -1.048575e-10, -1.05034e-10, -1.05208e-10, -1.057345e-10, 
    -1.060131e-10, -1.066371e-10, -1.065245e-10, -1.067152e-10, 
    -1.068975e-10, -1.072034e-10, -1.071531e-10, -1.072879e-10, 
    -1.067102e-10, -1.070941e-10, -1.064603e-10, -1.066337e-10, 
    -1.052553e-10, -1.047301e-10, -1.045069e-10, -1.043115e-10, 
    -1.038362e-10, -1.041645e-10, -1.040351e-10, -1.043429e-10, 
    -1.045385e-10, -1.044418e-10, -1.050388e-10, -1.048067e-10, 
    -1.060297e-10, -1.055029e-10, -1.068762e-10, -1.065476e-10, -1.06955e-10, 
    -1.067471e-10, -1.071033e-10, -1.067827e-10, -1.07338e-10, -1.07459e-10, 
    -1.073763e-10, -1.076937e-10, -1.067649e-10, -1.071216e-10, -1.04439e-10, 
    -1.044548e-10, -1.045283e-10, -1.042052e-10, -1.041854e-10, 
    -1.038893e-10, -1.041528e-10, -1.04265e-10, -1.045498e-10, -1.047183e-10, 
    -1.048785e-10, -1.052306e-10, -1.056239e-10, -1.061738e-10, 
    -1.065689e-10, -1.068337e-10, -1.066713e-10, -1.068147e-10, 
    -1.066544e-10, -1.065793e-10, -1.074137e-10, -1.069452e-10, 
    -1.076481e-10, -1.076092e-10, -1.072911e-10, -1.076136e-10, 
    -1.044659e-10, -1.043751e-10, -1.040599e-10, -1.043066e-10, 
    -1.038571e-10, -1.041087e-10, -1.042534e-10, -1.048116e-10, 
    -1.049342e-10, -1.050479e-10, -1.052725e-10, -1.055608e-10, 
    -1.060665e-10, -1.065064e-10, -1.069081e-10, -1.068786e-10, -1.06889e-10, 
    -1.069787e-10, -1.067565e-10, -1.070152e-10, -1.070586e-10, 
    -1.069451e-10, -1.07604e-10, -1.074157e-10, -1.076084e-10, -1.074858e-10, 
    -1.044046e-10, -1.045574e-10, -1.044748e-10, -1.046301e-10, 
    -1.045207e-10, -1.050071e-10, -1.051529e-10, -1.058351e-10, 
    -1.055551e-10, -1.060008e-10, -1.056004e-10, -1.056713e-10, 
    -1.060153e-10, -1.05622e-10, -1.064822e-10, -1.05899e-10, -1.069822e-10, 
    -1.063999e-10, -1.070187e-10, -1.069063e-10, -1.070924e-10, -1.07259e-10, 
    -1.074686e-10, -1.078555e-10, -1.077659e-10, -1.080894e-10, 
    -1.047852e-10, -1.049833e-10, -1.049659e-10, -1.051733e-10, 
    -1.053266e-10, -1.056591e-10, -1.061922e-10, -1.059917e-10, 
    -1.063598e-10, -1.064337e-10, -1.058745e-10, -1.062178e-10, -1.05116e-10, 
    -1.05294e-10, -1.05188e-10, -1.048008e-10, -1.060379e-10, -1.05403e-10, 
    -1.065754e-10, -1.062315e-10, -1.072353e-10, -1.067361e-10, 
    -1.077166e-10, -1.081358e-10, -1.085303e-10, -1.089913e-10, 
    -1.050915e-10, -1.049568e-10, -1.051979e-10, -1.055315e-10, -1.05841e-10, 
    -1.062525e-10, -1.062945e-10, -1.063716e-10, -1.065713e-10, 
    -1.067392e-10, -1.06396e-10, -1.067813e-10, -1.053353e-10, -1.060931e-10, 
    -1.049059e-10, -1.052634e-10, -1.055118e-10, -1.054029e-10, 
    -1.059688e-10, -1.061022e-10, -1.066443e-10, -1.06364e-10, -1.080323e-10, 
    -1.072942e-10, -1.093423e-10, -1.0877e-10, -1.049098e-10, -1.05091e-10, 
    -1.057218e-10, -1.054217e-10, -1.062799e-10, -1.064912e-10, 
    -1.066629e-10, -1.068824e-10, -1.069061e-10, -1.070362e-10, 
    -1.068231e-10, -1.070278e-10, -1.062533e-10, -1.065994e-10, 
    -1.056497e-10, -1.058808e-10, -1.057745e-10, -1.056578e-10, 
    -1.060179e-10, -1.064014e-10, -1.064096e-10, -1.065326e-10, 
    -1.068792e-10, -1.062834e-10, -1.081276e-10, -1.069887e-10, 
    -1.052886e-10, -1.056377e-10, -1.056876e-10, -1.055524e-10, -1.0647e-10, 
    -1.061375e-10, -1.07033e-10, -1.06791e-10, -1.071876e-10, -1.069905e-10, 
    -1.069615e-10, -1.067084e-10, -1.065509e-10, -1.061528e-10, 
    -1.058288e-10, -1.05572e-10, -1.056317e-10, -1.059139e-10, -1.064249e-10, 
    -1.069083e-10, -1.068024e-10, -1.071574e-10, -1.062177e-10, 
    -1.066117e-10, -1.064595e-10, -1.068566e-10, -1.059864e-10, 
    -1.067274e-10, -1.05797e-10, -1.058786e-10, -1.061309e-10, -1.066385e-10, 
    -1.067508e-10, -1.068707e-10, -1.067967e-10, -1.064378e-10, 
    -1.063791e-10, -1.061248e-10, -1.060546e-10, -1.058608e-10, 
    -1.057004e-10, -1.05847e-10, -1.060009e-10, -1.06438e-10, -1.068319e-10, 
    -1.072614e-10, -1.073665e-10, -1.078683e-10, -1.074598e-10, -1.08134e-10, 
    -1.075609e-10, -1.085529e-10, -1.067704e-10, -1.07544e-10, -1.061424e-10, 
    -1.062934e-10, -1.065665e-10, -1.071929e-10, -1.068547e-10, 
    -1.072502e-10, -1.063767e-10, -1.059236e-10, -1.058063e-10, 
    -1.055876e-10, -1.058113e-10, -1.057931e-10, -1.060072e-10, 
    -1.059384e-10, -1.064525e-10, -1.061764e-10, -1.069608e-10, 
    -1.072471e-10, -1.080555e-10, -1.085511e-10, -1.090555e-10, 
    -1.092782e-10, -1.09346e-10, -1.093744e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.62019e-12, -8.658122e-12, -8.650748e-12, -8.681344e-12, -8.664371e-12, 
    -8.684406e-12, -8.62788e-12, -8.659629e-12, -8.639361e-12, -8.623604e-12, 
    -8.740719e-12, -8.682708e-12, -8.800973e-12, -8.763977e-12, 
    -8.856911e-12, -8.795216e-12, -8.869351e-12, -8.85513e-12, -8.897928e-12, 
    -8.885667e-12, -8.940411e-12, -8.903587e-12, -8.968787e-12, 
    -8.931616e-12, -8.937432e-12, -8.902373e-12, -8.694382e-12, 
    -8.733497e-12, -8.692064e-12, -8.697642e-12, -8.695139e-12, 
    -8.664722e-12, -8.649395e-12, -8.61729e-12, -8.623118e-12, -8.646698e-12, 
    -8.700151e-12, -8.682005e-12, -8.727734e-12, -8.726701e-12, 
    -8.777611e-12, -8.754657e-12, -8.840223e-12, -8.815904e-12, 
    -8.886179e-12, -8.868506e-12, -8.885349e-12, -8.880241e-12, 
    -8.885416e-12, -8.859496e-12, -8.870601e-12, -8.847792e-12, 
    -8.758956e-12, -8.785065e-12, -8.707196e-12, -8.660375e-12, 
    -8.629273e-12, -8.607203e-12, -8.610323e-12, -8.616271e-12, 
    -8.646836e-12, -8.675572e-12, -8.697471e-12, -8.71212e-12, -8.726552e-12, 
    -8.770244e-12, -8.793366e-12, -8.845141e-12, -8.835797e-12, 
    -8.851626e-12, -8.866748e-12, -8.892136e-12, -8.887957e-12, 
    -8.899143e-12, -8.851208e-12, -8.883066e-12, -8.830474e-12, 
    -8.844858e-12, -8.730481e-12, -8.6869e-12, -8.668379e-12, -8.652166e-12, 
    -8.612722e-12, -8.639961e-12, -8.629223e-12, -8.654769e-12, 
    -8.671001e-12, -8.662972e-12, -8.712519e-12, -8.693257e-12, 
    -8.794737e-12, -8.751026e-12, -8.864983e-12, -8.837714e-12, -8.87152e-12, 
    -8.854269e-12, -8.883827e-12, -8.857226e-12, -8.903305e-12, -8.91334e-12, 
    -8.906482e-12, -8.932821e-12, -8.85575e-12, -8.885349e-12, -8.662748e-12, 
    -8.664057e-12, -8.670157e-12, -8.643344e-12, -8.641704e-12, -8.61713e-12, 
    -8.638995e-12, -8.648306e-12, -8.671942e-12, -8.685923e-12, 
    -8.699212e-12, -8.728433e-12, -8.761067e-12, -8.806699e-12, 
    -8.839482e-12, -8.861457e-12, -8.847982e-12, -8.859879e-12, -8.84658e-12, 
    -8.840346e-12, -8.909581e-12, -8.870705e-12, -8.929033e-12, 
    -8.925805e-12, -8.899409e-12, -8.92617e-12, -8.664977e-12, -8.657441e-12, 
    -8.631281e-12, -8.651754e-12, -8.614454e-12, -8.635334e-12, 
    -8.647339e-12, -8.69366e-12, -8.703837e-12, -8.713274e-12, -8.731912e-12, 
    -8.755831e-12, -8.797791e-12, -8.8343e-12, -8.867627e-12, -8.865185e-12, 
    -8.866045e-12, -8.87349e-12, -8.855048e-12, -8.876518e-12, -8.880121e-12, 
    -8.870699e-12, -8.925373e-12, -8.909753e-12, -8.925737e-12, 
    -8.915567e-12, -8.659891e-12, -8.672569e-12, -8.665718e-12, 
    -8.678601e-12, -8.669525e-12, -8.709882e-12, -8.721981e-12, 
    -8.778597e-12, -8.755361e-12, -8.79234e-12, -8.759117e-12, -8.765004e-12, 
    -8.793548e-12, -8.760912e-12, -8.832287e-12, -8.783899e-12, 
    -8.873779e-12, -8.82546e-12, -8.876807e-12, -8.867483e-12, -8.882921e-12, 
    -8.896749e-12, -8.914143e-12, -8.94624e-12, -8.938807e-12, -8.965649e-12, 
    -8.691469e-12, -8.707914e-12, -8.706465e-12, -8.723675e-12, 
    -8.736401e-12, -8.763985e-12, -8.808228e-12, -8.79159e-12, -8.822132e-12, 
    -8.828264e-12, -8.781862e-12, -8.810353e-12, -8.718919e-12, 
    -8.733693e-12, -8.724896e-12, -8.692767e-12, -8.795425e-12, 
    -8.742741e-12, -8.840024e-12, -8.811484e-12, -8.894777e-12, 
    -8.853355e-12, -8.934716e-12, -8.9695e-12, -9.002232e-12, -9.040489e-12, 
    -8.716888e-12, -8.705714e-12, -8.725721e-12, -8.753401e-12, 
    -8.779082e-12, -8.813225e-12, -8.816718e-12, -8.823114e-12, 
    -8.839682e-12, -8.853612e-12, -8.825138e-12, -8.857104e-12, -8.73712e-12, 
    -8.799997e-12, -8.701491e-12, -8.731155e-12, -8.751769e-12, 
    -8.742725e-12, -8.789689e-12, -8.800757e-12, -8.845737e-12, 
    -8.822485e-12, -8.960915e-12, -8.89967e-12, -9.069615e-12, -9.022123e-12, 
    -8.70181e-12, -8.716849e-12, -8.769189e-12, -8.744286e-12, -8.815504e-12, 
    -8.833034e-12, -8.847284e-12, -8.865501e-12, -8.867468e-12, 
    -8.878261e-12, -8.860574e-12, -8.877562e-12, -8.813297e-12, 
    -8.842016e-12, -8.763206e-12, -8.782388e-12, -8.773563e-12, 
    -8.763884e-12, -8.793758e-12, -8.825586e-12, -8.826265e-12, 
    -8.836471e-12, -8.865232e-12, -8.815792e-12, -8.968822e-12, 
    -8.874317e-12, -8.733248e-12, -8.762217e-12, -8.766352e-12, 
    -8.755131e-12, -8.831277e-12, -8.803687e-12, -8.877998e-12, 
    -8.857914e-12, -8.890821e-12, -8.874469e-12, -8.872063e-12, 
    -8.851061e-12, -8.837986e-12, -8.804952e-12, -8.778073e-12, 
    -8.756758e-12, -8.761714e-12, -8.785128e-12, -8.827532e-12, 
    -8.867646e-12, -8.858859e-12, -8.88832e-12, -8.81034e-12, -8.843039e-12, 
    -8.830402e-12, -8.863354e-12, -8.791148e-12, -8.852639e-12, 
    -8.775431e-12, -8.7822e-12, -8.803139e-12, -8.845258e-12, -8.854574e-12, 
    -8.864524e-12, -8.858385e-12, -8.828609e-12, -8.82373e-12, -8.80263e-12, 
    -8.796804e-12, -8.780726e-12, -8.767416e-12, -8.779578e-12, -8.79235e-12, 
    -8.828621e-12, -8.861308e-12, -8.896946e-12, -8.905666e-12, 
    -8.947308e-12, -8.913412e-12, -8.969349e-12, -8.921794e-12, 
    -9.004113e-12, -8.8562e-12, -8.920393e-12, -8.804091e-12, -8.816621e-12, 
    -8.839283e-12, -8.89126e-12, -8.863198e-12, -8.896016e-12, -8.823539e-12, 
    -8.785936e-12, -8.776206e-12, -8.758054e-12, -8.776622e-12, 
    -8.775112e-12, -8.792878e-12, -8.787169e-12, -8.829825e-12, 
    -8.806912e-12, -8.872003e-12, -8.895757e-12, -8.962837e-12, 
    -9.003959e-12, -9.045817e-12, -9.064297e-12, -9.069922e-12, -9.072273e-12 ;

 SMIN_NH4 =
  0.0004618175, 0.0004637462, 0.0004633711, 0.0004649268, 0.0004640637, 
    0.0004650823, 0.0004622081, 0.0004638225, 0.0004627918, 0.0004619905, 
    0.0004679451, 0.0004649957, 0.0004710071, 0.0004691266, 0.0004738494, 
    0.0004707145, 0.0004744813, 0.0004737586, 0.0004759328, 0.0004753099, 
    0.000478091, 0.0004762202, 0.000479532, 0.000477644, 0.0004779394, 
    0.0004761582, 0.0004655895, 0.0004675784, 0.0004654716, 0.0004657552, 
    0.0004656278, 0.0004640814, 0.0004633022, 0.0004616693, 0.0004619657, 
    0.0004631648, 0.0004658824, 0.0004649597, 0.0004672842, 0.0004672317, 
    0.0004698193, 0.0004686527, 0.0004730011, 0.0004717651, 0.0004753358, 
    0.0004744379, 0.0004752936, 0.000475034, 0.0004752968, 0.0004739799, 
    0.0004745441, 0.0004733852, 0.0004688718, 0.0004701988, 0.0004662407, 
    0.0004638605, 0.0004622788, 0.0004611565, 0.000461315, 0.0004616175, 
    0.0004631717, 0.0004646325, 0.0004657458, 0.0004664904, 0.000467224, 
    0.0004694453, 0.0004706201, 0.000473251, 0.000472776, 0.0004735803, 
    0.0004743485, 0.0004756383, 0.0004754259, 0.0004759941, 0.0004735587, 
    0.0004751774, 0.000472505, 0.000473236, 0.0004674249, 0.0004652088, 
    0.0004642674, 0.0004634428, 0.000461437, 0.0004628222, 0.0004622761, 
    0.0004635748, 0.0004644001, 0.0004639918, 0.0004665107, 0.0004655314, 
    0.0004706897, 0.0004684681, 0.000474259, 0.0004728733, 0.0004745908, 
    0.0004737144, 0.0004752161, 0.0004738645, 0.0004762055, 0.0004767153, 
    0.0004763668, 0.0004777047, 0.0004737892, 0.0004752931, 0.0004639807, 
    0.0004640473, 0.0004643573, 0.0004629941, 0.0004629106, 0.0004616609, 
    0.0004627727, 0.0004632462, 0.0004644477, 0.0004651585, 0.0004658341, 
    0.0004673195, 0.0004689783, 0.0004712974, 0.0004729631, 0.0004740795, 
    0.0004733948, 0.0004739992, 0.0004733235, 0.0004730066, 0.0004765242, 
    0.0004745492, 0.0004775121, 0.0004773482, 0.0004760073, 0.0004773665, 
    0.0004640939, 0.0004637107, 0.0004623806, 0.0004634215, 0.0004615247, 
    0.0004625865, 0.000463197, 0.000465552, 0.0004660691, 0.0004665489, 
    0.0004674962, 0.000468712, 0.0004708446, 0.0004726997, 0.0004743929, 
    0.0004742687, 0.0004743124, 0.0004746906, 0.0004737536, 0.0004748444, 
    0.0004750274, 0.0004745487, 0.000477326, 0.0004765326, 0.0004773445, 
    0.0004768277, 0.0004638352, 0.0004644797, 0.0004641313, 0.0004647864, 
    0.0004643248, 0.0004663767, 0.0004669917, 0.0004698693, 0.0004686881, 
    0.0004705676, 0.0004688788, 0.0004691781, 0.0004706291, 0.0004689699, 
    0.0004725974, 0.0004701384, 0.0004747053, 0.0004722504, 0.000474859, 
    0.0004743851, 0.0004751694, 0.000475872, 0.0004767555, 0.000478386, 
    0.0004780083, 0.0004793716, 0.0004654405, 0.0004662766, 0.0004662028, 
    0.0004670775, 0.0004677244, 0.0004691264, 0.0004713749, 0.0004705293, 
    0.0004720812, 0.0004723929, 0.0004700347, 0.0004714827, 0.0004668354, 
    0.0004675864, 0.0004671391, 0.0004655058, 0.0004707239, 0.0004680461, 
    0.00047299, 0.0004715396, 0.0004757717, 0.0004736673, 0.0004778004, 
    0.0004795674, 0.0004812293, 0.0004831721, 0.0004667326, 0.0004661645, 
    0.0004671814, 0.0004685886, 0.0004698936, 0.0004716288, 0.0004718061, 
    0.0004721311, 0.0004729729, 0.0004736807, 0.0004722339, 0.000473858, 
    0.0004677609, 0.0004709562, 0.0004659491, 0.0004674573, 0.0004685048, 
    0.0004680451, 0.0004704319, 0.0004709943, 0.00047328, 0.0004720984, 
    0.0004791313, 0.0004760202, 0.0004846506, 0.0004822394, 0.000465966, 
    0.0004667304, 0.0004693909, 0.000468125, 0.0004717444, 0.0004726352, 
    0.0004733591, 0.0004742848, 0.0004743845, 0.000474933, 0.0004740342, 
    0.0004748973, 0.0004716319, 0.0004730912, 0.000469086, 0.0004700609, 
    0.0004696123, 0.0004691203, 0.0004706385, 0.0004722561, 0.0004722904, 
    0.000472809, 0.000474271, 0.000471758, 0.000479533, 0.0004747322, 
    0.0004675639, 0.0004690365, 0.0004692464, 0.0004686761, 0.0004725457, 
    0.0004711438, 0.0004749196, 0.000473899, 0.0004755708, 0.0004747401, 
    0.0004746178, 0.0004735507, 0.0004728863, 0.0004712077, 0.0004698415, 
    0.0004687581, 0.0004690099, 0.0004702, 0.0004723548, 0.000474393, 
    0.0004739465, 0.0004754431, 0.0004714808, 0.0004731425, 0.0004725003, 
    0.0004741745, 0.0004705066, 0.0004736319, 0.0004697077, 0.0004700517, 
    0.0004711158, 0.0004732563, 0.0004737292, 0.0004742349, 0.0004739227, 
    0.0004724099, 0.0004721619, 0.0004710895, 0.0004707935, 0.0004699763, 
    0.0004692996, 0.0004699178, 0.0004705669, 0.00047241, 0.0004740709, 
    0.0004758813, 0.0004763242, 0.0004784398, 0.0004767179, 0.0004795595, 
    0.0004771441, 0.0004813247, 0.0004738124, 0.0004770737, 0.0004711641, 
    0.0004718007, 0.0004729525, 0.0004755933, 0.0004741673, 0.0004758348, 
    0.0004721521, 0.0004702413, 0.0004697465, 0.0004688239, 0.0004697675, 
    0.0004696907, 0.0004705936, 0.0004703033, 0.0004724711, 0.0004713066, 
    0.0004746141, 0.0004758209, 0.0004792282, 0.0004813166, 0.0004834418, 
    0.00048438, 0.0004846655, 0.0004847849 ;

 SMIN_NH4_vr =
  0.00302471, 0.003029867, 0.003028857, 0.003033014, 0.003030704, 
    0.003033421, 0.003025739, 0.003030051, 0.003027294, 0.003025146, 
    0.003041045, 0.003033175, 0.003049191, 0.00304418, 0.003056736, 
    0.003048406, 0.00305841, 0.003056486, 0.003062254, 0.003060597, 
    0.003067966, 0.003063007, 0.003071773, 0.003066776, 0.003067555, 
    0.003062829, 0.00303478, 0.00304009, 0.003034459, 0.003035217, 
    0.003034873, 0.00303074, 0.003028658, 0.003024285, 0.003025074, 
    0.003028281, 0.003035535, 0.003033067, 0.003039265, 0.003039125, 
    0.003046013, 0.003042907, 0.003054471, 0.003051181, 0.003060662, 
    0.003058275, 0.003060544, 0.003059851, 0.003060544, 0.003057051, 
    0.003058542, 0.003055465, 0.003043526, 0.003047054, 0.003036506, 
    0.003030149, 0.003025915, 0.003022914, 0.003023331, 0.003024142, 
    0.003028294, 0.003032191, 0.003035162, 0.003037144, 0.003039096, 
    0.003045018, 0.00304814, 0.003055128, 0.003053864, 0.003055997, 
    0.003058034, 0.003061452, 0.003060887, 0.00306239, 0.003055923, 
    0.003060221, 0.003053118, 0.003055061, 0.003039666, 0.003033745, 
    0.003031233, 0.003029023, 0.003023656, 0.003027362, 0.003025898, 
    0.003029364, 0.003031567, 0.003030472, 0.003037194, 0.003034577, 
    0.00304832, 0.003042405, 0.003057801, 0.003054116, 0.003058673, 
    0.003056347, 0.003060326, 0.003056739, 0.003062944, 0.003064297, 
    0.003063366, 0.003066912, 0.003056521, 0.003060514, 0.00303046, 
    0.003030638, 0.003031463, 0.003027817, 0.003027592, 0.003024245, 
    0.003027214, 0.003028481, 0.003031686, 0.00303358, 0.003035379, 
    0.003039342, 0.003043759, 0.003049926, 0.003054351, 0.003057311, 
    0.003055492, 0.003057092, 0.003055297, 0.00305445, 0.003063782, 
    0.003058544, 0.003066393, 0.003065959, 0.003062402, 0.003065999, 
    0.003030757, 0.003029728, 0.003026173, 0.00302895, 0.003023874, 
    0.003026715, 0.003028344, 0.003034629, 0.003036004, 0.003037285, 
    0.003039807, 0.003043042, 0.003048718, 0.003053645, 0.00305814, 
    0.003057806, 0.00305792, 0.00305892, 0.003056431, 0.003059322, 
    0.003059804, 0.003058534, 0.003065892, 0.00306379, 0.003065938, 
    0.003064564, 0.003030058, 0.003031775, 0.00303084, 0.003032591, 
    0.003031352, 0.00303683, 0.003038467, 0.003046129, 0.003042978, 
    0.003047983, 0.00304348, 0.003044278, 0.003048139, 0.003043715, 
    0.003053365, 0.003046822, 0.003058956, 0.003052434, 0.003059358, 
    0.003058095, 0.003060172, 0.003062037, 0.003064372, 0.003068693, 
    0.003067686, 0.003071295, 0.003034337, 0.003036564, 0.003036365, 
    0.003038693, 0.003040414, 0.00304415, 0.00305013, 0.003047875, 
    0.003051999, 0.003052828, 0.003046549, 0.003050403, 0.003038024, 
    0.003040022, 0.003038827, 0.003034466, 0.00304837, 0.003041236, 
    0.003054387, 0.003050528, 0.003061762, 0.003056179, 0.003067133, 
    0.003071813, 0.003076201, 0.00308133, 0.003037776, 0.003036256, 
    0.003038964, 0.003042717, 0.003046184, 0.003050801, 0.003051268, 
    0.003052128, 0.00305436, 0.003056241, 0.003052395, 0.003056703, 
    0.003040486, 0.003048987, 0.003035643, 0.003039667, 0.003042451, 
    0.003041226, 0.003047577, 0.003049069, 0.003055142, 0.003052002, 
    0.003070651, 0.00306241, 0.003085223, 0.003078862, 0.003035723, 
    0.003037757, 0.003044844, 0.003041473, 0.003051099, 0.003053468, 
    0.003055384, 0.003057844, 0.003058101, 0.003059558, 0.003057165, 
    0.003059457, 0.003050777, 0.003054656, 0.003043998, 0.00304659, 
    0.003045394, 0.003044079, 0.003048117, 0.003052421, 0.003052506, 
    0.003053881, 0.003057767, 0.003051081, 0.003071706, 0.00305898, 
    0.003039976, 0.003043897, 0.003044451, 0.003042932, 0.003053222, 
    0.003049495, 0.003059522, 0.003056808, 0.003061241, 0.003059037, 
    0.003058706, 0.003055874, 0.003054103, 0.003049642, 0.003046, 
    0.003043115, 0.003043779, 0.003046949, 0.003052674, 0.003058088, 
    0.003056899, 0.003060865, 0.003050338, 0.003054756, 0.003053043, 
    0.003057489, 0.003047803, 0.003056116, 0.003045673, 0.003046584, 
    0.003049412, 0.003055104, 0.003056351, 0.003057695, 0.003056859, 
    0.003052842, 0.003052179, 0.003049322, 0.003048531, 0.003046357, 
    0.003044549, 0.003046196, 0.003047917, 0.003052818, 0.003057227, 
    0.003062025, 0.003063198, 0.003068802, 0.003064238, 0.003071762, 
    0.003065365, 0.003076421, 0.003056585, 0.003065236, 0.003049541, 
    0.003051229, 0.00305429, 0.003061296, 0.003057507, 0.003061933, 
    0.00305215, 0.003047065, 0.003045742, 0.003043287, 0.003045792, 
    0.003045589, 0.003047988, 0.003047211, 0.003052972, 0.003049877, 
    0.003058658, 0.003061861, 0.003070882, 0.003076401, 0.00308201, 
    0.003084481, 0.003085232, 0.003085543,
  0.00181022, 0.001816974, 0.001815661, 0.001821105, 0.001818086, 0.00182165, 
    0.00181159, 0.001817243, 0.001813634, 0.001810828, 0.001831657, 
    0.001821348, 0.001842343, 0.001835782, 0.001852247, 0.001841323, 
    0.001854447, 0.001851931, 0.001859498, 0.001857331, 0.001867001, 
    0.001860497, 0.001872005, 0.001865448, 0.001866474, 0.001860283, 
    0.001823423, 0.001830375, 0.001823011, 0.001824003, 0.001823558, 
    0.001818148, 0.001815422, 0.001809703, 0.001810741, 0.001814941, 
    0.001824449, 0.001821222, 0.001829349, 0.001829165, 0.0018382, 
    0.001834128, 0.001849293, 0.001844987, 0.001857421, 0.001854297, 
    0.001857275, 0.001856372, 0.001857287, 0.001852703, 0.001854668, 
    0.001850633, 0.001834891, 0.001839522, 0.001825701, 0.001817376, 
    0.001811838, 0.001807906, 0.001808462, 0.001809522, 0.001814965, 
    0.001820078, 0.001823972, 0.001826575, 0.001829139, 0.001836895, 
    0.001840994, 0.001850164, 0.001848509, 0.001851311, 0.001853986, 
    0.001858474, 0.001857736, 0.001859713, 0.001851237, 0.001856872, 
    0.001847567, 0.001850113, 0.001829839, 0.001822093, 0.0018188, 
    0.001815914, 0.00180889, 0.001813742, 0.001811829, 0.001816377, 
    0.001819265, 0.001817837, 0.001826646, 0.001823223, 0.001841237, 
    0.001833484, 0.001853674, 0.001848849, 0.00185483, 0.001851778, 
    0.001857006, 0.001852301, 0.001860448, 0.001862221, 0.001861009, 
    0.00186566, 0.001852041, 0.001857275, 0.001817797, 0.00181803, 
    0.001819115, 0.001814344, 0.001814052, 0.001809675, 0.001813569, 
    0.001815227, 0.001819432, 0.001821919, 0.001824281, 0.001829473, 
    0.001835266, 0.001843357, 0.001849162, 0.00185305, 0.001850666, 
    0.001852771, 0.001850418, 0.001849314, 0.001861557, 0.001854686, 
    0.001864991, 0.001864421, 0.00185976, 0.001864486, 0.001818193, 
    0.001816852, 0.001812196, 0.00181584, 0.001809198, 0.001812917, 
    0.001815055, 0.001823295, 0.001825103, 0.00182678, 0.001830091, 
    0.001834337, 0.001841778, 0.001848245, 0.001854141, 0.001853709, 
    0.001853861, 0.001855178, 0.001851916, 0.001855714, 0.001856351, 
    0.001854685, 0.001864345, 0.001861587, 0.001864409, 0.001862613, 
    0.001817288, 0.001819544, 0.001818325, 0.001820617, 0.001819003, 
    0.001826178, 0.001828328, 0.001838376, 0.001834253, 0.001840812, 
    0.00183492, 0.001835964, 0.001841028, 0.001835238, 0.001847889, 
    0.001839316, 0.001855229, 0.001846681, 0.001855765, 0.001854116, 
    0.001856845, 0.001859289, 0.001862362, 0.001868028, 0.001866717, 
    0.001871451, 0.001822905, 0.001825828, 0.00182557, 0.001828628, 
    0.001830888, 0.001835783, 0.001843627, 0.001840679, 0.00184609, 
    0.001847176, 0.001838954, 0.001844004, 0.001827783, 0.001830408, 
    0.001828845, 0.001823136, 0.001841359, 0.001832014, 0.001849258, 
    0.001844204, 0.001858941, 0.001851617, 0.001865995, 0.001872131, 
    0.001877898, 0.001884633, 0.001827422, 0.001825437, 0.001828991, 
    0.001833906, 0.001838461, 0.001844512, 0.001845131, 0.001846264, 
    0.001849197, 0.001851662, 0.001846623, 0.00185228, 0.001831018, 
    0.001842169, 0.001824687, 0.001829957, 0.001833616, 0.001832011, 
    0.001840341, 0.001842303, 0.001850269, 0.001846152, 0.001870618, 
    0.001859807, 0.001889753, 0.001881401, 0.001824743, 0.001827415, 
    0.001836707, 0.001832288, 0.001844916, 0.00184802, 0.001850542, 
    0.001853766, 0.001854113, 0.001856022, 0.001852894, 0.001855898, 
    0.001844525, 0.00184961, 0.001835645, 0.001839047, 0.001837482, 
    0.001835765, 0.001841063, 0.001846702, 0.001846822, 0.001848629, 
    0.001853721, 0.001844967, 0.001872014, 0.001855327, 0.001830328, 
    0.001835471, 0.001836203, 0.001834212, 0.001847709, 0.001842822, 
    0.001855975, 0.001852423, 0.001858242, 0.001855351, 0.001854926, 
    0.001851211, 0.001848897, 0.001843047, 0.001838282, 0.001834501, 
    0.00183538, 0.001839533, 0.001847047, 0.001854145, 0.001852591, 
    0.0018578, 0.001844001, 0.001849792, 0.001847555, 0.001853386, 0.0018406, 
    0.001851493, 0.001837813, 0.001839014, 0.001842725, 0.001850185, 
    0.001851832, 0.001853593, 0.001852506, 0.001847237, 0.001846373, 
    0.001842635, 0.001841603, 0.001838752, 0.001836392, 0.001838549, 
    0.001840814, 0.001847239, 0.001853024, 0.001859325, 0.001860865, 
    0.001868218, 0.001862234, 0.001872107, 0.001863717, 0.001878231, 
    0.001852122, 0.001863468, 0.001842894, 0.001845114, 0.001849127, 
    0.001858321, 0.001853358, 0.001859161, 0.001846339, 0.001839677, 
    0.001837951, 0.001834731, 0.001838024, 0.001837757, 0.001840907, 
    0.001839894, 0.001847452, 0.001843394, 0.001854916, 0.001859115, 
    0.001870956, 0.001878203, 0.001885568, 0.001888818, 0.001889806, 
    0.001890219,
  0.001646094, 0.001653298, 0.001651898, 0.001657706, 0.001654484, 
    0.001658287, 0.001647554, 0.001653584, 0.001649735, 0.001646742, 
    0.001668967, 0.001657964, 0.001680378, 0.001673372, 0.00169096, 
    0.001679289, 0.001693311, 0.001690623, 0.00169871, 0.001696394, 
    0.001706732, 0.001699779, 0.001712085, 0.001705072, 0.00170617, 
    0.00169955, 0.001660179, 0.001667598, 0.001659739, 0.001660798, 
    0.001660323, 0.001654551, 0.001651641, 0.001645542, 0.00164665, 
    0.001651129, 0.001661274, 0.001657831, 0.001666504, 0.001666308, 
    0.001675955, 0.001671606, 0.001687804, 0.001683203, 0.001696491, 
    0.001693151, 0.001696334, 0.001695369, 0.001696347, 0.001691448, 
    0.001693547, 0.001689235, 0.001672421, 0.001677366, 0.00166261, 
    0.001653726, 0.001647819, 0.001643626, 0.001644219, 0.001645349, 
    0.001651155, 0.00165661, 0.001660765, 0.001663543, 0.00166628, 
    0.00167456, 0.001678938, 0.001688735, 0.001686967, 0.001689961, 
    0.001692819, 0.001697617, 0.001696827, 0.00169894, 0.001689881, 
    0.001695903, 0.00168596, 0.001688681, 0.001667026, 0.00165876, 
    0.001655246, 0.001652167, 0.001644675, 0.001649849, 0.00164781, 
    0.001652661, 0.001655742, 0.001654218, 0.001663619, 0.001659966, 
    0.001679198, 0.001670919, 0.001692486, 0.001687329, 0.001693721, 
    0.00169046, 0.001696047, 0.001691019, 0.001699726, 0.001701621, 
    0.001700326, 0.001705299, 0.00169074, 0.001696334, 0.001654176, 
    0.001654424, 0.001655582, 0.001650492, 0.00165018, 0.001645512, 
    0.001649666, 0.001651434, 0.001655921, 0.001658574, 0.001661095, 
    0.001666637, 0.001672821, 0.001681462, 0.001687664, 0.001691819, 
    0.001689271, 0.00169152, 0.001689006, 0.001687827, 0.001700912, 
    0.001693567, 0.001704584, 0.001703975, 0.00169899, 0.001704043, 
    0.001654599, 0.001653168, 0.001648201, 0.001652089, 0.001645004, 
    0.00164897, 0.001651251, 0.001660043, 0.001661972, 0.001663762, 
    0.001667296, 0.001671829, 0.001679776, 0.001686684, 0.001692985, 
    0.001692523, 0.001692686, 0.001694093, 0.001690607, 0.001694666, 
    0.001695347, 0.001693566, 0.001703893, 0.001700944, 0.001703962, 
    0.001702041, 0.001653633, 0.00165604, 0.00165474, 0.001657185, 
    0.001655462, 0.00166312, 0.001665414, 0.001676142, 0.00167174, 
    0.001678744, 0.001672452, 0.001673567, 0.001678973, 0.001672791, 
    0.001686304, 0.001677146, 0.001694148, 0.001685012, 0.00169472, 
    0.001692958, 0.001695875, 0.001698488, 0.001701773, 0.001707832, 
    0.001706429, 0.001711493, 0.001659626, 0.001662746, 0.001662471, 
    0.001665734, 0.001668147, 0.001673374, 0.001681751, 0.001678601, 
    0.001684382, 0.001685542, 0.00167676, 0.001682153, 0.001664833, 
    0.001667634, 0.001665966, 0.001659873, 0.001679328, 0.001669349, 
    0.001687766, 0.001682367, 0.001698115, 0.001690288, 0.001705657, 
    0.00171222, 0.001718389, 0.001725596, 0.001664448, 0.001662328, 
    0.001666122, 0.001671369, 0.001676233, 0.001682697, 0.001683357, 
    0.001684568, 0.001687702, 0.001690336, 0.001684951, 0.001690996, 
    0.001668284, 0.001680193, 0.001661528, 0.001667153, 0.00167106, 
    0.001669346, 0.001678241, 0.001680337, 0.001688847, 0.001684448, 
    0.001710601, 0.00169904, 0.001731078, 0.001722138, 0.001661588, 
    0.00166444, 0.00167436, 0.001669641, 0.001683128, 0.001686444, 
    0.001689139, 0.001692584, 0.001692955, 0.001694995, 0.001691652, 
    0.001694863, 0.00168271, 0.001688143, 0.001673226, 0.001676859, 
    0.001675188, 0.001673354, 0.001679012, 0.001685036, 0.001685164, 
    0.001687094, 0.001692535, 0.001683182, 0.001712093, 0.001694251, 
    0.001667549, 0.001673039, 0.001673822, 0.001671696, 0.001686112, 
    0.001680891, 0.001694945, 0.001691149, 0.001697368, 0.001694278, 
    0.001693824, 0.001689853, 0.001687381, 0.001681131, 0.001676042, 
    0.001672004, 0.001672943, 0.001677378, 0.001685404, 0.001692989, 
    0.001691328, 0.001696895, 0.00168215, 0.001688337, 0.001685946, 
    0.001692177, 0.001678518, 0.001690154, 0.001675542, 0.001676823, 
    0.001680788, 0.001688757, 0.001690518, 0.001692399, 0.001691238, 
    0.001685607, 0.001684684, 0.001680691, 0.001679589, 0.001676544, 
    0.001674023, 0.001676327, 0.001678745, 0.001685609, 0.001691791, 
    0.001698525, 0.001700172, 0.001708034, 0.001701636, 0.001712193, 
    0.00170322, 0.001718745, 0.001690826, 0.001702954, 0.001680968, 
    0.001683339, 0.001687627, 0.001697452, 0.001692148, 0.00169835, 
    0.001684648, 0.001677532, 0.001675688, 0.00167225, 0.001675767, 
    0.001675481, 0.001678845, 0.001677764, 0.001685837, 0.001681502, 
    0.001693812, 0.001698301, 0.001710962, 0.001718715, 0.001726599, 
    0.001730077, 0.001731135, 0.001731578,
  0.001514893, 0.001522024, 0.001520637, 0.001526388, 0.001523198, 
    0.001526964, 0.001516338, 0.001522307, 0.001518497, 0.001515534, 
    0.001537545, 0.001526645, 0.00154886, 0.001541913, 0.001559361, 
    0.00154778, 0.001561695, 0.001559026, 0.001567057, 0.001564757, 
    0.001575027, 0.001568119, 0.001580348, 0.001573377, 0.001574468, 
    0.001567891, 0.001528838, 0.001536189, 0.001528403, 0.001529451, 
    0.00152898, 0.001523264, 0.001520383, 0.001514347, 0.001515443, 
    0.001519876, 0.001529922, 0.001526512, 0.001535104, 0.00153491, 
    0.001544473, 0.001540162, 0.001556228, 0.001551663, 0.001564853, 
    0.001561536, 0.001564697, 0.001563739, 0.001564709, 0.001559846, 
    0.00156193, 0.001557649, 0.001540969, 0.001545873, 0.001531246, 
    0.001522448, 0.0015166, 0.001512451, 0.001513037, 0.001514156, 
    0.001519902, 0.001525303, 0.001529418, 0.001532171, 0.001534882, 
    0.00154309, 0.001547432, 0.001557152, 0.001555397, 0.001558369, 
    0.001561206, 0.00156597, 0.001565186, 0.001567285, 0.00155829, 
    0.001564269, 0.001554398, 0.001557098, 0.001535622, 0.001527432, 
    0.001523952, 0.001520904, 0.001513488, 0.00151861, 0.001516591, 
    0.001521393, 0.001524444, 0.001522935, 0.001532246, 0.001528627, 
    0.001547689, 0.00153948, 0.001560875, 0.001555757, 0.001562102, 
    0.001558865, 0.001564412, 0.001559419, 0.001568066, 0.001569949, 
    0.001568662, 0.001573603, 0.001559143, 0.001564697, 0.001522893, 
    0.001523139, 0.001524285, 0.001519246, 0.001518937, 0.001514317, 
    0.001518428, 0.001520178, 0.001524621, 0.001527248, 0.001529746, 
    0.001535236, 0.001541366, 0.001549935, 0.001556089, 0.001560214, 
    0.001557685, 0.001559917, 0.001557421, 0.001556251, 0.001569243, 
    0.001561949, 0.001572892, 0.001572287, 0.001567335, 0.001572355, 
    0.001523312, 0.001521895, 0.001516978, 0.001520826, 0.001513814, 
    0.00151774, 0.001519997, 0.001528703, 0.001530615, 0.001532388, 
    0.001535889, 0.001540383, 0.001548263, 0.001555117, 0.001561371, 
    0.001560913, 0.001561074, 0.001562472, 0.001559011, 0.00156304, 
    0.001563716, 0.001561948, 0.001572206, 0.001569276, 0.001572274, 
    0.001570366, 0.001522356, 0.001524739, 0.001523451, 0.001525873, 
    0.001524167, 0.001531751, 0.001534024, 0.001544659, 0.001540294, 
    0.001547239, 0.001541, 0.001542105, 0.001547467, 0.001541337, 
    0.001554739, 0.001545654, 0.001562526, 0.001553458, 0.001563094, 
    0.001561344, 0.001564241, 0.001566836, 0.001570099, 0.00157612, 
    0.001574725, 0.001579759, 0.001528291, 0.001531381, 0.001531108, 
    0.001534342, 0.001536733, 0.001541914, 0.001550222, 0.001547098, 
    0.001552832, 0.001553983, 0.001545271, 0.001550621, 0.001533449, 
    0.001536224, 0.001534571, 0.001528535, 0.001547819, 0.001537924, 
    0.001556191, 0.001550833, 0.001566466, 0.001558693, 0.001573958, 
    0.001580482, 0.001586618, 0.001593788, 0.001533067, 0.001530967, 
    0.001534726, 0.001539927, 0.001544749, 0.00155116, 0.001551816, 
    0.001553017, 0.001556127, 0.001558741, 0.001553397, 0.001559397, 
    0.001536869, 0.001548677, 0.001530174, 0.001535748, 0.00153962, 
    0.001537921, 0.001546741, 0.001548819, 0.001557264, 0.001552898, 
    0.001578872, 0.001567384, 0.001599245, 0.001590346, 0.001530234, 
    0.001533059, 0.001542892, 0.001538214, 0.001551588, 0.001554879, 
    0.001557554, 0.001560973, 0.001561342, 0.001563367, 0.001560048, 
    0.001563236, 0.001551174, 0.001556565, 0.001541768, 0.00154537, 
    0.001543713, 0.001541895, 0.001547505, 0.001553481, 0.001553608, 
    0.001555524, 0.001560924, 0.001551642, 0.001580356, 0.001562629, 
    0.00153614, 0.001541582, 0.001542359, 0.001540251, 0.001554549, 
    0.001549369, 0.001563318, 0.001559549, 0.001565724, 0.001562655, 
    0.001562204, 0.001558263, 0.001555808, 0.001549607, 0.00154456, 
    0.001540557, 0.001541487, 0.001545885, 0.001553847, 0.001561375, 
    0.001559726, 0.001565254, 0.001550618, 0.001556757, 0.001554385, 
    0.00156057, 0.001547015, 0.00155856, 0.001544063, 0.001545335, 
    0.001549267, 0.001557174, 0.001558922, 0.001560789, 0.001559637, 
    0.001554048, 0.001553132, 0.001549171, 0.001548077, 0.001545058, 
    0.001542558, 0.001544842, 0.001547241, 0.00155405, 0.001560186, 
    0.001566873, 0.001568509, 0.001576321, 0.001569963, 0.001580455, 
    0.001571536, 0.001586972, 0.001559228, 0.001571273, 0.001549445, 
    0.001551797, 0.001556052, 0.001565807, 0.001560541, 0.001566699, 
    0.001553096, 0.001546037, 0.001544209, 0.0015408, 0.001544287, 
    0.001544003, 0.00154734, 0.001546268, 0.001554277, 0.001549975, 
    0.001562193, 0.00156665, 0.001579232, 0.001586942, 0.001594786, 
    0.001598249, 0.001599302, 0.001599743,
  0.0013795, 0.001385892, 0.001384649, 0.001389807, 0.001386945, 0.001390323, 
    0.001380795, 0.001386146, 0.00138273, 0.001380075, 0.001399825, 
    0.001390037, 0.001409999, 0.00140375, 0.001419454, 0.001409026, 
    0.001421557, 0.001419152, 0.001426391, 0.001424317, 0.001433584, 
    0.001427349, 0.00143839, 0.001432094, 0.001433079, 0.001427144, 
    0.001392005, 0.001398606, 0.001391615, 0.001392556, 0.001392133, 
    0.001387005, 0.001384421, 0.001379011, 0.001379993, 0.001383967, 
    0.001392979, 0.001389918, 0.001397632, 0.001397458, 0.001406052, 
    0.001402176, 0.001416632, 0.001412521, 0.001424404, 0.001421414, 
    0.001424263, 0.001423399, 0.001424274, 0.00141989, 0.001421768, 
    0.001417911, 0.001402902, 0.001407311, 0.001394167, 0.001386272, 
    0.00138103, 0.001377312, 0.001377838, 0.00137884, 0.00138399, 
    0.001388833, 0.001392526, 0.001394997, 0.001397433, 0.001404809, 
    0.001408714, 0.001417463, 0.001415883, 0.00141856, 0.001421117, 
    0.001425412, 0.001424704, 0.001426597, 0.001418489, 0.001423877, 
    0.001414983, 0.001417415, 0.001398097, 0.001390744, 0.001387622, 
    0.001384888, 0.001378242, 0.001382831, 0.001381022, 0.001385326, 
    0.001388063, 0.001386709, 0.001395065, 0.001391816, 0.001408945, 
    0.001401564, 0.001420818, 0.001416207, 0.001421924, 0.001419006, 
    0.001424006, 0.001419506, 0.001427302, 0.001429, 0.001427839, 
    0.001432298, 0.001419257, 0.001424263, 0.001386671, 0.001386892, 
    0.00138792, 0.001383401, 0.001383125, 0.001378985, 0.001382668, 
    0.001384238, 0.001388221, 0.001390579, 0.00139282, 0.00139775, 
    0.001403259, 0.001410966, 0.001416506, 0.001420222, 0.001417943, 
    0.001419955, 0.001417706, 0.001416652, 0.001428364, 0.001421786, 
    0.001431657, 0.00143111, 0.001426642, 0.001431172, 0.001387047, 
    0.001385777, 0.001381369, 0.001384818, 0.001378534, 0.001382051, 
    0.001384075, 0.001391884, 0.0013936, 0.001395192, 0.001398337, 
    0.001402374, 0.001409461, 0.00141563, 0.001421265, 0.001420852, 
    0.001420998, 0.001422257, 0.001419138, 0.001422769, 0.001423379, 
    0.001421785, 0.001431037, 0.001428393, 0.001431098, 0.001429377, 
    0.00138619, 0.001388327, 0.001387172, 0.001389344, 0.001387814, 
    0.00139462, 0.001396662, 0.001406219, 0.001402295, 0.00140854, 
    0.001402929, 0.001403923, 0.001408745, 0.001403232, 0.001415291, 
    0.001407115, 0.001422306, 0.001414137, 0.001422818, 0.001421241, 
    0.001423852, 0.001426192, 0.001429136, 0.001434571, 0.001433312, 
    0.001437858, 0.001391514, 0.001394288, 0.001394044, 0.001396947, 
    0.001399095, 0.001403751, 0.001411224, 0.001408413, 0.001413573, 
    0.00141461, 0.00140677, 0.001411583, 0.001396145, 0.001398638, 
    0.001397153, 0.001391733, 0.001409061, 0.001400165, 0.001416598, 
    0.001411774, 0.001425858, 0.001418852, 0.001432619, 0.001438511, 
    0.001444058, 0.001450546, 0.001395802, 0.001393917, 0.001397292, 
    0.001401965, 0.0014063, 0.001412068, 0.001412658, 0.00141374, 0.00141654, 
    0.001418895, 0.001414082, 0.001419486, 0.001399217, 0.001409834, 
    0.001393205, 0.00139821, 0.001401689, 0.001400162, 0.001408092, 
    0.001409962, 0.001417564, 0.001413633, 0.001437057, 0.001426687, 
    0.001455488, 0.001447431, 0.001393258, 0.001395795, 0.00140463, 
    0.001400425, 0.001412453, 0.001415416, 0.001417825, 0.001420906, 
    0.001421238, 0.001423064, 0.001420072, 0.001422946, 0.001412081, 
    0.001416935, 0.001403619, 0.001406859, 0.001405368, 0.001403734, 
    0.001408779, 0.001414158, 0.001414272, 0.001415997, 0.001420862, 
    0.001412502, 0.001438398, 0.001422399, 0.001398562, 0.001403453, 
    0.001404151, 0.001402256, 0.001415119, 0.001410457, 0.00142302, 
    0.001419623, 0.001425189, 0.001422423, 0.001422016, 0.001418464, 
    0.001416253, 0.001410671, 0.00140613, 0.001402531, 0.001403367, 
    0.001407322, 0.001414487, 0.001421269, 0.001419783, 0.001424766, 
    0.001411581, 0.001417108, 0.001414971, 0.001420543, 0.001408338, 
    0.001418732, 0.001405684, 0.001406827, 0.001410364, 0.001417483, 
    0.001419058, 0.001420741, 0.001419702, 0.001414668, 0.001413844, 
    0.001410278, 0.001409294, 0.001406578, 0.00140433, 0.001406384, 
    0.001408542, 0.00141467, 0.001420197, 0.001426225, 0.001427701, 
    0.001434752, 0.001429013, 0.001438487, 0.001430433, 0.001444378, 
    0.001419334, 0.001430195, 0.001410525, 0.001412642, 0.001416473, 
    0.001425264, 0.001420516, 0.001426069, 0.001413811, 0.001407459, 
    0.001405815, 0.00140275, 0.001405885, 0.00140563, 0.00140863, 
    0.001407666, 0.001414874, 0.001411001, 0.001422006, 0.001426024, 
    0.001437382, 0.001444351, 0.001451449, 0.001454585, 0.001455539, 
    0.001455938,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.348949e-06, 1.360497e-06, 1.358248e-06, 1.367592e-06, 1.362404e-06, 
    1.368528e-06, 1.351285e-06, 1.360956e-06, 1.354778e-06, 1.349985e-06, 
    1.385818e-06, 1.368008e-06, 1.404436e-06, 1.392987e-06, 1.421834e-06, 
    1.402651e-06, 1.425718e-06, 1.421277e-06, 1.43466e-06, 1.430819e-06, 
    1.448008e-06, 1.436434e-06, 1.456957e-06, 1.445238e-06, 1.447069e-06, 
    1.436052e-06, 1.371582e-06, 1.383595e-06, 1.370872e-06, 1.372582e-06, 
    1.371814e-06, 1.362511e-06, 1.357835e-06, 1.348066e-06, 1.349837e-06, 
    1.357012e-06, 1.37335e-06, 1.367792e-06, 1.381818e-06, 1.3815e-06, 
    1.3972e-06, 1.39011e-06, 1.416631e-06, 1.409067e-06, 1.430979e-06, 
    1.425452e-06, 1.430719e-06, 1.429121e-06, 1.43074e-06, 1.422638e-06, 
    1.426106e-06, 1.418988e-06, 1.391438e-06, 1.399507e-06, 1.375511e-06, 
    1.361184e-06, 1.351708e-06, 1.345005e-06, 1.345951e-06, 1.347757e-06, 
    1.357054e-06, 1.365824e-06, 1.372527e-06, 1.37702e-06, 1.381454e-06, 
    1.394924e-06, 1.402077e-06, 1.418163e-06, 1.415252e-06, 1.420184e-06, 
    1.424903e-06, 1.432844e-06, 1.431535e-06, 1.43504e-06, 1.420052e-06, 
    1.430004e-06, 1.413594e-06, 1.418073e-06, 1.382666e-06, 1.36929e-06, 
    1.363628e-06, 1.358679e-06, 1.346679e-06, 1.35496e-06, 1.351693e-06, 
    1.359472e-06, 1.364427e-06, 1.361975e-06, 1.377143e-06, 1.371236e-06, 
    1.402501e-06, 1.38899e-06, 1.424352e-06, 1.415849e-06, 1.426394e-06, 
    1.421008e-06, 1.430242e-06, 1.42193e-06, 1.436344e-06, 1.439493e-06, 
    1.437341e-06, 1.445616e-06, 1.421469e-06, 1.430718e-06, 1.361907e-06, 
    1.362307e-06, 1.36417e-06, 1.35599e-06, 1.35549e-06, 1.348017e-06, 
    1.354665e-06, 1.357502e-06, 1.364714e-06, 1.36899e-06, 1.37306e-06, 
    1.382032e-06, 1.392088e-06, 1.40621e-06, 1.416399e-06, 1.42325e-06, 
    1.419047e-06, 1.422757e-06, 1.41861e-06, 1.416667e-06, 1.438313e-06, 
    1.426138e-06, 1.444424e-06, 1.443409e-06, 1.435122e-06, 1.443523e-06, 
    1.362587e-06, 1.360287e-06, 1.352318e-06, 1.358552e-06, 1.347204e-06, 
    1.353551e-06, 1.357207e-06, 1.37136e-06, 1.374478e-06, 1.377374e-06, 
    1.383102e-06, 1.390471e-06, 1.403447e-06, 1.414786e-06, 1.425177e-06, 
    1.424414e-06, 1.424682e-06, 1.427009e-06, 1.42125e-06, 1.427955e-06, 
    1.429082e-06, 1.426136e-06, 1.443273e-06, 1.438366e-06, 1.443387e-06, 
    1.440191e-06, 1.361034e-06, 1.364906e-06, 1.362813e-06, 1.36675e-06, 
    1.363976e-06, 1.376334e-06, 1.38005e-06, 1.397504e-06, 1.390326e-06, 
    1.401758e-06, 1.391485e-06, 1.393302e-06, 1.402133e-06, 1.392038e-06, 
    1.41416e-06, 1.399144e-06, 1.427099e-06, 1.412036e-06, 1.428045e-06, 
    1.425131e-06, 1.429957e-06, 1.434288e-06, 1.439744e-06, 1.449841e-06, 
    1.447499e-06, 1.455963e-06, 1.370688e-06, 1.375729e-06, 1.375284e-06, 
    1.380569e-06, 1.384484e-06, 1.392988e-06, 1.406683e-06, 1.401525e-06, 
    1.411001e-06, 1.412907e-06, 1.398513e-06, 1.407343e-06, 1.379107e-06, 
    1.38365e-06, 1.380943e-06, 1.371084e-06, 1.402712e-06, 1.386435e-06, 
    1.416566e-06, 1.407692e-06, 1.433669e-06, 1.420721e-06, 1.446211e-06, 
    1.45718e-06, 1.467538e-06, 1.479694e-06, 1.378484e-06, 1.375054e-06, 
    1.381197e-06, 1.389722e-06, 1.397653e-06, 1.408234e-06, 1.409319e-06, 
    1.411306e-06, 1.41646e-06, 1.420802e-06, 1.411935e-06, 1.421891e-06, 
    1.384706e-06, 1.404129e-06, 1.373757e-06, 1.382868e-06, 1.389217e-06, 
    1.386429e-06, 1.400934e-06, 1.404364e-06, 1.418346e-06, 1.411108e-06, 
    1.454469e-06, 1.435203e-06, 1.488981e-06, 1.473852e-06, 1.373856e-06, 
    1.378471e-06, 1.394595e-06, 1.386911e-06, 1.408941e-06, 1.414391e-06, 
    1.418829e-06, 1.424513e-06, 1.425126e-06, 1.4285e-06, 1.422973e-06, 
    1.428281e-06, 1.408255e-06, 1.417187e-06, 1.392745e-06, 1.398674e-06, 
    1.395945e-06, 1.392954e-06, 1.402194e-06, 1.412073e-06, 1.412283e-06, 
    1.415459e-06, 1.42443e-06, 1.409028e-06, 1.456967e-06, 1.427267e-06, 
    1.383512e-06, 1.392442e-06, 1.393718e-06, 1.390254e-06, 1.413844e-06, 
    1.405273e-06, 1.428418e-06, 1.422143e-06, 1.43243e-06, 1.427314e-06, 
    1.426562e-06, 1.420005e-06, 1.415931e-06, 1.405665e-06, 1.397339e-06, 
    1.390755e-06, 1.392284e-06, 1.399522e-06, 1.412678e-06, 1.425181e-06, 
    1.422437e-06, 1.431646e-06, 1.407335e-06, 1.417504e-06, 1.413569e-06, 
    1.423839e-06, 1.401387e-06, 1.420501e-06, 1.396523e-06, 1.398617e-06, 
    1.405103e-06, 1.418198e-06, 1.421101e-06, 1.424207e-06, 1.42229e-06, 
    1.413014e-06, 1.411496e-06, 1.404944e-06, 1.403138e-06, 1.398159e-06, 
    1.394044e-06, 1.397804e-06, 1.401757e-06, 1.413016e-06, 1.423201e-06, 
    1.434348e-06, 1.437082e-06, 1.450177e-06, 1.439514e-06, 1.457133e-06, 
    1.442149e-06, 1.468135e-06, 1.42161e-06, 1.44171e-06, 1.405398e-06, 
    1.409287e-06, 1.416336e-06, 1.432569e-06, 1.423792e-06, 1.434059e-06, 
    1.411437e-06, 1.399773e-06, 1.396761e-06, 1.391154e-06, 1.396889e-06, 
    1.396422e-06, 1.401921e-06, 1.400152e-06, 1.41339e-06, 1.406271e-06, 
    1.426541e-06, 1.433975e-06, 1.455073e-06, 1.468085e-06, 1.481388e-06, 
    1.487281e-06, 1.489077e-06, 1.489828e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.308049e-06, 8.344628e-06, 8.337494e-06, 8.367022e-06, 8.350627e-06, 
    8.369953e-06, 8.315417e-06, 8.34603e-06, 8.326471e-06, 8.311266e-06, 
    8.424324e-06, 8.368273e-06, 8.482571e-06, 8.446762e-06, 8.536712e-06, 
    8.476982e-06, 8.548755e-06, 8.534956e-06, 8.576433e-06, 8.564532e-06, 
    8.617637e-06, 8.581898e-06, 8.645161e-06, 8.609079e-06, 8.614716e-06, 
    8.580681e-06, 8.379595e-06, 8.417405e-06, 8.377342e-06, 8.382733e-06, 
    8.380302e-06, 8.350934e-06, 8.336152e-06, 8.305174e-06, 8.310782e-06, 
    8.333524e-06, 8.385096e-06, 8.36756e-06, 8.411709e-06, 8.410713e-06, 
    8.459914e-06, 8.437717e-06, 8.520507e-06, 8.496943e-06, 8.565019e-06, 
    8.547877e-06, 8.5642e-06, 8.559235e-06, 8.56424e-06, 8.539122e-06, 
    8.549866e-06, 8.527767e-06, 8.441973e-06, 8.467213e-06, 8.39194e-06, 
    8.346746e-06, 8.316728e-06, 8.295457e-06, 8.298445e-06, 8.304181e-06, 
    8.33364e-06, 8.361345e-06, 8.38248e-06, 8.396614e-06, 8.410546e-06, 
    8.452802e-06, 8.475149e-06, 8.525257e-06, 8.516196e-06, 8.531521e-06, 
    8.546163e-06, 8.570762e-06, 8.566705e-06, 8.577541e-06, 8.531067e-06, 
    8.561946e-06, 8.510967e-06, 8.524903e-06, 8.414453e-06, 8.372322e-06, 
    8.354458e-06, 8.338793e-06, 8.300753e-06, 8.327015e-06, 8.316651e-06, 
    8.341267e-06, 8.356926e-06, 8.349165e-06, 8.396992e-06, 8.378379e-06, 
    8.476462e-06, 8.434185e-06, 8.544466e-06, 8.518035e-06, 8.550775e-06, 
    8.534061e-06, 8.562692e-06, 8.536908e-06, 8.581559e-06, 8.591297e-06, 
    8.584626e-06, 8.610177e-06, 8.53543e-06, 8.56412e-06, 8.348997e-06, 
    8.350263e-06, 8.356136e-06, 8.330265e-06, 8.328678e-06, 8.304973e-06, 
    8.32604e-06, 8.335024e-06, 8.357809e-06, 8.371293e-06, 8.384113e-06, 
    8.41234e-06, 8.443877e-06, 8.488008e-06, 8.519738e-06, 8.541012e-06, 
    8.527953e-06, 8.539466e-06, 8.526579e-06, 8.520527e-06, 8.587627e-06, 
    8.549936e-06, 8.606477e-06, 8.603347e-06, 8.577736e-06, 8.603676e-06, 
    8.351133e-06, 8.34385e-06, 8.318621e-06, 8.338348e-06, 8.302377e-06, 
    8.322509e-06, 8.334078e-06, 8.378764e-06, 8.388572e-06, 8.39769e-06, 
    8.415684e-06, 8.438791e-06, 8.479376e-06, 8.514704e-06, 8.546981e-06, 
    8.544602e-06, 8.545431e-06, 8.552636e-06, 8.534761e-06, 8.555555e-06, 
    8.559039e-06, 8.549906e-06, 8.602904e-06, 8.587753e-06, 8.603248e-06, 
    8.593367e-06, 8.346203e-06, 8.358425e-06, 8.351803e-06, 8.364239e-06, 
    8.355463e-06, 8.394431e-06, 8.406109e-06, 8.460825e-06, 8.438337e-06, 
    8.474108e-06, 8.441951e-06, 8.447648e-06, 8.475263e-06, 8.443663e-06, 
    8.512736e-06, 8.465892e-06, 8.552908e-06, 8.506102e-06, 8.555826e-06, 
    8.546774e-06, 8.561727e-06, 8.575137e-06, 8.591987e-06, 8.623139e-06, 
    8.615904e-06, 8.641962e-06, 8.376658e-06, 8.39253e-06, 8.391121e-06, 
    8.407733e-06, 8.420021e-06, 8.446686e-06, 8.489478e-06, 8.473363e-06, 
    8.502911e-06, 8.508852e-06, 8.463923e-06, 8.4915e-06, 8.403074e-06, 
    8.417342e-06, 8.408831e-06, 8.37779e-06, 8.477014e-06, 8.426053e-06, 
    8.520165e-06, 8.492519e-06, 8.573203e-06, 8.533062e-06, 8.611928e-06, 
    8.645708e-06, 8.677477e-06, 8.714662e-06, 8.401185e-06, 8.390377e-06, 
    8.409692e-06, 8.436456e-06, 8.461264e-06, 8.494304e-06, 8.497671e-06, 
    8.503853e-06, 8.519883e-06, 8.53338e-06, 8.505798e-06, 8.536738e-06, 
    8.420657e-06, 8.481434e-06, 8.386195e-06, 8.41486e-06, 8.434759e-06, 
    8.426016e-06, 8.471415e-06, 8.482113e-06, 8.525657e-06, 8.503135e-06, 
    8.63735e-06, 8.577918e-06, 8.742964e-06, 8.696789e-06, 8.386599e-06, 
    8.40111e-06, 8.451694e-06, 8.427615e-06, 8.496483e-06, 8.51346e-06, 
    8.52724e-06, 8.544897e-06, 8.546781e-06, 8.557246e-06, 8.540083e-06, 
    8.55655e-06, 8.494286e-06, 8.522093e-06, 8.445811e-06, 8.464354e-06, 
    8.455811e-06, 8.446438e-06, 8.475323e-06, 8.506142e-06, 8.506779e-06, 
    8.516653e-06, 8.544542e-06, 8.49661e-06, 8.645014e-06, 8.553312e-06, 
    8.416945e-06, 8.444945e-06, 8.448925e-06, 8.438074e-06, 8.511734e-06, 
    8.485027e-06, 8.556989e-06, 8.537511e-06, 8.569396e-06, 8.553547e-06, 
    8.551197e-06, 8.530847e-06, 8.518166e-06, 8.486189e-06, 8.460164e-06, 
    8.43955e-06, 8.444324e-06, 8.466975e-06, 8.508001e-06, 8.546856e-06, 
    8.538333e-06, 8.566867e-06, 8.491317e-06, 8.522984e-06, 8.510729e-06, 
    8.542645e-06, 8.472903e-06, 8.532465e-06, 8.457687e-06, 8.464222e-06, 
    8.484473e-06, 8.525264e-06, 8.53426e-06, 8.543906e-06, 8.537934e-06, 
    8.509102e-06, 8.504365e-06, 8.483925e-06, 8.478281e-06, 8.462722e-06, 
    8.449831e-06, 8.461597e-06, 8.473939e-06, 8.509045e-06, 8.540698e-06, 
    8.575229e-06, 8.583678e-06, 8.624089e-06, 8.59119e-06, 8.645486e-06, 
    8.599327e-06, 8.679227e-06, 8.535879e-06, 8.598119e-06, 8.485394e-06, 
    8.497508e-06, 8.519459e-06, 8.569817e-06, 8.542595e-06, 8.574417e-06, 
    8.504173e-06, 8.467776e-06, 8.458343e-06, 8.440793e-06, 8.458728e-06, 
    8.457269e-06, 8.474445e-06, 8.468908e-06, 8.510187e-06, 8.488005e-06, 
    8.551032e-06, 8.574065e-06, 8.639139e-06, 8.679073e-06, 8.719749e-06, 
    8.737708e-06, 8.743176e-06, 8.745455e-06,
  4.946846e-06, 4.984e-06, 4.976769e-06, 5.006795e-06, 4.990129e-06, 
    5.009803e-06, 4.954369e-06, 4.985479e-06, 4.96561e-06, 4.950185e-06, 
    5.065255e-06, 5.008135e-06, 5.124812e-06, 5.088208e-06, 5.180328e-06, 
    5.119112e-06, 5.192701e-06, 5.178554e-06, 5.221163e-06, 5.208944e-06, 
    5.263584e-06, 5.226806e-06, 5.291979e-06, 5.25479e-06, 5.260604e-06, 
    5.225595e-06, 5.019608e-06, 5.058133e-06, 5.01733e-06, 5.022816e-06, 
    5.020353e-06, 4.990475e-06, 4.975445e-06, 4.944008e-06, 4.949709e-06, 
    4.9728e-06, 5.025283e-06, 5.007443e-06, 5.052441e-06, 5.051423e-06, 
    5.101685e-06, 5.079001e-06, 5.16374e-06, 5.139605e-06, 5.209453e-06, 
    5.191857e-06, 5.208627e-06, 5.203539e-06, 5.208693e-06, 5.182895e-06, 
    5.193943e-06, 5.17126e-06, 5.083248e-06, 5.109061e-06, 5.032215e-06, 
    4.986213e-06, 4.955733e-06, 4.934148e-06, 4.937197e-06, 4.943013e-06, 
    4.972935e-06, 5.001124e-06, 5.022644e-06, 5.03706e-06, 5.051277e-06, 
    5.094407e-06, 5.117279e-06, 5.168628e-06, 5.159344e-06, 5.175072e-06, 
    5.190107e-06, 5.21539e-06, 5.211225e-06, 5.222375e-06, 5.174654e-06, 
    5.206354e-06, 5.15406e-06, 5.168345e-06, 5.055158e-06, 5.012253e-06, 
    4.994068e-06, 4.978159e-06, 4.939543e-06, 4.9662e-06, 4.955685e-06, 
    4.98071e-06, 4.996636e-06, 4.988756e-06, 5.037454e-06, 5.018502e-06, 
    5.118636e-06, 5.075419e-06, 5.188353e-06, 5.161249e-06, 5.194856e-06, 
    5.177697e-06, 5.207112e-06, 5.180636e-06, 5.226526e-06, 5.236539e-06, 
    5.229696e-06, 5.255994e-06, 5.17917e-06, 5.208628e-06, 4.988536e-06, 
    4.989821e-06, 4.995807e-06, 4.969514e-06, 4.967906e-06, 4.943853e-06, 
    4.965252e-06, 4.974376e-06, 4.997559e-06, 5.011292e-06, 5.024358e-06, 
    5.053131e-06, 5.085335e-06, 5.130484e-06, 5.163005e-06, 5.184845e-06, 
    5.171447e-06, 5.183274e-06, 5.170054e-06, 5.163862e-06, 5.232787e-06, 
    5.194046e-06, 5.252208e-06, 5.248984e-06, 5.222641e-06, 5.249347e-06, 
    4.990723e-06, 4.983331e-06, 4.9577e-06, 4.977754e-06, 4.941236e-06, 
    4.961667e-06, 4.973429e-06, 5.018901e-06, 5.028908e-06, 5.038198e-06, 
    5.05656e-06, 5.080162e-06, 5.121659e-06, 5.15786e-06, 5.190982e-06, 
    5.188553e-06, 5.189408e-06, 5.196818e-06, 5.178471e-06, 5.199832e-06, 
    5.203422e-06, 5.194041e-06, 5.248552e-06, 5.232958e-06, 5.248915e-06, 
    5.238759e-06, 4.985733e-06, 4.998175e-06, 4.991451e-06, 5.004099e-06, 
    4.995188e-06, 5.03486e-06, 5.046777e-06, 5.102664e-06, 5.079698e-06, 
    5.116261e-06, 5.083406e-06, 5.089224e-06, 5.117462e-06, 5.085179e-06, 
    5.155864e-06, 5.10791e-06, 5.197106e-06, 5.14909e-06, 5.200121e-06, 
    5.190839e-06, 5.206208e-06, 5.219988e-06, 5.237339e-06, 5.26941e-06, 
    5.261977e-06, 5.288834e-06, 5.016744e-06, 5.032922e-06, 5.031494e-06, 
    5.048441e-06, 5.060987e-06, 5.088215e-06, 5.131997e-06, 5.115517e-06, 
    5.145783e-06, 5.151867e-06, 5.10589e-06, 5.134104e-06, 5.043757e-06, 
    5.058318e-06, 5.049645e-06, 5.018021e-06, 5.119316e-06, 5.067243e-06, 
    5.163543e-06, 5.135224e-06, 5.218023e-06, 5.176791e-06, 5.257888e-06, 
    5.292695e-06, 5.325513e-06, 5.363966e-06, 5.041756e-06, 5.030755e-06, 
    5.050457e-06, 5.077764e-06, 5.103141e-06, 5.136951e-06, 5.140413e-06, 
    5.146758e-06, 5.163202e-06, 5.177044e-06, 5.148767e-06, 5.180515e-06, 
    5.061703e-06, 5.123844e-06, 5.0266e-06, 5.055817e-06, 5.076152e-06, 
    5.067226e-06, 5.113634e-06, 5.124594e-06, 5.169219e-06, 5.146132e-06, 
    5.284099e-06, 5.222904e-06, 5.393298e-06, 5.345496e-06, 5.026914e-06, 
    5.041717e-06, 5.09336e-06, 5.068765e-06, 5.139209e-06, 5.156602e-06, 
    5.170754e-06, 5.188869e-06, 5.190824e-06, 5.201568e-06, 5.183966e-06, 
    5.200872e-06, 5.137023e-06, 5.165521e-06, 5.087445e-06, 5.106411e-06, 
    5.097682e-06, 5.088115e-06, 5.117663e-06, 5.149212e-06, 5.149883e-06, 
    5.160015e-06, 5.188611e-06, 5.139495e-06, 5.292024e-06, 5.197651e-06, 
    5.057877e-06, 5.086471e-06, 5.090555e-06, 5.079469e-06, 5.154858e-06, 
    5.127497e-06, 5.201306e-06, 5.181321e-06, 5.214079e-06, 5.197792e-06, 
    5.195398e-06, 5.174508e-06, 5.161519e-06, 5.128751e-06, 5.102143e-06, 
    5.081076e-06, 5.085972e-06, 5.109123e-06, 5.151143e-06, 5.191003e-06, 
    5.182263e-06, 5.211587e-06, 5.134089e-06, 5.166539e-06, 5.15399e-06, 
    5.186731e-06, 5.11508e-06, 5.176087e-06, 5.099529e-06, 5.106224e-06, 
    5.126954e-06, 5.168745e-06, 5.178e-06, 5.187897e-06, 5.181788e-06, 
    5.152211e-06, 5.147369e-06, 5.126449e-06, 5.120681e-06, 5.104765e-06, 
    5.091605e-06, 5.10363e-06, 5.11627e-06, 5.152222e-06, 5.184698e-06, 
    5.220185e-06, 5.22888e-06, 5.270484e-06, 5.236614e-06, 5.292552e-06, 
    5.24499e-06, 5.327409e-06, 5.179623e-06, 5.243585e-06, 5.127897e-06, 
    5.140316e-06, 5.16281e-06, 5.214521e-06, 5.186577e-06, 5.219261e-06, 
    5.147179e-06, 5.109924e-06, 5.100296e-06, 5.082356e-06, 5.100706e-06, 
    5.099213e-06, 5.116791e-06, 5.11114e-06, 5.153417e-06, 5.130692e-06, 
    5.195339e-06, 5.219001e-06, 5.286019e-06, 5.32725e-06, 5.369324e-06, 
    5.387936e-06, 5.393605e-06, 5.395976e-06,
  4.461328e-06, 4.500614e-06, 4.492965e-06, 4.524734e-06, 4.507098e-06, 
    4.527918e-06, 4.469281e-06, 4.502177e-06, 4.481165e-06, 4.464858e-06, 
    4.586655e-06, 4.526153e-06, 4.649839e-06, 4.610998e-06, 4.708818e-06, 
    4.643787e-06, 4.721975e-06, 4.706934e-06, 4.752256e-06, 4.739254e-06, 
    4.797421e-06, 4.758261e-06, 4.827682e-06, 4.788056e-06, 4.794248e-06, 
    4.756972e-06, 4.538299e-06, 4.579105e-06, 4.535887e-06, 4.541695e-06, 
    4.539088e-06, 4.507463e-06, 4.491563e-06, 4.45833e-06, 4.464356e-06, 
    4.488767e-06, 4.544308e-06, 4.525421e-06, 4.573079e-06, 4.572e-06, 
    4.625295e-06, 4.601234e-06, 4.691189e-06, 4.665549e-06, 4.739796e-06, 
    4.721079e-06, 4.738917e-06, 4.733504e-06, 4.738987e-06, 4.711549e-06, 
    4.723297e-06, 4.699181e-06, 4.605737e-06, 4.633121e-06, 4.551649e-06, 
    4.502952e-06, 4.470722e-06, 4.447911e-06, 4.451133e-06, 4.457278e-06, 
    4.48891e-06, 4.518733e-06, 4.541515e-06, 4.556782e-06, 4.571845e-06, 
    4.617571e-06, 4.641842e-06, 4.696382e-06, 4.686518e-06, 4.703232e-06, 
    4.719218e-06, 4.746112e-06, 4.741681e-06, 4.753545e-06, 4.702789e-06, 
    4.736498e-06, 4.680903e-06, 4.696083e-06, 4.575953e-06, 4.530512e-06, 
    4.511263e-06, 4.494435e-06, 4.453611e-06, 4.481788e-06, 4.470671e-06, 
    4.497134e-06, 4.513983e-06, 4.505646e-06, 4.5572e-06, 4.537128e-06, 
    4.643282e-06, 4.597434e-06, 4.717353e-06, 4.688542e-06, 4.724269e-06, 
    4.706023e-06, 4.737304e-06, 4.709148e-06, 4.757963e-06, 4.76862e-06, 
    4.761337e-06, 4.789338e-06, 4.70759e-06, 4.738918e-06, 4.505413e-06, 
    4.506772e-06, 4.513106e-06, 4.485291e-06, 4.483592e-06, 4.458166e-06, 
    4.480786e-06, 4.490434e-06, 4.51496e-06, 4.529495e-06, 4.54333e-06, 
    4.573809e-06, 4.607949e-06, 4.655862e-06, 4.690407e-06, 4.713622e-06, 
    4.699381e-06, 4.711953e-06, 4.6979e-06, 4.691319e-06, 4.764627e-06, 
    4.723407e-06, 4.785306e-06, 4.781872e-06, 4.753827e-06, 4.782259e-06, 
    4.507727e-06, 4.499906e-06, 4.472801e-06, 4.494007e-06, 4.4554e-06, 
    4.476995e-06, 4.489432e-06, 4.53755e-06, 4.548147e-06, 4.557987e-06, 
    4.577444e-06, 4.602464e-06, 4.646493e-06, 4.68494e-06, 4.720149e-06, 
    4.717565e-06, 4.718475e-06, 4.726355e-06, 4.706847e-06, 4.729561e-06, 
    4.733378e-06, 4.723401e-06, 4.781412e-06, 4.76481e-06, 4.781799e-06, 
    4.770986e-06, 4.502448e-06, 4.515613e-06, 4.508497e-06, 4.521882e-06, 
    4.512451e-06, 4.554451e-06, 4.567074e-06, 4.626332e-06, 4.601972e-06, 
    4.640763e-06, 4.605905e-06, 4.612074e-06, 4.642035e-06, 4.607786e-06, 
    4.682819e-06, 4.631897e-06, 4.726661e-06, 4.67562e-06, 4.729868e-06, 
    4.719996e-06, 4.736343e-06, 4.751004e-06, 4.769473e-06, 4.80363e-06, 
    4.795711e-06, 4.824332e-06, 4.535267e-06, 4.552398e-06, 4.550887e-06, 
    4.568839e-06, 4.582135e-06, 4.611006e-06, 4.657469e-06, 4.639974e-06, 
    4.67211e-06, 4.678574e-06, 4.629757e-06, 4.659707e-06, 4.563877e-06, 
    4.579305e-06, 4.570115e-06, 4.536618e-06, 4.644005e-06, 4.588766e-06, 
    4.690979e-06, 4.660896e-06, 4.748913e-06, 4.705058e-06, 4.791355e-06, 
    4.828445e-06, 4.863449e-06, 4.904494e-06, 4.561757e-06, 4.550104e-06, 
    4.570976e-06, 4.599921e-06, 4.626839e-06, 4.662729e-06, 4.666406e-06, 
    4.673146e-06, 4.690618e-06, 4.705329e-06, 4.675279e-06, 4.70902e-06, 
    4.58289e-06, 4.648812e-06, 4.545703e-06, 4.576654e-06, 4.598211e-06, 
    4.588748e-06, 4.637976e-06, 4.64961e-06, 4.697011e-06, 4.672482e-06, 
    4.819282e-06, 4.754106e-06, 4.935832e-06, 4.884773e-06, 4.546036e-06, 
    4.561716e-06, 4.616462e-06, 4.59038e-06, 4.665128e-06, 4.683604e-06, 
    4.698644e-06, 4.717901e-06, 4.719981e-06, 4.731407e-06, 4.712689e-06, 
    4.730667e-06, 4.662806e-06, 4.693082e-06, 4.610189e-06, 4.63031e-06, 
    4.621048e-06, 4.6109e-06, 4.642251e-06, 4.675752e-06, 4.676466e-06, 
    4.68723e-06, 4.717621e-06, 4.665432e-06, 4.827726e-06, 4.727235e-06, 
    4.578839e-06, 4.609154e-06, 4.613487e-06, 4.60173e-06, 4.68175e-06, 
    4.652691e-06, 4.731128e-06, 4.709876e-06, 4.744717e-06, 4.727391e-06, 
    4.724845e-06, 4.702634e-06, 4.688828e-06, 4.654023e-06, 4.625781e-06, 
    4.603434e-06, 4.608626e-06, 4.633187e-06, 4.677803e-06, 4.72017e-06, 
    4.710877e-06, 4.742065e-06, 4.659692e-06, 4.694162e-06, 4.680828e-06, 
    4.715629e-06, 4.63951e-06, 4.704306e-06, 4.623007e-06, 4.630112e-06, 
    4.652115e-06, 4.696506e-06, 4.706346e-06, 4.716867e-06, 4.710373e-06, 
    4.678938e-06, 4.673795e-06, 4.651579e-06, 4.645454e-06, 4.628564e-06, 
    4.614601e-06, 4.627359e-06, 4.640773e-06, 4.67895e-06, 4.713465e-06, 
    4.751214e-06, 4.760469e-06, 4.804771e-06, 4.768699e-06, 4.828288e-06, 
    4.777613e-06, 4.865467e-06, 4.708068e-06, 4.77612e-06, 4.653116e-06, 
    4.666304e-06, 4.690199e-06, 4.745185e-06, 4.715464e-06, 4.750229e-06, 
    4.673593e-06, 4.634036e-06, 4.623821e-06, 4.604792e-06, 4.624257e-06, 
    4.622672e-06, 4.641327e-06, 4.635328e-06, 4.68022e-06, 4.656084e-06, 
    4.724781e-06, 4.749953e-06, 4.82133e-06, 4.8653e-06, 4.910219e-06, 
    4.930103e-06, 4.936162e-06, 4.938695e-06,
  4.331477e-06, 4.372477e-06, 4.364491e-06, 4.397667e-06, 4.379247e-06, 
    4.400993e-06, 4.339774e-06, 4.37411e-06, 4.352175e-06, 4.335159e-06, 
    4.46239e-06, 4.399149e-06, 4.528519e-06, 4.487857e-06, 4.590327e-06, 
    4.522182e-06, 4.604125e-06, 4.58835e-06, 4.635895e-06, 4.62225e-06, 
    4.683322e-06, 4.642198e-06, 4.715122e-06, 4.673483e-06, 4.679987e-06, 
    4.640845e-06, 4.411838e-06, 4.454495e-06, 4.409318e-06, 4.415387e-06, 
    4.412662e-06, 4.379629e-06, 4.363028e-06, 4.328349e-06, 4.334635e-06, 
    4.360109e-06, 4.418117e-06, 4.398383e-06, 4.448191e-06, 4.447063e-06, 
    4.502821e-06, 4.47764e-06, 4.571844e-06, 4.544975e-06, 4.62282e-06, 
    4.603184e-06, 4.621897e-06, 4.616219e-06, 4.621971e-06, 4.593189e-06, 
    4.605511e-06, 4.580222e-06, 4.482352e-06, 4.511013e-06, 4.425789e-06, 
    4.374919e-06, 4.341277e-06, 4.317481e-06, 4.320842e-06, 4.327252e-06, 
    4.360259e-06, 4.391397e-06, 4.415198e-06, 4.431154e-06, 4.446901e-06, 
    4.494736e-06, 4.520145e-06, 4.577288e-06, 4.566947e-06, 4.584469e-06, 
    4.601233e-06, 4.629447e-06, 4.624797e-06, 4.637248e-06, 4.584004e-06, 
    4.619359e-06, 4.561063e-06, 4.576973e-06, 4.451198e-06, 4.403702e-06, 
    4.383597e-06, 4.366026e-06, 4.323426e-06, 4.352824e-06, 4.341225e-06, 
    4.368843e-06, 4.386437e-06, 4.377731e-06, 4.431591e-06, 4.410615e-06, 
    4.521653e-06, 4.473665e-06, 4.599276e-06, 4.569069e-06, 4.60653e-06, 
    4.587396e-06, 4.620205e-06, 4.590672e-06, 4.641885e-06, 4.653074e-06, 
    4.645427e-06, 4.67483e-06, 4.589038e-06, 4.621898e-06, 4.377488e-06, 
    4.378907e-06, 4.385521e-06, 4.356481e-06, 4.354707e-06, 4.328178e-06, 
    4.351779e-06, 4.361849e-06, 4.387457e-06, 4.40264e-06, 4.417095e-06, 
    4.448955e-06, 4.484667e-06, 4.534827e-06, 4.571024e-06, 4.595364e-06, 
    4.580431e-06, 4.593614e-06, 4.578879e-06, 4.571979e-06, 4.648881e-06, 
    4.605626e-06, 4.670595e-06, 4.666988e-06, 4.637545e-06, 4.667395e-06, 
    4.379904e-06, 4.371738e-06, 4.343447e-06, 4.36558e-06, 4.325293e-06, 
    4.347823e-06, 4.360804e-06, 4.411055e-06, 4.42213e-06, 4.432414e-06, 
    4.452756e-06, 4.478928e-06, 4.525015e-06, 4.565294e-06, 4.602209e-06, 
    4.599499e-06, 4.600453e-06, 4.608718e-06, 4.588259e-06, 4.612081e-06, 
    4.616086e-06, 4.60562e-06, 4.666505e-06, 4.649072e-06, 4.666912e-06, 
    4.655556e-06, 4.374391e-06, 4.388139e-06, 4.380708e-06, 4.394687e-06, 
    4.384837e-06, 4.428718e-06, 4.441914e-06, 4.503906e-06, 4.478412e-06, 
    4.519015e-06, 4.482528e-06, 4.488984e-06, 4.520347e-06, 4.484496e-06, 
    4.563071e-06, 4.509733e-06, 4.60904e-06, 4.555528e-06, 4.612403e-06, 
    4.602049e-06, 4.619197e-06, 4.634582e-06, 4.653969e-06, 4.689844e-06, 
    4.681524e-06, 4.711599e-06, 4.40867e-06, 4.426572e-06, 4.424992e-06, 
    4.443759e-06, 4.457663e-06, 4.487865e-06, 4.53651e-06, 4.518188e-06, 
    4.551849e-06, 4.558622e-06, 4.507491e-06, 4.538855e-06, 4.438571e-06, 
    4.454704e-06, 4.445093e-06, 4.410082e-06, 4.52241e-06, 4.464598e-06, 
    4.571624e-06, 4.5401e-06, 4.632387e-06, 4.586384e-06, 4.676948e-06, 
    4.715924e-06, 4.752733e-06, 4.795932e-06, 4.436355e-06, 4.424174e-06, 
    4.445993e-06, 4.476267e-06, 4.504437e-06, 4.542021e-06, 4.545873e-06, 
    4.552934e-06, 4.571245e-06, 4.586668e-06, 4.55517e-06, 4.590538e-06, 
    4.458453e-06, 4.527444e-06, 4.419575e-06, 4.451931e-06, 4.474479e-06, 
    4.464579e-06, 4.516095e-06, 4.528279e-06, 4.577947e-06, 4.552238e-06, 
    4.706292e-06, 4.637838e-06, 4.828938e-06, 4.775171e-06, 4.419923e-06, 
    4.436311e-06, 4.493576e-06, 4.466286e-06, 4.544534e-06, 4.563894e-06, 
    4.579658e-06, 4.599851e-06, 4.602032e-06, 4.614019e-06, 4.594385e-06, 
    4.613241e-06, 4.542101e-06, 4.573827e-06, 4.48701e-06, 4.50807e-06, 
    4.498375e-06, 4.487754e-06, 4.520573e-06, 4.555665e-06, 4.556413e-06, 
    4.567694e-06, 4.59956e-06, 4.544852e-06, 4.715168e-06, 4.609644e-06, 
    4.454215e-06, 4.485928e-06, 4.490462e-06, 4.47816e-06, 4.561951e-06, 
    4.531506e-06, 4.613726e-06, 4.591435e-06, 4.627983e-06, 4.609805e-06, 
    4.607134e-06, 4.583841e-06, 4.569369e-06, 4.532901e-06, 4.503329e-06, 
    4.479943e-06, 4.485375e-06, 4.511082e-06, 4.557815e-06, 4.602231e-06, 
    4.592485e-06, 4.625201e-06, 4.538839e-06, 4.574961e-06, 4.560985e-06, 
    4.597468e-06, 4.517702e-06, 4.585597e-06, 4.500426e-06, 4.507862e-06, 
    4.530903e-06, 4.577418e-06, 4.587734e-06, 4.598767e-06, 4.591957e-06, 
    4.559004e-06, 4.553614e-06, 4.530341e-06, 4.523927e-06, 4.506242e-06, 
    4.491628e-06, 4.504981e-06, 4.519025e-06, 4.559016e-06, 4.5952e-06, 
    4.634802e-06, 4.644516e-06, 4.691044e-06, 4.653156e-06, 4.71576e-06, 
    4.662518e-06, 4.754858e-06, 4.58954e-06, 4.660949e-06, 4.531951e-06, 
    4.545766e-06, 4.570807e-06, 4.628476e-06, 4.597296e-06, 4.633769e-06, 
    4.553403e-06, 4.511972e-06, 4.501278e-06, 4.481363e-06, 4.501733e-06, 
    4.500075e-06, 4.519604e-06, 4.513324e-06, 4.560347e-06, 4.535059e-06, 
    4.607068e-06, 4.633479e-06, 4.708444e-06, 4.754681e-06, 4.801959e-06, 
    4.822903e-06, 4.829285e-06, 4.831955e-06,
  4.364439e-06, 4.40508e-06, 4.397161e-06, 4.430066e-06, 4.411794e-06, 
    4.433366e-06, 4.372659e-06, 4.4067e-06, 4.38495e-06, 4.368086e-06, 
    4.494324e-06, 4.431537e-06, 4.56006e-06, 4.519628e-06, 4.621583e-06, 
    4.553758e-06, 4.635328e-06, 4.619614e-06, 4.666991e-06, 4.653389e-06, 
    4.714299e-06, 4.673276e-06, 4.746046e-06, 4.704481e-06, 4.710971e-06, 
    4.671926e-06, 4.444128e-06, 4.486481e-06, 4.441627e-06, 4.44765e-06, 
    4.444946e-06, 4.412173e-06, 4.395712e-06, 4.361338e-06, 4.367566e-06, 
    4.392817e-06, 4.45036e-06, 4.430776e-06, 4.480218e-06, 4.479098e-06, 
    4.534503e-06, 4.509474e-06, 4.603176e-06, 4.576431e-06, 4.653956e-06, 
    4.63439e-06, 4.653037e-06, 4.647378e-06, 4.653111e-06, 4.624434e-06, 
    4.636708e-06, 4.611518e-06, 4.514156e-06, 4.542649e-06, 4.457975e-06, 
    4.407503e-06, 4.37415e-06, 4.350572e-06, 4.3539e-06, 4.360251e-06, 
    4.392965e-06, 4.423845e-06, 4.447462e-06, 4.4633e-06, 4.478937e-06, 
    4.526468e-06, 4.551731e-06, 4.608597e-06, 4.598301e-06, 4.615748e-06, 
    4.632446e-06, 4.660563e-06, 4.655928e-06, 4.66834e-06, 4.615285e-06, 
    4.650508e-06, 4.592443e-06, 4.608284e-06, 4.483208e-06, 4.436054e-06, 
    4.41611e-06, 4.398683e-06, 4.356461e-06, 4.385595e-06, 4.374097e-06, 
    4.401476e-06, 4.418926e-06, 4.41029e-06, 4.463734e-06, 4.442913e-06, 
    4.553231e-06, 4.505524e-06, 4.630497e-06, 4.600413e-06, 4.637724e-06, 
    4.618662e-06, 4.651351e-06, 4.621926e-06, 4.672963e-06, 4.684121e-06, 
    4.676495e-06, 4.705824e-06, 4.620298e-06, 4.653039e-06, 4.410048e-06, 
    4.411456e-06, 4.418017e-06, 4.389221e-06, 4.387462e-06, 4.361168e-06, 
    4.384558e-06, 4.394542e-06, 4.419937e-06, 4.435e-06, 4.449344e-06, 
    4.480977e-06, 4.516458e-06, 4.566336e-06, 4.60236e-06, 4.626599e-06, 
    4.611727e-06, 4.624856e-06, 4.610181e-06, 4.603311e-06, 4.67994e-06, 
    4.636824e-06, 4.701599e-06, 4.698001e-06, 4.668636e-06, 4.698406e-06, 
    4.412445e-06, 4.404346e-06, 4.376299e-06, 4.39824e-06, 4.35831e-06, 
    4.380638e-06, 4.393506e-06, 4.443351e-06, 4.454342e-06, 4.464552e-06, 
    4.484752e-06, 4.510753e-06, 4.556574e-06, 4.596656e-06, 4.633418e-06, 
    4.630719e-06, 4.631669e-06, 4.639904e-06, 4.619522e-06, 4.643255e-06, 
    4.647246e-06, 4.636817e-06, 4.697519e-06, 4.68013e-06, 4.697924e-06, 
    4.686597e-06, 4.406977e-06, 4.420613e-06, 4.413242e-06, 4.427109e-06, 
    4.417338e-06, 4.460883e-06, 4.473985e-06, 4.535583e-06, 4.510242e-06, 
    4.550607e-06, 4.514331e-06, 4.520748e-06, 4.551933e-06, 4.516286e-06, 
    4.594443e-06, 4.541377e-06, 4.640224e-06, 4.586936e-06, 4.643576e-06, 
    4.633258e-06, 4.650346e-06, 4.665682e-06, 4.685014e-06, 4.720809e-06, 
    4.712505e-06, 4.742528e-06, 4.440984e-06, 4.458752e-06, 4.457184e-06, 
    4.475817e-06, 4.489626e-06, 4.519636e-06, 4.568009e-06, 4.549784e-06, 
    4.583273e-06, 4.590013e-06, 4.539146e-06, 4.570342e-06, 4.470665e-06, 
    4.486687e-06, 4.477141e-06, 4.442385e-06, 4.553984e-06, 4.496516e-06, 
    4.602957e-06, 4.571581e-06, 4.663494e-06, 4.617656e-06, 4.707938e-06, 
    4.746848e-06, 4.783622e-06, 4.826822e-06, 4.468464e-06, 4.456371e-06, 
    4.478034e-06, 4.50811e-06, 4.53611e-06, 4.573492e-06, 4.577325e-06, 
    4.584353e-06, 4.602579e-06, 4.617938e-06, 4.586578e-06, 4.621792e-06, 
    4.490413e-06, 4.55899e-06, 4.451807e-06, 4.483933e-06, 4.506333e-06, 
    4.496496e-06, 4.547702e-06, 4.55982e-06, 4.609254e-06, 4.58366e-06, 
    4.73723e-06, 4.668929e-06, 4.859856e-06, 4.806057e-06, 4.452151e-06, 
    4.468421e-06, 4.525313e-06, 4.498192e-06, 4.575993e-06, 4.595261e-06, 
    4.610957e-06, 4.63107e-06, 4.633242e-06, 4.645186e-06, 4.625624e-06, 
    4.644411e-06, 4.573572e-06, 4.605151e-06, 4.518786e-06, 4.539722e-06, 
    4.530083e-06, 4.519525e-06, 4.552156e-06, 4.587072e-06, 4.587815e-06, 
    4.599045e-06, 4.630783e-06, 4.576309e-06, 4.746096e-06, 4.640829e-06, 
    4.486201e-06, 4.517712e-06, 4.522217e-06, 4.50999e-06, 4.593328e-06, 
    4.563031e-06, 4.644894e-06, 4.622686e-06, 4.659104e-06, 4.640987e-06, 
    4.638325e-06, 4.615123e-06, 4.600713e-06, 4.564419e-06, 4.535008e-06, 
    4.511761e-06, 4.517161e-06, 4.542718e-06, 4.589211e-06, 4.633441e-06, 
    4.623732e-06, 4.65633e-06, 4.570326e-06, 4.60628e-06, 4.592366e-06, 
    4.628695e-06, 4.549301e-06, 4.616874e-06, 4.532121e-06, 4.539515e-06, 
    4.562431e-06, 4.608728e-06, 4.618999e-06, 4.62999e-06, 4.623205e-06, 
    4.590394e-06, 4.58503e-06, 4.561872e-06, 4.555493e-06, 4.537905e-06, 
    4.523376e-06, 4.536651e-06, 4.550616e-06, 4.590406e-06, 4.626436e-06, 
    4.665901e-06, 4.675586e-06, 4.722008e-06, 4.684205e-06, 4.746687e-06, 
    4.693545e-06, 4.78575e-06, 4.620801e-06, 4.691978e-06, 4.563474e-06, 
    4.577219e-06, 4.602144e-06, 4.659596e-06, 4.628524e-06, 4.664872e-06, 
    4.584819e-06, 4.543603e-06, 4.532968e-06, 4.513174e-06, 4.533421e-06, 
    4.531772e-06, 4.551192e-06, 4.544946e-06, 4.591731e-06, 4.566566e-06, 
    4.63826e-06, 4.664583e-06, 4.739378e-06, 4.785571e-06, 4.832852e-06, 
    4.853813e-06, 4.860203e-06, 4.862876e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SNOW_SOURCES =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SOIL1C =
  5.777962, 5.777942, 5.777946, 5.77793, 5.777939, 5.777928, 5.777958, 
    5.777941, 5.777952, 5.77796, 5.777898, 5.777929, 5.777866, 5.777886, 
    5.777836, 5.777869, 5.77783, 5.777837, 5.777814, 5.777821, 5.777792, 
    5.777812, 5.777777, 5.777797, 5.777793, 5.777812, 5.777923, 5.777902, 
    5.777924, 5.777921, 5.777923, 5.777938, 5.777947, 5.777964, 5.777961, 
    5.777948, 5.77792, 5.777929, 5.777905, 5.777905, 5.777878, 5.777891, 
    5.777845, 5.777858, 5.777821, 5.77783, 5.777821, 5.777824, 5.777821, 
    5.777835, 5.777829, 5.777841, 5.777888, 5.777874, 5.777916, 5.777941, 
    5.777957, 5.777969, 5.777967, 5.777965, 5.777948, 5.777933, 5.777921, 
    5.777914, 5.777905, 5.777883, 5.77787, 5.777843, 5.777848, 5.777839, 
    5.777831, 5.777818, 5.77782, 5.777814, 5.777839, 5.777822, 5.77785, 
    5.777843, 5.777904, 5.777927, 5.777936, 5.777945, 5.777966, 5.777952, 
    5.777957, 5.777944, 5.777935, 5.777939, 5.777913, 5.777924, 5.777869, 
    5.777893, 5.777832, 5.777846, 5.777829, 5.777838, 5.777822, 5.777836, 
    5.777812, 5.777806, 5.77781, 5.777796, 5.777837, 5.777821, 5.77794, 
    5.777939, 5.777936, 5.77795, 5.777951, 5.777964, 5.777952, 5.777947, 
    5.777935, 5.777927, 5.77792, 5.777905, 5.777887, 5.777863, 5.777845, 
    5.777834, 5.777841, 5.777835, 5.777842, 5.777845, 5.777808, 5.777829, 
    5.777798, 5.7778, 5.777814, 5.7778, 5.777938, 5.777943, 5.777956, 
    5.777946, 5.777966, 5.777954, 5.777948, 5.777923, 5.777918, 5.777913, 
    5.777903, 5.77789, 5.777868, 5.777848, 5.777831, 5.777832, 5.777832, 
    5.777828, 5.777837, 5.777826, 5.777824, 5.777829, 5.7778, 5.777808, 
    5.7778, 5.777805, 5.777941, 5.777935, 5.777938, 5.777931, 5.777936, 
    5.777915, 5.777908, 5.777878, 5.77789, 5.777871, 5.777888, 5.777885, 
    5.77787, 5.777887, 5.777849, 5.777875, 5.777827, 5.777853, 5.777826, 
    5.777831, 5.777822, 5.777815, 5.777806, 5.777789, 5.777793, 5.777779, 
    5.777925, 5.777915, 5.777916, 5.777907, 5.7779, 5.777886, 5.777862, 
    5.777871, 5.777855, 5.777852, 5.777876, 5.777861, 5.77791, 5.777902, 
    5.777906, 5.777924, 5.777869, 5.777897, 5.777845, 5.777861, 5.777816, 
    5.777838, 5.777795, 5.777776, 5.777759, 5.777739, 5.777911, 5.777917, 
    5.777906, 5.777891, 5.777878, 5.77786, 5.777858, 5.777854, 5.777845, 
    5.777838, 5.777853, 5.777836, 5.7779, 5.777866, 5.777919, 5.777903, 
    5.777892, 5.777897, 5.777872, 5.777866, 5.777842, 5.777854, 5.777781, 
    5.777813, 5.777723, 5.777749, 5.777919, 5.777911, 5.777883, 5.777896, 
    5.777858, 5.777849, 5.777842, 5.777832, 5.777831, 5.777825, 5.777834, 
    5.777825, 5.77786, 5.777844, 5.777886, 5.777876, 5.777881, 5.777886, 
    5.77787, 5.777853, 5.777853, 5.777847, 5.777832, 5.777858, 5.777777, 
    5.777827, 5.777902, 5.777887, 5.777884, 5.777891, 5.77785, 5.777864, 
    5.777825, 5.777836, 5.777818, 5.777827, 5.777828, 5.77784, 5.777846, 
    5.777864, 5.777878, 5.77789, 5.777887, 5.777874, 5.777852, 5.777831, 
    5.777835, 5.77782, 5.777861, 5.777843, 5.777851, 5.777833, 5.777871, 
    5.777839, 5.77788, 5.777876, 5.777865, 5.777843, 5.777838, 5.777833, 
    5.777835, 5.777852, 5.777854, 5.777865, 5.777868, 5.777877, 5.777884, 
    5.777877, 5.777871, 5.777852, 5.777834, 5.777815, 5.777811, 5.777788, 
    5.777806, 5.777777, 5.777802, 5.777758, 5.777837, 5.777802, 5.777864, 
    5.777858, 5.777846, 5.777818, 5.777833, 5.777815, 5.777854, 5.777874, 
    5.777879, 5.777889, 5.777879, 5.77788, 5.77787, 5.777874, 5.777851, 
    5.777863, 5.777828, 5.777816, 5.77778, 5.777758, 5.777736, 5.777726, 
    5.777723, 5.777722 ;

 SOIL1C_TO_SOIL2C =
  3.180418e-08, 3.194395e-08, 3.191678e-08, 3.202952e-08, 3.196698e-08, 
    3.20408e-08, 3.183252e-08, 3.19495e-08, 3.187482e-08, 3.181676e-08, 
    3.224829e-08, 3.203455e-08, 3.24703e-08, 3.233398e-08, 3.267639e-08, 
    3.244909e-08, 3.272223e-08, 3.266983e-08, 3.282751e-08, 3.278234e-08, 
    3.298403e-08, 3.284836e-08, 3.308857e-08, 3.295163e-08, 3.297305e-08, 
    3.284389e-08, 3.207756e-08, 3.222168e-08, 3.206902e-08, 3.208957e-08, 
    3.208035e-08, 3.196827e-08, 3.191179e-08, 3.179349e-08, 3.181497e-08, 
    3.190186e-08, 3.209881e-08, 3.203195e-08, 3.220045e-08, 3.219664e-08, 
    3.238422e-08, 3.229965e-08, 3.261491e-08, 3.252531e-08, 3.278423e-08, 
    3.271911e-08, 3.278117e-08, 3.276235e-08, 3.278141e-08, 3.268592e-08, 
    3.272683e-08, 3.26428e-08, 3.231548e-08, 3.241168e-08, 3.212477e-08, 
    3.195225e-08, 3.183765e-08, 3.175633e-08, 3.176782e-08, 3.178974e-08, 
    3.190236e-08, 3.200825e-08, 3.208894e-08, 3.214291e-08, 3.219609e-08, 
    3.235708e-08, 3.244227e-08, 3.263303e-08, 3.25986e-08, 3.265692e-08, 
    3.271263e-08, 3.280617e-08, 3.279078e-08, 3.283199e-08, 3.265538e-08, 
    3.277276e-08, 3.257899e-08, 3.263199e-08, 3.221056e-08, 3.204999e-08, 
    3.198175e-08, 3.1922e-08, 3.177666e-08, 3.187703e-08, 3.183747e-08, 
    3.19316e-08, 3.199141e-08, 3.196183e-08, 3.214439e-08, 3.207341e-08, 
    3.244732e-08, 3.228627e-08, 3.270614e-08, 3.260567e-08, 3.273022e-08, 
    3.266666e-08, 3.277556e-08, 3.267755e-08, 3.284732e-08, 3.288429e-08, 
    3.285903e-08, 3.295607e-08, 3.267212e-08, 3.278117e-08, 3.196099e-08, 
    3.196582e-08, 3.19883e-08, 3.18895e-08, 3.188345e-08, 3.179291e-08, 
    3.187347e-08, 3.190778e-08, 3.199487e-08, 3.204639e-08, 3.209535e-08, 
    3.220302e-08, 3.232326e-08, 3.24914e-08, 3.261218e-08, 3.269314e-08, 
    3.26435e-08, 3.268733e-08, 3.263833e-08, 3.261536e-08, 3.287044e-08, 
    3.272721e-08, 3.294211e-08, 3.293022e-08, 3.283297e-08, 3.293156e-08, 
    3.196921e-08, 3.194144e-08, 3.184505e-08, 3.192049e-08, 3.178305e-08, 
    3.185998e-08, 3.190422e-08, 3.20749e-08, 3.21124e-08, 3.214717e-08, 
    3.221584e-08, 3.230397e-08, 3.245858e-08, 3.259309e-08, 3.271587e-08, 
    3.270688e-08, 3.271004e-08, 3.273748e-08, 3.266953e-08, 3.274863e-08, 
    3.276191e-08, 3.27272e-08, 3.292863e-08, 3.287108e-08, 3.292997e-08, 
    3.28925e-08, 3.195047e-08, 3.199719e-08, 3.197194e-08, 3.201941e-08, 
    3.198597e-08, 3.213467e-08, 3.217925e-08, 3.238785e-08, 3.230224e-08, 
    3.243849e-08, 3.231608e-08, 3.233777e-08, 3.244294e-08, 3.232269e-08, 
    3.258567e-08, 3.240739e-08, 3.273854e-08, 3.256052e-08, 3.27497e-08, 
    3.271535e-08, 3.277222e-08, 3.282317e-08, 3.288725e-08, 3.300551e-08, 
    3.297812e-08, 3.307701e-08, 3.206683e-08, 3.212742e-08, 3.212208e-08, 
    3.218549e-08, 3.223238e-08, 3.233402e-08, 3.249702e-08, 3.243573e-08, 
    3.254826e-08, 3.257085e-08, 3.239989e-08, 3.250486e-08, 3.216797e-08, 
    3.22224e-08, 3.218999e-08, 3.207161e-08, 3.244985e-08, 3.225574e-08, 
    3.261418e-08, 3.250902e-08, 3.28159e-08, 3.266329e-08, 3.296305e-08, 
    3.30912e-08, 3.321179e-08, 3.335272e-08, 3.216049e-08, 3.211931e-08, 
    3.219303e-08, 3.229502e-08, 3.238964e-08, 3.251544e-08, 3.252831e-08, 
    3.255187e-08, 3.261292e-08, 3.266424e-08, 3.255933e-08, 3.267711e-08, 
    3.223503e-08, 3.24667e-08, 3.210375e-08, 3.221305e-08, 3.228901e-08, 
    3.225568e-08, 3.242872e-08, 3.24695e-08, 3.263522e-08, 3.254956e-08, 
    3.305957e-08, 3.283393e-08, 3.346003e-08, 3.328507e-08, 3.210493e-08, 
    3.216034e-08, 3.235319e-08, 3.226143e-08, 3.252384e-08, 3.258842e-08, 
    3.264093e-08, 3.270804e-08, 3.271529e-08, 3.275505e-08, 3.268989e-08, 
    3.275248e-08, 3.251571e-08, 3.262151e-08, 3.233114e-08, 3.240182e-08, 
    3.236931e-08, 3.233365e-08, 3.244371e-08, 3.256098e-08, 3.256348e-08, 
    3.260108e-08, 3.270705e-08, 3.25249e-08, 3.30887e-08, 3.274052e-08, 
    3.222076e-08, 3.23275e-08, 3.234274e-08, 3.230139e-08, 3.258195e-08, 
    3.248029e-08, 3.275408e-08, 3.268009e-08, 3.280133e-08, 3.274108e-08, 
    3.273222e-08, 3.265484e-08, 3.260667e-08, 3.248496e-08, 3.238592e-08, 
    3.230739e-08, 3.232565e-08, 3.241192e-08, 3.256815e-08, 3.271595e-08, 
    3.268357e-08, 3.279212e-08, 3.250481e-08, 3.262528e-08, 3.257872e-08, 
    3.270013e-08, 3.24341e-08, 3.266065e-08, 3.237619e-08, 3.240113e-08, 
    3.247828e-08, 3.263346e-08, 3.266778e-08, 3.270445e-08, 3.268182e-08, 
    3.257212e-08, 3.255414e-08, 3.24764e-08, 3.245494e-08, 3.23957e-08, 
    3.234666e-08, 3.239147e-08, 3.243852e-08, 3.257216e-08, 3.269259e-08, 
    3.282389e-08, 3.285602e-08, 3.300944e-08, 3.288456e-08, 3.309064e-08, 
    3.291544e-08, 3.321871e-08, 3.267377e-08, 3.291028e-08, 3.248179e-08, 
    3.252795e-08, 3.261145e-08, 3.280295e-08, 3.269956e-08, 3.282047e-08, 
    3.255344e-08, 3.24149e-08, 3.237905e-08, 3.231217e-08, 3.238057e-08, 
    3.237501e-08, 3.244047e-08, 3.241944e-08, 3.25766e-08, 3.249218e-08, 
    3.2732e-08, 3.281951e-08, 3.306665e-08, 3.321815e-08, 3.337236e-08, 
    3.344044e-08, 3.346116e-08, 3.346982e-08 ;

 SOIL1C_TO_SOIL3C =
  3.772076e-10, 3.788659e-10, 3.785436e-10, 3.798811e-10, 3.791391e-10, 
    3.80015e-10, 3.775438e-10, 3.789318e-10, 3.780457e-10, 3.773569e-10, 
    3.824769e-10, 3.799408e-10, 3.851109e-10, 3.834936e-10, 3.875563e-10, 
    3.848593e-10, 3.881002e-10, 3.874785e-10, 3.893494e-10, 3.888135e-10, 
    3.912066e-10, 3.895968e-10, 3.92447e-10, 3.908221e-10, 3.910763e-10, 
    3.895437e-10, 3.804511e-10, 3.821611e-10, 3.803498e-10, 3.805937e-10, 
    3.804842e-10, 3.791545e-10, 3.784844e-10, 3.770808e-10, 3.773356e-10, 
    3.783665e-10, 3.807033e-10, 3.7991e-10, 3.819092e-10, 3.81864e-10, 
    3.840896e-10, 3.830862e-10, 3.868268e-10, 3.857637e-10, 3.888358e-10, 
    3.880632e-10, 3.887995e-10, 3.885763e-10, 3.888024e-10, 3.876693e-10, 
    3.881548e-10, 3.871577e-10, 3.832741e-10, 3.844155e-10, 3.810113e-10, 
    3.789644e-10, 3.776047e-10, 3.766399e-10, 3.767762e-10, 3.770363e-10, 
    3.783725e-10, 3.796288e-10, 3.805861e-10, 3.812266e-10, 3.818575e-10, 
    3.837676e-10, 3.847784e-10, 3.870418e-10, 3.866333e-10, 3.873253e-10, 
    3.879863e-10, 3.890962e-10, 3.889135e-10, 3.894025e-10, 3.87307e-10, 
    3.886997e-10, 3.864006e-10, 3.870295e-10, 3.820292e-10, 3.80124e-10, 
    3.793144e-10, 3.786055e-10, 3.768811e-10, 3.78072e-10, 3.776025e-10, 
    3.787193e-10, 3.79429e-10, 3.79078e-10, 3.812441e-10, 3.80402e-10, 
    3.848383e-10, 3.829275e-10, 3.879093e-10, 3.867171e-10, 3.88195e-10, 
    3.874409e-10, 3.88733e-10, 3.875701e-10, 3.895845e-10, 3.900232e-10, 
    3.897234e-10, 3.908748e-10, 3.875056e-10, 3.887995e-10, 3.790681e-10, 
    3.791254e-10, 3.793921e-10, 3.782198e-10, 3.781481e-10, 3.770738e-10, 
    3.780297e-10, 3.784368e-10, 3.794701e-10, 3.800813e-10, 3.806623e-10, 
    3.819397e-10, 3.833664e-10, 3.853613e-10, 3.867944e-10, 3.877551e-10, 
    3.87166e-10, 3.876861e-10, 3.871047e-10, 3.868322e-10, 3.898588e-10, 
    3.881593e-10, 3.907092e-10, 3.905681e-10, 3.894142e-10, 3.90584e-10, 
    3.791656e-10, 3.788362e-10, 3.776925e-10, 3.785876e-10, 3.769569e-10, 
    3.778697e-10, 3.783945e-10, 3.804196e-10, 3.808645e-10, 3.81277e-10, 
    3.820918e-10, 3.831375e-10, 3.849719e-10, 3.865679e-10, 3.880248e-10, 
    3.879181e-10, 3.879556e-10, 3.882811e-10, 3.874749e-10, 3.884135e-10, 
    3.88571e-10, 3.881591e-10, 3.905492e-10, 3.898664e-10, 3.905651e-10, 
    3.901205e-10, 3.789432e-10, 3.794975e-10, 3.79198e-10, 3.797612e-10, 
    3.793645e-10, 3.811287e-10, 3.816577e-10, 3.841328e-10, 3.83117e-10, 
    3.847336e-10, 3.832812e-10, 3.835385e-10, 3.847864e-10, 3.833596e-10, 
    3.864799e-10, 3.843645e-10, 3.882938e-10, 3.861814e-10, 3.884261e-10, 
    3.880185e-10, 3.886934e-10, 3.892979e-10, 3.900583e-10, 3.914614e-10, 
    3.911365e-10, 3.923099e-10, 3.803238e-10, 3.810427e-10, 3.809794e-10, 
    3.817317e-10, 3.822881e-10, 3.83494e-10, 3.854281e-10, 3.847008e-10, 
    3.86036e-10, 3.86304e-10, 3.842755e-10, 3.85521e-10, 3.815238e-10, 
    3.821697e-10, 3.817851e-10, 3.803805e-10, 3.848684e-10, 3.825653e-10, 
    3.868181e-10, 3.855705e-10, 3.892117e-10, 3.874009e-10, 3.909576e-10, 
    3.924782e-10, 3.939091e-10, 3.955815e-10, 3.81435e-10, 3.809466e-10, 
    3.818212e-10, 3.830313e-10, 3.84154e-10, 3.856466e-10, 3.857993e-10, 
    3.860789e-10, 3.868031e-10, 3.874121e-10, 3.861673e-10, 3.875648e-10, 
    3.823195e-10, 3.850683e-10, 3.807619e-10, 3.820587e-10, 3.829599e-10, 
    3.825646e-10, 3.846176e-10, 3.851015e-10, 3.870678e-10, 3.860514e-10, 
    3.921029e-10, 3.894256e-10, 3.968547e-10, 3.947786e-10, 3.807759e-10, 
    3.814333e-10, 3.837215e-10, 3.826328e-10, 3.857462e-10, 3.865125e-10, 
    3.871355e-10, 3.879319e-10, 3.880178e-10, 3.884897e-10, 3.877165e-10, 
    3.884591e-10, 3.856497e-10, 3.869052e-10, 3.834599e-10, 3.842985e-10, 
    3.839127e-10, 3.834895e-10, 3.847955e-10, 3.861869e-10, 3.862166e-10, 
    3.866628e-10, 3.879201e-10, 3.857588e-10, 3.924486e-10, 3.883173e-10, 
    3.821503e-10, 3.834166e-10, 3.835975e-10, 3.831069e-10, 3.864357e-10, 
    3.852296e-10, 3.884782e-10, 3.876002e-10, 3.890387e-10, 3.883239e-10, 
    3.882187e-10, 3.873006e-10, 3.86729e-10, 3.852849e-10, 3.841099e-10, 
    3.83178e-10, 3.833947e-10, 3.844183e-10, 3.86272e-10, 3.880256e-10, 
    3.876415e-10, 3.889294e-10, 3.855204e-10, 3.869499e-10, 3.863974e-10, 
    3.87838e-10, 3.846815e-10, 3.873696e-10, 3.839944e-10, 3.842903e-10, 
    3.852056e-10, 3.870469e-10, 3.874542e-10, 3.878892e-10, 3.876207e-10, 
    3.863191e-10, 3.861058e-10, 3.851834e-10, 3.849287e-10, 3.842258e-10, 
    3.836439e-10, 3.841756e-10, 3.84734e-10, 3.863196e-10, 3.877486e-10, 
    3.893065e-10, 3.896877e-10, 3.915081e-10, 3.900263e-10, 3.924716e-10, 
    3.903927e-10, 3.939913e-10, 3.875253e-10, 3.903315e-10, 3.852473e-10, 
    3.85795e-10, 3.867857e-10, 3.89058e-10, 3.878312e-10, 3.892659e-10, 
    3.860975e-10, 3.844536e-10, 3.840283e-10, 3.832347e-10, 3.840464e-10, 
    3.839804e-10, 3.847571e-10, 3.845075e-10, 3.863723e-10, 3.853706e-10, 
    3.882161e-10, 3.892545e-10, 3.921869e-10, 3.939846e-10, 3.958144e-10, 
    3.966222e-10, 3.968681e-10, 3.969709e-10 ;

 SOIL1C_vr =
  19.97934, 19.97928, 19.97929, 19.97925, 19.97927, 19.97925, 19.97933, 
    19.97928, 19.97931, 19.97933, 19.97917, 19.97925, 19.97908, 19.97913, 
    19.979, 19.97909, 19.97898, 19.979, 19.97894, 19.97896, 19.97888, 
    19.97894, 19.97884, 19.9789, 19.97889, 19.97894, 19.97923, 19.97918, 
    19.97923, 19.97923, 19.97923, 19.97927, 19.9793, 19.97934, 19.97933, 
    19.9793, 19.97922, 19.97925, 19.97918, 19.97919, 19.97911, 19.97915, 
    19.97902, 19.97906, 19.97896, 19.97898, 19.97896, 19.97897, 19.97896, 
    19.979, 19.97898, 19.97901, 19.97914, 19.9791, 19.97921, 19.97928, 
    19.97932, 19.97935, 19.97935, 19.97934, 19.9793, 19.97926, 19.97923, 
    19.97921, 19.97919, 19.97912, 19.97909, 19.97902, 19.97903, 19.97901, 
    19.97899, 19.97895, 19.97896, 19.97894, 19.97901, 19.97896, 19.97904, 
    19.97902, 19.97918, 19.97924, 19.97927, 19.97929, 19.97935, 19.97931, 
    19.97932, 19.97929, 19.97927, 19.97928, 19.97921, 19.97923, 19.97909, 
    19.97915, 19.97899, 19.97903, 19.97898, 19.979, 19.97896, 19.979, 
    19.97894, 19.97892, 19.97893, 19.97889, 19.979, 19.97896, 19.97928, 
    19.97927, 19.97927, 19.9793, 19.97931, 19.97934, 19.97931, 19.9793, 
    19.97926, 19.97924, 19.97923, 19.97918, 19.97914, 19.97907, 19.97902, 
    19.97899, 19.97901, 19.979, 19.97902, 19.97902, 19.97893, 19.97898, 
    19.9789, 19.9789, 19.97894, 19.9789, 19.97927, 19.97928, 19.97932, 
    19.97929, 19.97935, 19.97931, 19.9793, 19.97923, 19.97922, 19.9792, 
    19.97918, 19.97914, 19.97908, 19.97903, 19.97898, 19.97899, 19.97899, 
    19.97898, 19.979, 19.97897, 19.97897, 19.97898, 19.9789, 19.97893, 
    19.9789, 19.97892, 19.97928, 19.97926, 19.97927, 19.97925, 19.97927, 
    19.97921, 19.97919, 19.97911, 19.97915, 19.97909, 19.97914, 19.97913, 
    19.97909, 19.97914, 19.97904, 19.9791, 19.97898, 19.97905, 19.97897, 
    19.97899, 19.97896, 19.97894, 19.97892, 19.97887, 19.97889, 19.97885, 
    19.97923, 19.97921, 19.97921, 19.97919, 19.97917, 19.97913, 19.97907, 
    19.97909, 19.97905, 19.97904, 19.97911, 19.97907, 19.9792, 19.97918, 
    19.97919, 19.97923, 19.97909, 19.97916, 19.97902, 19.97906, 19.97895, 
    19.97901, 19.97889, 19.97884, 19.9788, 19.97874, 19.9792, 19.97922, 
    19.97919, 19.97915, 19.97911, 19.97906, 19.97906, 19.97905, 19.97902, 
    19.97901, 19.97905, 19.979, 19.97917, 19.97908, 19.97922, 19.97918, 
    19.97915, 19.97916, 19.9791, 19.97908, 19.97902, 19.97905, 19.97885, 
    19.97894, 19.9787, 19.97877, 19.97922, 19.9792, 19.97912, 19.97916, 
    19.97906, 19.97903, 19.97902, 19.97899, 19.97899, 19.97897, 19.979, 
    19.97897, 19.97906, 19.97902, 19.97913, 19.97911, 19.97912, 19.97913, 
    19.97909, 19.97905, 19.97904, 19.97903, 19.97899, 19.97906, 19.97884, 
    19.97898, 19.97918, 19.97914, 19.97913, 19.97915, 19.97904, 19.97908, 
    19.97897, 19.979, 19.97895, 19.97898, 19.97898, 19.97901, 19.97903, 
    19.97907, 19.97911, 19.97914, 19.97914, 19.9791, 19.97904, 19.97898, 
    19.979, 19.97896, 19.97907, 19.97902, 19.97904, 19.97899, 19.97909, 
    19.97901, 19.97912, 19.97911, 19.97908, 19.97902, 19.979, 19.97899, 
    19.979, 19.97904, 19.97905, 19.97908, 19.97909, 19.97911, 19.97913, 
    19.97911, 19.97909, 19.97904, 19.97899, 19.97894, 19.97893, 19.97887, 
    19.97892, 19.97884, 19.97891, 19.97879, 19.979, 19.97891, 19.97908, 
    19.97906, 19.97902, 19.97895, 19.97899, 19.97894, 19.97905, 19.9791, 
    19.97911, 19.97914, 19.97911, 19.97912, 19.97909, 19.9791, 19.97904, 
    19.97907, 19.97898, 19.97895, 19.97885, 19.97879, 19.97873, 19.97871, 
    19.9787, 19.9787,
  19.981, 19.98093, 19.98095, 19.98089, 19.98092, 19.98088, 19.98099, 
    19.98093, 19.98097, 19.981, 19.98078, 19.98089, 19.98067, 19.98074, 
    19.98056, 19.98068, 19.98054, 19.98057, 19.98049, 19.98051, 19.98041, 
    19.98048, 19.98036, 19.98042, 19.98041, 19.98048, 19.98087, 19.98079, 
    19.98087, 19.98086, 19.98087, 19.98092, 19.98095, 19.98101, 19.981, 
    19.98096, 19.98086, 19.98089, 19.9808, 19.98081, 19.98071, 19.98075, 
    19.98059, 19.98064, 19.98051, 19.98054, 19.98051, 19.98052, 19.98051, 
    19.98056, 19.98054, 19.98058, 19.98075, 19.9807, 19.98084, 19.98093, 
    19.98099, 19.98103, 19.98102, 19.98101, 19.98096, 19.9809, 19.98086, 
    19.98083, 19.98081, 19.98072, 19.98068, 19.98059, 19.9806, 19.98057, 
    19.98055, 19.9805, 19.9805, 19.98048, 19.98057, 19.98051, 19.98061, 
    19.98059, 19.9808, 19.98088, 19.98092, 19.98095, 19.98102, 19.98097, 
    19.98099, 19.98094, 19.98091, 19.98092, 19.98083, 19.98087, 19.98068, 
    19.98076, 19.98055, 19.9806, 19.98054, 19.98057, 19.98051, 19.98056, 
    19.98048, 19.98046, 19.98047, 19.98042, 19.98057, 19.98051, 19.98093, 
    19.98092, 19.98091, 19.98096, 19.98096, 19.98101, 19.98097, 19.98095, 
    19.98091, 19.98088, 19.98086, 19.9808, 19.98074, 19.98066, 19.9806, 
    19.98055, 19.98058, 19.98056, 19.98058, 19.98059, 19.98046, 19.98054, 
    19.98043, 19.98043, 19.98048, 19.98043, 19.98092, 19.98094, 19.98099, 
    19.98095, 19.98102, 19.98098, 19.98096, 19.98087, 19.98085, 19.98083, 
    19.9808, 19.98075, 19.98067, 19.98061, 19.98054, 19.98055, 19.98055, 
    19.98053, 19.98057, 19.98053, 19.98052, 19.98054, 19.98044, 19.98046, 
    19.98043, 19.98045, 19.98093, 19.98091, 19.98092, 19.9809, 19.98091, 
    19.98084, 19.98082, 19.98071, 19.98075, 19.98068, 19.98075, 19.98073, 
    19.98068, 19.98074, 19.98061, 19.9807, 19.98053, 19.98062, 19.98053, 
    19.98054, 19.98051, 19.98049, 19.98046, 19.9804, 19.98041, 19.98036, 
    19.98087, 19.98084, 19.98084, 19.98081, 19.98079, 19.98074, 19.98065, 
    19.98068, 19.98063, 19.98062, 19.9807, 19.98065, 19.98082, 19.98079, 
    19.98081, 19.98087, 19.98068, 19.98078, 19.98059, 19.98065, 19.98049, 
    19.98057, 19.98042, 19.98035, 19.98029, 19.98022, 19.98083, 19.98084, 
    19.98081, 19.98076, 19.98071, 19.98064, 19.98064, 19.98063, 19.98059, 
    19.98057, 19.98062, 19.98056, 19.98079, 19.98067, 19.98085, 19.9808, 
    19.98076, 19.98078, 19.98069, 19.98067, 19.98058, 19.98063, 19.98037, 
    19.98048, 19.98017, 19.98026, 19.98085, 19.98083, 19.98073, 19.98077, 
    19.98064, 19.98061, 19.98058, 19.98055, 19.98054, 19.98052, 19.98056, 
    19.98052, 19.98064, 19.98059, 19.98074, 19.9807, 19.98072, 19.98074, 
    19.98068, 19.98062, 19.98062, 19.9806, 19.98055, 19.98064, 19.98036, 
    19.98053, 19.98079, 19.98074, 19.98073, 19.98075, 19.98061, 19.98066, 
    19.98052, 19.98056, 19.9805, 19.98053, 19.98054, 19.98057, 19.9806, 
    19.98066, 19.98071, 19.98075, 19.98074, 19.9807, 19.98062, 19.98054, 
    19.98056, 19.9805, 19.98065, 19.98059, 19.98061, 19.98055, 19.98069, 
    19.98057, 19.98071, 19.9807, 19.98066, 19.98059, 19.98057, 19.98055, 
    19.98056, 19.98062, 19.98063, 19.98067, 19.98067, 19.98071, 19.98073, 
    19.98071, 19.98068, 19.98062, 19.98055, 19.98049, 19.98047, 19.98039, 
    19.98046, 19.98035, 19.98044, 19.98029, 19.98056, 19.98045, 19.98066, 
    19.98064, 19.9806, 19.9805, 19.98055, 19.98049, 19.98063, 19.9807, 
    19.98071, 19.98075, 19.98071, 19.98072, 19.98068, 19.98069, 19.98061, 
    19.98066, 19.98054, 19.98049, 19.98037, 19.98029, 19.98021, 19.98018, 
    19.98017, 19.98016,
  19.98273, 19.98265, 19.98267, 19.9826, 19.98264, 19.9826, 19.98271, 
    19.98265, 19.98269, 19.98272, 19.98249, 19.9826, 19.98237, 19.98244, 
    19.98226, 19.98238, 19.98223, 19.98226, 19.98217, 19.9822, 19.98209, 
    19.98216, 19.98203, 19.98211, 19.9821, 19.98217, 19.98258, 19.9825, 
    19.98258, 19.98257, 19.98258, 19.98264, 19.98267, 19.98273, 19.98272, 
    19.98268, 19.98257, 19.9826, 19.98251, 19.98252, 19.98241, 19.98246, 
    19.98229, 19.98234, 19.9822, 19.98223, 19.9822, 19.98221, 19.9822, 
    19.98225, 19.98223, 19.98228, 19.98245, 19.9824, 19.98255, 19.98265, 
    19.98271, 19.98275, 19.98275, 19.98274, 19.98268, 19.98262, 19.98257, 
    19.98254, 19.98252, 19.98243, 19.98238, 19.98228, 19.9823, 19.98227, 
    19.98224, 19.98219, 19.98219, 19.98217, 19.98227, 19.9822, 19.98231, 
    19.98228, 19.98251, 19.9826, 19.98263, 19.98266, 19.98274, 19.98269, 
    19.98271, 19.98266, 19.98263, 19.98264, 19.98254, 19.98258, 19.98238, 
    19.98247, 19.98224, 19.98229, 19.98223, 19.98226, 19.9822, 19.98226, 
    19.98216, 19.98214, 19.98216, 19.98211, 19.98226, 19.9822, 19.98264, 
    19.98264, 19.98263, 19.98268, 19.98269, 19.98273, 19.98269, 19.98267, 
    19.98262, 19.9826, 19.98257, 19.98251, 19.98245, 19.98236, 19.98229, 
    19.98225, 19.98227, 19.98225, 19.98228, 19.98229, 19.98215, 19.98223, 
    19.98211, 19.98212, 19.98217, 19.98212, 19.98264, 19.98265, 19.98271, 
    19.98266, 19.98274, 19.9827, 19.98267, 19.98258, 19.98256, 19.98254, 
    19.98251, 19.98246, 19.98237, 19.9823, 19.98223, 19.98224, 19.98224, 
    19.98222, 19.98226, 19.98222, 19.98221, 19.98223, 19.98212, 19.98215, 
    19.98212, 19.98214, 19.98265, 19.98262, 19.98264, 19.98261, 19.98263, 
    19.98255, 19.98252, 19.98241, 19.98246, 19.98238, 19.98245, 19.98244, 
    19.98238, 19.98245, 19.98231, 19.9824, 19.98222, 19.98232, 19.98222, 
    19.98223, 19.9822, 19.98218, 19.98214, 19.98208, 19.98209, 19.98204, 
    19.98259, 19.98255, 19.98256, 19.98252, 19.9825, 19.98244, 19.98235, 
    19.98239, 19.98232, 19.98231, 19.9824, 19.98235, 19.98253, 19.9825, 
    19.98252, 19.98258, 19.98238, 19.98248, 19.98229, 19.98235, 19.98218, 
    19.98226, 19.9821, 19.98203, 19.98197, 19.98189, 19.98253, 19.98256, 
    19.98252, 19.98246, 19.98241, 19.98234, 19.98234, 19.98232, 19.98229, 
    19.98226, 19.98232, 19.98226, 19.98249, 19.98237, 19.98256, 19.98251, 
    19.98247, 19.98248, 19.98239, 19.98237, 19.98228, 19.98232, 19.98205, 
    19.98217, 19.98183, 19.98193, 19.98256, 19.98253, 19.98243, 19.98248, 
    19.98234, 19.9823, 19.98228, 19.98224, 19.98223, 19.98221, 19.98225, 
    19.98221, 19.98234, 19.98229, 19.98244, 19.9824, 19.98242, 19.98244, 
    19.98238, 19.98232, 19.98232, 19.9823, 19.98224, 19.98234, 19.98203, 
    19.98222, 19.9825, 19.98244, 19.98244, 19.98246, 19.98231, 19.98236, 
    19.98221, 19.98225, 19.98219, 19.98222, 19.98223, 19.98227, 19.98229, 
    19.98236, 19.98241, 19.98246, 19.98244, 19.9824, 19.98232, 19.98223, 
    19.98225, 19.98219, 19.98235, 19.98228, 19.98231, 19.98224, 19.98239, 
    19.98226, 19.98242, 19.9824, 19.98236, 19.98228, 19.98226, 19.98224, 
    19.98225, 19.98231, 19.98232, 19.98236, 19.98238, 19.98241, 19.98243, 
    19.98241, 19.98238, 19.98231, 19.98225, 19.98218, 19.98216, 19.98208, 
    19.98214, 19.98203, 19.98213, 19.98196, 19.98226, 19.98213, 19.98236, 
    19.98234, 19.98229, 19.98219, 19.98224, 19.98218, 19.98232, 19.9824, 
    19.98242, 19.98245, 19.98242, 19.98242, 19.98238, 19.9824, 19.98231, 
    19.98236, 19.98223, 19.98218, 19.98205, 19.98196, 19.98188, 19.98184, 
    19.98183, 19.98183,
  19.9841, 19.98403, 19.98404, 19.98398, 19.98401, 19.98397, 19.98409, 
    19.98402, 19.98406, 19.98409, 19.98386, 19.98398, 19.98375, 19.98382, 
    19.98363, 19.98376, 19.98361, 19.98364, 19.98355, 19.98358, 19.98347, 
    19.98354, 19.98341, 19.98349, 19.98347, 19.98355, 19.98396, 19.98388, 
    19.98396, 19.98395, 19.98395, 19.98401, 19.98405, 19.98411, 19.9841, 
    19.98405, 19.98394, 19.98398, 19.98389, 19.98389, 19.98379, 19.98384, 
    19.98367, 19.98372, 19.98358, 19.98361, 19.98358, 19.98359, 19.98358, 
    19.98363, 19.98361, 19.98365, 19.98383, 19.98378, 19.98393, 19.98402, 
    19.98409, 19.98413, 19.98412, 19.98411, 19.98405, 19.98399, 19.98395, 
    19.98392, 19.98389, 19.9838, 19.98376, 19.98366, 19.98368, 19.98364, 
    19.98361, 19.98356, 19.98357, 19.98355, 19.98365, 19.98358, 19.98369, 
    19.98366, 19.98388, 19.98397, 19.98401, 19.98404, 19.98412, 19.98406, 
    19.98409, 19.98403, 19.984, 19.98402, 19.98392, 19.98396, 19.98376, 
    19.98384, 19.98362, 19.98367, 19.98361, 19.98364, 19.98358, 19.98363, 
    19.98354, 19.98352, 19.98354, 19.98348, 19.98364, 19.98358, 19.98402, 
    19.98402, 19.984, 19.98406, 19.98406, 19.98411, 19.98407, 19.98405, 
    19.984, 19.98397, 19.98395, 19.98389, 19.98382, 19.98373, 19.98367, 
    19.98363, 19.98365, 19.98363, 19.98365, 19.98367, 19.98353, 19.98361, 
    19.98349, 19.9835, 19.98355, 19.9835, 19.98401, 19.98403, 19.98408, 
    19.98404, 19.98411, 19.98407, 19.98405, 19.98396, 19.98394, 19.98392, 
    19.98388, 19.98383, 19.98375, 19.98368, 19.98361, 19.98362, 19.98362, 
    19.9836, 19.98364, 19.98359, 19.98359, 19.98361, 19.9835, 19.98353, 
    19.9835, 19.98352, 19.98402, 19.984, 19.98401, 19.98399, 19.984, 
    19.98392, 19.9839, 19.98379, 19.98384, 19.98376, 19.98383, 19.98382, 
    19.98376, 19.98382, 19.98368, 19.98378, 19.9836, 19.9837, 19.98359, 
    19.98361, 19.98358, 19.98355, 19.98352, 19.98346, 19.98347, 19.98342, 
    19.98396, 19.98393, 19.98393, 19.9839, 19.98387, 19.98382, 19.98373, 
    19.98376, 19.9837, 19.98369, 19.98378, 19.98373, 19.98391, 19.98388, 
    19.98389, 19.98396, 19.98376, 19.98386, 19.98367, 19.98372, 19.98356, 
    19.98364, 19.98348, 19.98341, 19.98335, 19.98327, 19.98391, 19.98393, 
    19.98389, 19.98384, 19.98379, 19.98372, 19.98371, 19.9837, 19.98367, 
    19.98364, 19.9837, 19.98363, 19.98387, 19.98375, 19.98394, 19.98388, 
    19.98384, 19.98386, 19.98377, 19.98375, 19.98366, 19.9837, 19.98343, 
    19.98355, 19.98322, 19.98331, 19.98394, 19.98391, 19.98381, 19.98386, 
    19.98372, 19.98368, 19.98365, 19.98362, 19.98361, 19.98359, 19.98363, 
    19.98359, 19.98372, 19.98366, 19.98382, 19.98378, 19.9838, 19.98382, 
    19.98376, 19.9837, 19.98369, 19.98368, 19.98362, 19.98372, 19.98341, 
    19.9836, 19.98388, 19.98382, 19.98381, 19.98384, 19.98368, 19.98374, 
    19.98359, 19.98363, 19.98357, 19.9836, 19.9836, 19.98365, 19.98367, 
    19.98374, 19.98379, 19.98383, 19.98382, 19.98378, 19.98369, 19.98361, 
    19.98363, 19.98357, 19.98373, 19.98366, 19.98369, 19.98362, 19.98376, 
    19.98364, 19.9838, 19.98378, 19.98374, 19.98366, 19.98364, 19.98362, 
    19.98363, 19.98369, 19.9837, 19.98374, 19.98375, 19.98379, 19.98381, 
    19.98379, 19.98376, 19.98369, 19.98363, 19.98355, 19.98354, 19.98346, 
    19.98352, 19.98341, 19.98351, 19.98334, 19.98363, 19.98351, 19.98374, 
    19.98371, 19.98367, 19.98357, 19.98362, 19.98356, 19.9837, 19.98377, 
    19.98379, 19.98383, 19.98379, 19.9838, 19.98376, 19.98377, 19.98369, 
    19.98373, 19.9836, 19.98356, 19.98343, 19.98334, 19.98326, 19.98322, 
    19.98321, 19.98321,
  19.98571, 19.98564, 19.98565, 19.9856, 19.98563, 19.98559, 19.98569, 
    19.98564, 19.98567, 19.9857, 19.98549, 19.9856, 19.98539, 19.98545, 
    19.98529, 19.9854, 19.98527, 19.98529, 19.98522, 19.98524, 19.98514, 
    19.98521, 19.98509, 19.98516, 19.98515, 19.98521, 19.98558, 19.98551, 
    19.98558, 19.98557, 19.98557, 19.98563, 19.98565, 19.98571, 19.9857, 
    19.98566, 19.98557, 19.9856, 19.98552, 19.98552, 19.98543, 19.98547, 
    19.98532, 19.98536, 19.98524, 19.98527, 19.98524, 19.98525, 19.98524, 
    19.98529, 19.98527, 19.98531, 19.98546, 19.98542, 19.98555, 19.98564, 
    19.98569, 19.98573, 19.98572, 19.98571, 19.98566, 19.98561, 19.98557, 
    19.98554, 19.98552, 19.98544, 19.9854, 19.98531, 19.98533, 19.9853, 
    19.98527, 19.98523, 19.98524, 19.98522, 19.9853, 19.98524, 19.98534, 
    19.98531, 19.98551, 19.98559, 19.98562, 19.98565, 19.98572, 19.98567, 
    19.98569, 19.98565, 19.98562, 19.98563, 19.98554, 19.98558, 19.9854, 
    19.98548, 19.98528, 19.98532, 19.98527, 19.98529, 19.98524, 19.98529, 
    19.98521, 19.98519, 19.9852, 19.98516, 19.98529, 19.98524, 19.98563, 
    19.98563, 19.98562, 19.98567, 19.98567, 19.98571, 19.98567, 19.98566, 
    19.98561, 19.98559, 19.98557, 19.98552, 19.98546, 19.98538, 19.98532, 
    19.98528, 19.98531, 19.98528, 19.98531, 19.98532, 19.9852, 19.98527, 
    19.98516, 19.98517, 19.98522, 19.98517, 19.98563, 19.98564, 19.98569, 
    19.98565, 19.98572, 19.98568, 19.98566, 19.98558, 19.98556, 19.98554, 
    19.98551, 19.98547, 19.98539, 19.98533, 19.98527, 19.98528, 19.98528, 
    19.98526, 19.98529, 19.98526, 19.98525, 19.98527, 19.98517, 19.9852, 
    19.98517, 19.98519, 19.98564, 19.98561, 19.98563, 19.9856, 19.98562, 
    19.98555, 19.98553, 19.98543, 19.98547, 19.9854, 19.98546, 19.98545, 
    19.9854, 19.98546, 19.98533, 19.98542, 19.98526, 19.98535, 19.98526, 
    19.98527, 19.98524, 19.98522, 19.98519, 19.98513, 19.98515, 19.9851, 
    19.98558, 19.98555, 19.98556, 19.98553, 19.9855, 19.98545, 19.98538, 
    19.9854, 19.98535, 19.98534, 19.98542, 19.98537, 19.98553, 19.98551, 
    19.98552, 19.98558, 19.9854, 19.98549, 19.98532, 19.98537, 19.98522, 
    19.9853, 19.98515, 19.98509, 19.98503, 19.98497, 19.98554, 19.98556, 
    19.98552, 19.98547, 19.98543, 19.98537, 19.98536, 19.98535, 19.98532, 
    19.9853, 19.98535, 19.98529, 19.9855, 19.98539, 19.98556, 19.98551, 
    19.98548, 19.98549, 19.98541, 19.98539, 19.98531, 19.98535, 19.98511, 
    19.98522, 19.98492, 19.985, 19.98556, 19.98554, 19.98545, 19.98549, 
    19.98536, 19.98533, 19.98531, 19.98528, 19.98527, 19.98525, 19.98528, 
    19.98525, 19.98537, 19.98532, 19.98545, 19.98542, 19.98544, 19.98545, 
    19.9854, 19.98535, 19.98534, 19.98533, 19.98528, 19.98536, 19.98509, 
    19.98526, 19.98551, 19.98546, 19.98545, 19.98547, 19.98534, 19.98538, 
    19.98525, 19.98529, 19.98523, 19.98526, 19.98526, 19.9853, 19.98532, 
    19.98538, 19.98543, 19.98547, 19.98546, 19.98542, 19.98534, 19.98527, 
    19.98529, 19.98524, 19.98537, 19.98532, 19.98534, 19.98528, 19.98541, 
    19.9853, 19.98543, 19.98542, 19.98539, 19.98531, 19.98529, 19.98528, 
    19.98529, 19.98534, 19.98535, 19.98539, 19.9854, 19.98542, 19.98545, 
    19.98543, 19.9854, 19.98534, 19.98528, 19.98522, 19.9852, 19.98513, 
    19.98519, 19.98509, 19.98518, 19.98503, 19.98529, 19.98518, 19.98538, 
    19.98536, 19.98532, 19.98523, 19.98528, 19.98522, 19.98535, 19.98541, 
    19.98543, 19.98546, 19.98543, 19.98543, 19.9854, 19.98541, 19.98534, 
    19.98538, 19.98526, 19.98522, 19.9851, 19.98503, 19.98496, 19.98493, 
    19.98491, 19.98491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222453, 0.7222428, 0.7222432, 0.7222412, 0.7222424, 0.722241, 0.7222448, 
    0.7222427, 0.722244, 0.722245, 0.7222373, 0.7222411, 0.7222332, 
    0.7222357, 0.7222295, 0.7222337, 0.7222287, 0.7222297, 0.7222268, 
    0.7222276, 0.722224, 0.7222264, 0.7222221, 0.7222246, 0.7222242, 
    0.7222265, 0.7222403, 0.7222378, 0.7222405, 0.7222401, 0.7222403, 
    0.7222423, 0.7222434, 0.7222455, 0.7222451, 0.7222435, 0.72224, 
    0.7222412, 0.7222381, 0.7222382, 0.7222348, 0.7222363, 0.7222307, 
    0.7222323, 0.7222276, 0.7222288, 0.7222276, 0.722228, 0.7222276, 
    0.7222294, 0.7222286, 0.7222301, 0.722236, 0.7222343, 0.7222395, 
    0.7222426, 0.7222447, 0.7222462, 0.7222459, 0.7222456, 0.7222435, 
    0.7222416, 0.7222401, 0.7222392, 0.7222382, 0.7222353, 0.7222338, 
    0.7222303, 0.722231, 0.7222299, 0.7222289, 0.7222272, 0.7222275, 
    0.7222267, 0.7222299, 0.7222278, 0.7222313, 0.7222303, 0.7222379, 
    0.7222409, 0.7222421, 0.7222431, 0.7222458, 0.722244, 0.7222447, 
    0.722243, 0.7222419, 0.7222424, 0.7222391, 0.7222404, 0.7222337, 
    0.7222366, 0.722229, 0.7222308, 0.7222286, 0.7222297, 0.7222278, 
    0.7222295, 0.7222264, 0.7222258, 0.7222263, 0.7222245, 0.7222296, 
    0.7222276, 0.7222425, 0.7222424, 0.7222419, 0.7222437, 0.7222438, 
    0.7222455, 0.722244, 0.7222434, 0.7222418, 0.7222409, 0.72224, 0.7222381, 
    0.7222359, 0.7222329, 0.7222307, 0.7222292, 0.7222301, 0.7222294, 
    0.7222303, 0.7222306, 0.722226, 0.7222286, 0.7222248, 0.722225, 
    0.7222267, 0.722225, 0.7222423, 0.7222428, 0.7222446, 0.7222432, 
    0.7222457, 0.7222443, 0.7222435, 0.7222404, 0.7222397, 0.7222391, 
    0.7222378, 0.7222363, 0.7222335, 0.722231, 0.7222288, 0.722229, 
    0.7222289, 0.7222285, 0.7222297, 0.7222282, 0.722228, 0.7222286, 
    0.722225, 0.722226, 0.722225, 0.7222257, 0.7222427, 0.7222418, 0.7222422, 
    0.7222414, 0.722242, 0.7222393, 0.7222385, 0.7222347, 0.7222363, 
    0.7222338, 0.722236, 0.7222357, 0.7222338, 0.7222359, 0.7222311, 
    0.7222344, 0.7222284, 0.7222316, 0.7222282, 0.7222288, 0.7222278, 
    0.7222269, 0.7222257, 0.7222236, 0.7222241, 0.7222223, 0.7222406, 
    0.7222394, 0.7222396, 0.7222384, 0.7222375, 0.7222357, 0.7222328, 
    0.7222339, 0.7222319, 0.7222314, 0.7222345, 0.7222326, 0.7222387, 
    0.7222377, 0.7222383, 0.7222404, 0.7222337, 0.7222371, 0.7222307, 
    0.7222326, 0.722227, 0.7222298, 0.7222244, 0.722222, 0.7222199, 
    0.7222173, 0.7222388, 0.7222396, 0.7222382, 0.7222364, 0.7222347, 
    0.7222325, 0.7222322, 0.7222318, 0.7222307, 0.7222298, 0.7222316, 
    0.7222295, 0.7222375, 0.7222333, 0.7222399, 0.7222379, 0.7222365, 
    0.7222371, 0.722234, 0.7222333, 0.7222303, 0.7222318, 0.7222226, 
    0.7222267, 0.7222154, 0.7222186, 0.7222399, 0.7222388, 0.7222354, 
    0.7222371, 0.7222323, 0.7222311, 0.7222302, 0.7222289, 0.7222288, 
    0.7222281, 0.7222293, 0.7222282, 0.7222325, 0.7222306, 0.7222358, 
    0.7222345, 0.7222351, 0.7222357, 0.7222337, 0.7222316, 0.7222316, 
    0.7222309, 0.722229, 0.7222323, 0.7222221, 0.7222284, 0.7222378, 
    0.7222359, 0.7222356, 0.7222363, 0.7222313, 0.7222331, 0.7222281, 
    0.7222295, 0.7222273, 0.7222283, 0.7222285, 0.72223, 0.7222308, 0.722233, 
    0.7222348, 0.7222362, 0.7222359, 0.7222343, 0.7222315, 0.7222288, 
    0.7222294, 0.7222275, 0.7222326, 0.7222304, 0.7222313, 0.7222291, 
    0.7222339, 0.7222298, 0.722235, 0.7222345, 0.7222331, 0.7222303, 
    0.7222297, 0.7222291, 0.7222294, 0.7222314, 0.7222317, 0.7222332, 
    0.7222335, 0.7222346, 0.7222355, 0.7222347, 0.7222338, 0.7222314, 
    0.7222292, 0.7222269, 0.7222263, 0.7222235, 0.7222258, 0.7222221, 
    0.7222252, 0.7222198, 0.7222296, 0.7222253, 0.7222331, 0.7222322, 
    0.7222307, 0.7222273, 0.7222291, 0.7222269, 0.7222317, 0.7222342, 
    0.7222349, 0.7222361, 0.7222349, 0.722235, 0.7222338, 0.7222342, 
    0.7222313, 0.7222329, 0.7222285, 0.722227, 0.7222225, 0.7222198, 
    0.722217, 0.7222158, 0.7222154, 0.7222152 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  1.027984e-20, 1.027984e-20, -2.006177e-36, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 2.569961e-20, 5.653913e-20, 2.055969e-20, 
    -2.006177e-36, 3.597945e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    3.083953e-20, 5.139921e-21, 5.139921e-21, 4.111937e-20, 3.597945e-20, 
    -3.083953e-20, 3.597945e-20, -1.027984e-20, -2.055969e-20, -1.541976e-20, 
    5.139921e-21, 2.055969e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -3.597945e-20, -1.541976e-20, -3.083953e-20, -1.541976e-20, 2.569961e-20, 
    3.597945e-20, 0, -1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 1.541976e-20, 1.027984e-20, 0, 
    -2.055969e-20, 0, 1.541976e-20, 0, 0, 2.055969e-20, 5.139921e-21, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -2.569961e-20, -1.027984e-20, 
    -4.111937e-20, -3.597945e-20, -2.569961e-20, -5.139921e-21, 1.027984e-20, 
    -1.541976e-20, -1.541976e-20, 3.597945e-20, -1.027984e-20, -1.541976e-20, 
    1.541976e-20, 1.541976e-20, -5.139921e-20, -2.055969e-20, 5.139921e-21, 
    0, 5.139921e-21, 5.139921e-21, 3.597945e-20, -5.139921e-21, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    1.541976e-20, 2.569961e-20, 4.625929e-20, 3.083953e-20, 0, 1.027984e-20, 
    -4.111937e-20, 2.569961e-20, 1.541976e-20, -5.139921e-21, 2.569961e-20, 
    3.083953e-20, 1.541976e-20, 1.027984e-20, 1.541976e-20, 0, 2.055969e-20, 
    -1.027984e-20, 1.541976e-20, 1.027984e-20, -5.139921e-21, 2.055969e-20, 
    4.625929e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -1.541976e-20, -2.055969e-20, -5.139921e-21, 
    -2.569961e-20, 2.569961e-20, 5.139921e-21, 2.055969e-20, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, -2.569961e-20, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 2.569961e-20, 
    -4.111937e-20, 1.027984e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    3.597945e-20, 2.006177e-36, 2.055969e-20, 1.027984e-20, -3.597945e-20, 
    -2.006177e-36, -2.006177e-36, -2.569961e-20, 1.027984e-20, 1.027984e-20, 
    0, 1.027984e-20, -1.027984e-20, 2.006177e-36, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 3.083953e-20, 1.027984e-20, 0, 
    -5.139921e-21, 0, 1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.006177e-36, 1.541976e-20, -1.027984e-20, -2.569961e-20, 
    -1.027984e-20, 5.139921e-21, 2.055969e-20, 0, 3.597945e-20, 
    -1.541976e-20, 0, -2.569961e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -3.597945e-20, -1.541976e-20, 0, 
    5.139921e-21, -2.569961e-20, -2.569961e-20, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 4.111937e-20, 1.027984e-20, -2.055969e-20, -2.055969e-20, 
    2.055969e-20, 0, -2.006177e-36, -5.139921e-20, 2.055969e-20, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, 2.055969e-20, -2.569961e-20, 
    -3.083953e-20, -2.006177e-36, 5.139921e-21, 0, -2.055969e-20, 
    -1.541976e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, -2.006177e-36, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, -1.027984e-20, -4.111937e-20, -1.027984e-20, 2.055969e-20, 
    1.027984e-20, 3.083953e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 0, 2.006177e-36, 5.139921e-21, 
    -2.055969e-20, -1.027984e-20, -2.569961e-20, 5.139921e-21, -4.111937e-20, 
    -3.083953e-20, -1.541976e-20, 5.139921e-21, -4.111937e-20, 3.083953e-20, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, -2.569961e-20, 2.006177e-36, 
    -5.139921e-21, -1.541976e-20, 2.569961e-20, -5.139921e-21, 0, 
    -2.055969e-20, 1.541976e-20, -3.597945e-20, -2.569961e-20, 1.541976e-20, 
    -2.569961e-20, 1.541976e-20, 1.027984e-20, -2.055969e-20, 2.006177e-36, 
    0, 1.541976e-20, 2.569961e-20, -5.139921e-21, -1.541976e-20, 
    1.541976e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, -2.006177e-36, 
    -5.139921e-21, -3.083953e-20, -1.541976e-20, -3.597945e-20, 0, 
    1.027984e-20, -3.083953e-20, 2.569961e-20, 5.139921e-21, 1.541976e-20, 0, 
    -1.541976e-20, 1.541976e-20, 1.541976e-20, 1.541976e-20, -2.006177e-36, 
    -1.027984e-20, 1.541976e-20, 5.139921e-21, 0, -1.027984e-20, 0, 
    2.569961e-20, 4.111937e-20, 2.006177e-36, -2.055969e-20, 0, 1.541976e-20, 
    1.027984e-20, 3.083953e-20, -1.027984e-20, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, 2.569961e-20, 1.541976e-20, 1.027984e-20, 
    2.569961e-20, -2.006177e-36, -2.569961e-20, -1.541976e-20, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, -2.055969e-20, 5.139921e-21, 2.055969e-20, 
    5.139921e-21, 2.055969e-20, 0, -2.055969e-20, -2.569961e-20, 
    -1.541976e-20, 0, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    2.569961e-20, -1.541976e-20, -2.055969e-20, -2.569961e-20, 5.139921e-21, 
    3.597945e-20, 1.541976e-20, 5.139921e-21, -3.083953e-20,
  -1.541976e-20, -3.083953e-20, 1.541976e-20, -4.111937e-20, -3.083953e-20, 
    -1.541976e-20, 2.055969e-20, 2.569961e-20, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -1.541976e-20, 5.139921e-21, 
    2.055969e-20, -2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 2.569961e-20, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, -5.139921e-21, 2.569961e-20, 
    -1.027984e-20, 2.055969e-20, 1.027984e-20, 0, 1.027984e-20, 3.083953e-20, 
    -1.027984e-20, -5.139921e-21, 2.055969e-20, 2.006177e-36, -5.139921e-21, 
    5.139921e-21, 3.083953e-20, -2.006177e-36, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, 0, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -2.055969e-20, -1.027984e-20, 2.055969e-20, 5.139921e-21, 5.139921e-21, 
    -5.139921e-20, 1.027984e-20, -3.083953e-20, -3.597945e-20, -3.083953e-20, 
    0, 2.055969e-20, 5.139921e-21, -1.027984e-20, -3.083953e-20, 0, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, -2.055969e-20, 
    -2.055969e-20, 3.597945e-20, -5.139921e-21, -3.597945e-20, 0, 
    -5.139921e-21, 0, -1.027984e-20, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, 0, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 3.597945e-20, -5.139921e-21, 5.139921e-21, 
    3.597945e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    0, -5.139921e-21, -5.139921e-21, 0, -2.055969e-20, 5.139921e-21, 
    2.055969e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.027984e-20, 0, 0, 
    -1.541976e-20, -1.541976e-20, 2.569961e-20, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 3.597945e-20, 5.139921e-21, 3.083953e-20, 0, 
    -1.027984e-20, -5.139921e-21, -2.055969e-20, 1.027984e-20, 1.027984e-20, 
    0, 1.541976e-20, 5.139921e-21, -1.541976e-20, 0, -1.027984e-20, 0, 
    5.139921e-21, -3.083953e-20, -2.006177e-36, -1.027984e-20, -1.027984e-20, 
    -2.006177e-36, -5.139921e-21, 5.139921e-20, 5.139921e-21, -1.027984e-20, 
    0, -1.541976e-20, -1.541976e-20, 1.541976e-20, -1.027984e-20, 
    -2.055969e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, -1.027984e-20, -2.569961e-20, 1.027984e-20, 
    2.006177e-36, -1.027984e-20, -2.006177e-36, 1.027984e-20, -2.055969e-20, 
    2.006177e-36, 0, -1.541976e-20, 2.569961e-20, 1.027984e-20, 0, 
    2.569961e-20, -2.006177e-36, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 0, 
    2.569961e-20, -2.006177e-36, 1.541976e-20, 0, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, -2.055969e-20, 2.569961e-20, 
    -1.541976e-20, 2.055969e-20, 1.541976e-20, 2.006177e-36, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, 2.055969e-20, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    3.083953e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 3.083953e-20, -2.055969e-20, 5.139921e-21, 
    -1.541976e-20, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -2.006177e-36, 5.139921e-21, 1.027984e-20, 1.541976e-20, 1.027984e-20, 0, 
    -2.006177e-36, -5.139921e-21, -1.541976e-20, -1.541976e-20, 0, 
    4.111937e-20, 2.569961e-20, 1.541976e-20, 1.541976e-20, 2.055969e-20, 0, 
    2.055969e-20, -1.027984e-20, -2.569961e-20, -2.006177e-36, -3.083953e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 2.006177e-36, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, 2.055969e-20, 2.055969e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 2.569961e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, -3.083953e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, -1.541976e-20, -3.597945e-20, 
    2.006177e-36, 1.541976e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, 
    2.006177e-36, -2.569961e-20, 1.541976e-20, 0, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -2.055969e-20, -4.111937e-20, -1.541976e-20, 2.055969e-20, 
    -2.055969e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, -1.541976e-20, 
    1.027984e-20, 2.569961e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 1.027984e-20, 
    -1.541976e-20, 1.027984e-20, 0, -3.083953e-20, -3.083953e-20, 0, 
    5.139921e-21, -2.569961e-20, -1.027984e-20, 2.006177e-36, -1.027984e-20, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 0, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, -2.055969e-20, 
    1.027984e-20, 2.569961e-20, -1.027984e-20, -2.006177e-36, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20,
  -1.027984e-20, 2.055969e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, 5.139921e-21, -3.083953e-20, 
    -2.569961e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -3.083953e-20, 2.006177e-36, -5.139921e-21, 0, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, 2.055969e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-20, -2.569961e-20, 
    -1.027984e-20, 0, 0, 5.139921e-21, -2.006177e-36, 1.541976e-20, 
    2.569961e-20, -3.083953e-20, 1.027984e-20, -1.541976e-20, -2.055969e-20, 
    1.027984e-20, -5.139921e-21, 0, -5.139921e-21, 2.569961e-20, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, 2.055969e-20, 1.541976e-20, 
    5.139921e-21, -2.006177e-36, -1.027984e-20, -1.027984e-20, -2.055969e-20, 
    2.569961e-20, 4.111937e-20, 1.541976e-20, -1.541976e-20, -2.006177e-36, 
    1.541976e-20, -2.569961e-20, 2.055969e-20, -1.027984e-20, 0, 
    -2.055969e-20, 1.027984e-20, 0, -2.055969e-20, -2.055969e-20, 
    -1.541976e-20, 1.027984e-20, 3.083953e-20, -2.055969e-20, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, 0, -3.083953e-20, 
    -3.083953e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 1.541976e-20, 
    -3.083953e-20, -1.541976e-20, 1.541976e-20, -1.541976e-20, -1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-20, 
    -3.597945e-20, -2.006177e-36, -5.139921e-21, 5.139921e-21, -3.597945e-20, 
    1.541976e-20, -3.083953e-20, 1.541976e-20, -2.055969e-20, 2.006177e-36, 
    2.569961e-20, 5.139921e-21, 2.055969e-20, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -2.055969e-20, 0, -1.027984e-20, 0, 5.139921e-21, 
    2.055969e-20, -4.625929e-20, -1.027984e-20, 5.139921e-21, 2.569961e-20, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 2.569961e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -3.083953e-20, 1.027984e-20, 1.027984e-20, 
    4.111937e-20, -1.027984e-20, 5.139921e-21, -2.006177e-36, 3.083953e-20, 
    1.541976e-20, 1.541976e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 
    -2.569961e-20, -1.027984e-20, 0, -4.625929e-20, 2.006177e-36, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, 1.027984e-20, 0, 2.055969e-20, 
    -5.139921e-21, -1.027984e-20, 3.083953e-20, 2.055969e-20, 5.139921e-21, 
    0, 1.027984e-20, -1.541976e-20, 1.027984e-20, -2.569961e-20, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, 2.006177e-36, 
    -2.006177e-36, -5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 0, -1.541976e-20, 
    -2.569961e-20, 1.541976e-20, 1.027984e-20, 2.569961e-20, 3.083953e-20, 
    1.027984e-20, 0, 2.569961e-20, 1.027984e-20, -5.139921e-21, 
    -2.006177e-36, 3.083953e-20, -1.027984e-20, -1.541976e-20, -1.541976e-20, 
    -2.055969e-20, 2.055969e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 2.569961e-20, 2.055969e-20, 2.006177e-36, 
    0, -2.055969e-20, 1.541976e-20, -3.083953e-20, -1.027984e-20, 
    2.006177e-36, 2.569961e-20, 2.055969e-20, 2.055969e-20, 1.541976e-20, 
    -2.055969e-20, -1.027984e-20, 2.055969e-20, 1.541976e-20, 2.055969e-20, 
    2.055969e-20, 3.083953e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    1.027984e-20, 0, -2.569961e-20, -3.083953e-20, 1.541976e-20, 
    3.597945e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -2.055969e-20, 0, -2.055969e-20, -1.541976e-20, 5.139921e-21, 
    1.027984e-20, -2.055969e-20, 0, -5.139921e-21, 1.541976e-20, 
    1.027984e-20, 0, 0, -1.027984e-20, 2.006177e-36, 2.006177e-36, 
    2.006177e-36, -2.006177e-36, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -3.083953e-20, 4.111937e-20, 5.139921e-21, -5.139921e-21, 
    3.083953e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, -2.569961e-20, 
    2.055969e-20, -5.139921e-21, 2.569961e-20, -1.027984e-20, 1.027984e-20, 
    3.597945e-20, 5.139921e-21, 2.006177e-36, 3.597945e-20, -1.541976e-20, 
    1.027984e-20, 0, 2.055969e-20, 1.541976e-20, -5.139921e-21, 
    -1.541976e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-20, 0, -1.027984e-20, 0, 5.139921e-21, 
    2.055969e-20, 2.055969e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, 3.597945e-20, -2.569961e-20, 
    1.027984e-20, -2.055969e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -2.006177e-36, 2.569961e-20, -1.027984e-20, 2.569961e-20, 5.139921e-21, 
    0, -1.027984e-20, 1.541976e-20, -2.006177e-36, 0, -5.139921e-21, 
    -2.006177e-36, 5.139921e-21, -1.027984e-20, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, -1.027984e-20, 0, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 0, 2.055969e-20, 2.006177e-36, 2.006177e-36, 1.027984e-20, 
    -3.083953e-20, -3.083953e-20, -1.541976e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21,
  2.569961e-20, -1.027984e-20, 0, -5.139921e-21, 0, 1.541976e-20, 
    2.055969e-20, 3.083953e-20, -2.055969e-20, 0, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.006177e-36, 2.055969e-20, 
    -1.027984e-20, 2.006177e-36, 2.569961e-20, 5.653913e-20, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -2.055969e-20, -2.006177e-36, 5.139921e-21, 
    -1.541976e-20, 2.055969e-20, -2.006177e-36, -1.541976e-20, 1.027984e-20, 
    -1.541976e-20, -2.055969e-20, 2.055969e-20, 1.541976e-20, 1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -3.083953e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, -1.541976e-20, 
    -2.569961e-20, -2.569961e-20, 5.139921e-21, 0, -1.027984e-20, 0, 
    -5.139921e-21, -4.111937e-20, -3.597945e-20, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, 2.569961e-20, -5.139921e-20, 5.139921e-21, -2.006177e-36, 
    1.027984e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, -4.111937e-20, 
    2.055969e-20, -5.139921e-21, -3.597945e-20, 1.027984e-20, -1.027984e-20, 
    2.569961e-20, 1.027984e-20, -1.541976e-20, -2.055969e-20, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 1.541976e-20, -3.083953e-20, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 0, -2.569961e-20, -3.083953e-20, 1.027984e-20, 
    -1.027984e-20, 1.541976e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, 
    -2.006177e-36, 1.027984e-20, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    -5.139921e-21, -2.055969e-20, -4.111937e-20, -3.083953e-20, 2.055969e-20, 
    1.541976e-20, 5.139921e-21, 3.597945e-20, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, 1.541976e-20, 0, -2.055969e-20, -2.055969e-20, 
    -2.569961e-20, -2.569961e-20, 1.027984e-20, 2.569961e-20, 5.139921e-21, 
    3.083953e-20, 2.006177e-36, 0, 0, -2.055969e-20, 2.055969e-20, 
    1.541976e-20, 1.541976e-20, 5.653913e-20, 2.055969e-20, 2.055969e-20, 
    -4.111937e-20, 5.139921e-20, 3.597945e-20, 5.139921e-21, -1.027984e-20, 
    -1.541976e-20, 3.597945e-20, 0, -1.541976e-20, -2.055969e-20, 
    2.006177e-36, -2.055969e-20, 5.139921e-21, 2.569961e-20, -1.541976e-20, 
    5.139921e-21, -3.083953e-20, -1.027984e-20, -2.055969e-20, -3.597945e-20, 
    1.541976e-20, -2.055969e-20, 3.597945e-20, 0, -1.027984e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -2.055969e-20, -2.569961e-20, 1.541976e-20, 
    5.139921e-21, -1.541976e-20, 2.055969e-20, -2.569961e-20, -1.027984e-20, 
    -1.541976e-20, -2.055969e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, -3.083953e-20, 3.597945e-20, 
    5.139921e-21, 0, -1.541976e-20, 1.027984e-20, -1.027984e-20, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, 1.541976e-20, -3.083953e-20, 
    -5.139921e-21, 1.541976e-20, 1.541976e-20, -2.569961e-20, -1.027984e-20, 
    1.027984e-20, 4.111937e-20, 1.541976e-20, -3.597945e-20, -1.027984e-20, 
    1.027984e-20, 1.541976e-20, 1.027984e-20, -2.055969e-20, -2.055969e-20, 
    -1.027984e-20, 3.083953e-20, 0, 2.055969e-20, 2.569961e-20, 
    -2.569961e-20, 1.027984e-20, 5.139921e-21, -1.541976e-20, 2.055969e-20, 
    1.027984e-20, -3.597945e-20, -1.027984e-20, 0, 2.055969e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 3.083953e-20, 
    3.083953e-20, 5.139921e-21, 2.055969e-20, -3.083953e-20, -1.027984e-20, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    -1.027984e-20, -2.569961e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, 
    2.006177e-36, -1.541976e-20, 1.027984e-20, 2.569961e-20, 3.083953e-20, 
    1.541976e-20, -1.541976e-20, -1.541976e-20, -5.139921e-21, 3.597945e-20, 
    5.139921e-21, -4.111937e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, 
    3.597945e-20, -1.541976e-20, -1.027984e-20, -5.139921e-21, 2.055969e-20, 
    3.083953e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 1.541976e-20, 0, -2.055969e-20, 5.139921e-21, 
    2.055969e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 2.055969e-20, -2.055969e-20, -1.541976e-20, 2.569961e-20, 
    -2.006177e-36, 2.006177e-36, -2.569961e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, 2.569961e-20, 2.055969e-20, 5.139921e-21, 
    -2.569961e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    3.083953e-20, -5.139921e-21, -1.027984e-20, 0, 5.139921e-21, 
    5.139921e-20, 5.139921e-21, -4.111937e-20, -5.139921e-21, 1.027984e-20, 
    -1.541976e-20, 5.139921e-21, -2.055969e-20, -1.541976e-20, -5.139921e-21, 
    -1.027984e-20, -2.055969e-20, 5.139921e-21, -3.083953e-20, -1.027984e-20, 
    2.569961e-20, 2.006177e-36, 5.139921e-21, 2.006177e-36, 5.139921e-21, 
    -2.569961e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -2.569961e-20, -5.139921e-21, 3.083953e-20, -1.541976e-20, 1.541976e-20,
  -2.006177e-36, -1.027984e-20, -4.625929e-20, 1.027984e-20, 1.027984e-20, 
    -2.006177e-36, 5.139921e-21, 0, 1.027984e-20, -1.027984e-20, 0, 
    1.541976e-20, 1.027984e-20, -2.569961e-20, 0, 2.055969e-20, 
    -1.541976e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 2.006177e-36, 
    -5.139921e-21, 5.139921e-21, -3.597945e-20, -1.541976e-20, -1.027984e-20, 
    5.139921e-21, 2.569961e-20, -2.569961e-20, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 5.139921e-21, 2.569961e-20, -1.027984e-20, 
    5.139921e-21, 4.111937e-20, 5.139921e-21, 1.027984e-20, -2.055969e-20, 
    5.139921e-21, 2.006177e-36, -5.139921e-21, -1.027984e-20, -3.083953e-20, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, -2.055969e-20, 3.597945e-20, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    -4.625929e-20, 5.139921e-21, 2.055969e-20, 5.139921e-21, 1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -4.111937e-20, 5.139921e-21, 2.569961e-20, 
    2.569961e-20, -5.139921e-21, 5.139921e-21, -3.083953e-20, 1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, -2.569961e-20, 
    1.541976e-20, -2.569961e-20, -1.541976e-20, 3.083953e-20, 1.027984e-20, 
    0, 1.027984e-20, -3.597945e-20, 0, -2.006177e-36, 3.083953e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, 2.006177e-36, 3.083953e-20, 
    2.055969e-20, -5.139921e-21, 3.597945e-20, 1.027984e-20, 5.139921e-21, 
    2.055969e-20, -1.027984e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 2.006177e-36, 1.027984e-20, 0, -5.139921e-21, 
    5.139921e-21, 2.055969e-20, -1.541976e-20, 5.653913e-20, 5.139921e-21, 
    -5.139921e-21, -3.597945e-20, 5.139921e-21, -1.541976e-20, 2.055969e-20, 
    -3.083953e-20, 2.006177e-36, -5.139921e-21, -2.055969e-20, 2.055969e-20, 
    2.569961e-20, 4.111937e-20, 1.027984e-20, -2.055969e-20, -2.055969e-20, 
    1.541976e-20, 1.027984e-20, 2.055969e-20, -1.027984e-20, -1.541976e-20, 
    2.055969e-20, 1.027984e-20, 3.083953e-20, 2.569961e-20, -2.055969e-20, 
    5.139921e-21, -3.597945e-20, 1.541976e-20, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 1.027984e-20, -2.569961e-20, -1.541976e-20, 0, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, 2.055969e-20, 2.006177e-36, 3.083953e-20, 1.541976e-20, 
    2.006177e-36, 2.569961e-20, 0, 2.569961e-20, 2.569961e-20, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, 2.055969e-20, -1.027984e-20, 2.055969e-20, 
    1.027984e-20, -2.006177e-36, 5.139921e-21, 2.569961e-20, 2.006177e-36, 
    -5.139921e-21, 0, -5.139921e-21, 2.055969e-20, -5.139921e-21, 
    5.139921e-21, -2.569961e-20, 1.027984e-20, -2.006177e-36, -1.027984e-20, 
    2.055969e-20, -1.027984e-20, 0, 2.006177e-36, 2.569961e-20, 3.597945e-20, 
    2.055969e-20, -1.027984e-20, -3.597945e-20, 5.139921e-21, -3.597945e-20, 
    -3.597945e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 0, 
    -2.055969e-20, -2.055969e-20, 1.541976e-20, -1.541976e-20, 1.541976e-20, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    3.597945e-20, -2.055969e-20, 5.139921e-21, 1.027984e-20, 1.541976e-20, 0, 
    2.569961e-20, -5.139921e-21, 0, -2.006177e-36, -5.139921e-21, 
    2.006177e-36, 5.139921e-21, 0, -5.139921e-21, -5.139921e-20, 
    2.055969e-20, 2.569961e-20, 1.027984e-20, -2.569961e-20, 2.055969e-20, 
    1.541976e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, -2.006177e-36, 1.541976e-20, 
    3.083953e-20, -5.139921e-21, 2.569961e-20, 5.139921e-21, -5.139921e-21, 
    2.055969e-20, -2.055969e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 2.055969e-20, -3.597945e-20, 1.027984e-20, 3.597945e-20, 
    -1.027984e-20, -1.541976e-20, 1.541976e-20, -2.006177e-36, 1.541976e-20, 
    5.139921e-21, -2.006177e-36, 2.569961e-20, -1.541976e-20, -2.569961e-20, 
    2.006177e-36, 1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    4.111937e-20, 2.569961e-20, 5.139921e-21, 2.055969e-20, -1.027984e-20, 
    2.055969e-20, -1.027984e-20, 5.139921e-21, 2.569961e-20, -5.139921e-21, 
    -5.139921e-21, 0, 0, -3.083953e-20, 2.569961e-20, 1.541976e-20, 
    4.625929e-20, 2.055969e-20, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -3.083953e-20, -2.055969e-20, -1.541976e-20, 2.055969e-20, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, -3.083953e-20, 5.139921e-21, 
    3.083953e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -2.055969e-20, -5.139921e-21, -2.006177e-36, 2.569961e-20, 2.055969e-20, 
    -2.006177e-36, 5.139921e-21, 2.569961e-20, -2.055969e-20, -2.055969e-20, 
    -1.027984e-20, 0, 3.597945e-20, -2.055969e-20, -2.055969e-20, 
    -3.597945e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, -2.569961e-20, 
    5.139921e-21, -1.027984e-20,
  8.598664e-29, 8.598635e-29, 8.598641e-29, 8.598618e-29, 8.59863e-29, 
    8.598615e-29, 8.598658e-29, 8.598634e-29, 8.598649e-29, 8.598662e-29, 
    8.598573e-29, 8.598617e-29, 8.598527e-29, 8.598556e-29, 8.598485e-29, 
    8.598532e-29, 8.598476e-29, 8.598486e-29, 8.598454e-29, 8.598463e-29, 
    8.598422e-29, 8.59845e-29, 8.5984e-29, 8.598429e-29, 8.598424e-29, 
    8.598451e-29, 8.598608e-29, 8.598578e-29, 8.59861e-29, 8.598606e-29, 
    8.598607e-29, 8.59863e-29, 8.598642e-29, 8.598666e-29, 8.598662e-29, 
    8.598644e-29, 8.598604e-29, 8.598617e-29, 8.598583e-29, 8.598583e-29, 
    8.598545e-29, 8.598562e-29, 8.598498e-29, 8.598516e-29, 8.598463e-29, 
    8.598476e-29, 8.598463e-29, 8.598468e-29, 8.598463e-29, 8.598483e-29, 
    8.598475e-29, 8.598492e-29, 8.598559e-29, 8.598539e-29, 8.598598e-29, 
    8.598633e-29, 8.598657e-29, 8.598674e-29, 8.598671e-29, 8.598667e-29, 
    8.598643e-29, 8.598622e-29, 8.598606e-29, 8.598595e-29, 8.598584e-29, 
    8.598551e-29, 8.598533e-29, 8.598494e-29, 8.598501e-29, 8.598489e-29, 
    8.598478e-29, 8.598459e-29, 8.598462e-29, 8.598453e-29, 8.598489e-29, 
    8.598465e-29, 8.598505e-29, 8.598494e-29, 8.598581e-29, 8.598613e-29, 
    8.598627e-29, 8.59864e-29, 8.598669e-29, 8.598649e-29, 8.598657e-29, 
    8.598638e-29, 8.598625e-29, 8.598631e-29, 8.598594e-29, 8.598609e-29, 
    8.598532e-29, 8.598565e-29, 8.598479e-29, 8.5985e-29, 8.598474e-29, 
    8.598487e-29, 8.598465e-29, 8.598485e-29, 8.59845e-29, 8.598442e-29, 
    8.598448e-29, 8.598427e-29, 8.598486e-29, 8.598463e-29, 8.598632e-29, 
    8.598631e-29, 8.598626e-29, 8.598646e-29, 8.598648e-29, 8.598666e-29, 
    8.598649e-29, 8.598643e-29, 8.598625e-29, 8.598614e-29, 8.598604e-29, 
    8.598582e-29, 8.598557e-29, 8.598523e-29, 8.598498e-29, 8.598482e-29, 
    8.598492e-29, 8.598483e-29, 8.598493e-29, 8.598498e-29, 8.598445e-29, 
    8.598475e-29, 8.59843e-29, 8.598433e-29, 8.598453e-29, 8.598433e-29, 
    8.59863e-29, 8.598636e-29, 8.598655e-29, 8.59864e-29, 8.598668e-29, 
    8.598652e-29, 8.598643e-29, 8.598609e-29, 8.598601e-29, 8.598593e-29, 
    8.59858e-29, 8.598562e-29, 8.59853e-29, 8.598502e-29, 8.598477e-29, 
    8.598479e-29, 8.598478e-29, 8.598473e-29, 8.598486e-29, 8.59847e-29, 
    8.598468e-29, 8.598475e-29, 8.598433e-29, 8.598445e-29, 8.598433e-29, 
    8.598441e-29, 8.598634e-29, 8.598624e-29, 8.59863e-29, 8.59862e-29, 
    8.598627e-29, 8.598596e-29, 8.598587e-29, 8.598544e-29, 8.598562e-29, 
    8.598534e-29, 8.598559e-29, 8.598554e-29, 8.598533e-29, 8.598557e-29, 
    8.598504e-29, 8.598541e-29, 8.598473e-29, 8.598509e-29, 8.59847e-29, 
    8.598477e-29, 8.598465e-29, 8.598455e-29, 8.598442e-29, 8.598418e-29, 
    8.598423e-29, 8.598403e-29, 8.59861e-29, 8.598598e-29, 8.598599e-29, 
    8.598586e-29, 8.598576e-29, 8.598556e-29, 8.598522e-29, 8.598535e-29, 
    8.598512e-29, 8.598507e-29, 8.598542e-29, 8.59852e-29, 8.598589e-29, 
    8.598578e-29, 8.598585e-29, 8.598609e-29, 8.598532e-29, 8.598571e-29, 
    8.598498e-29, 8.598519e-29, 8.598456e-29, 8.598488e-29, 8.598426e-29, 
    8.5984e-29, 8.598375e-29, 8.598346e-29, 8.598591e-29, 8.5986e-29, 
    8.598584e-29, 8.598563e-29, 8.598544e-29, 8.598518e-29, 8.598515e-29, 
    8.59851e-29, 8.598498e-29, 8.598488e-29, 8.598509e-29, 8.598485e-29, 
    8.598575e-29, 8.598528e-29, 8.598603e-29, 8.59858e-29, 8.598565e-29, 
    8.598571e-29, 8.598536e-29, 8.598527e-29, 8.598494e-29, 8.598511e-29, 
    8.598406e-29, 8.598453e-29, 8.598324e-29, 8.59836e-29, 8.598603e-29, 
    8.598591e-29, 8.598551e-29, 8.59857e-29, 8.598516e-29, 8.598503e-29, 
    8.598492e-29, 8.598479e-29, 8.598477e-29, 8.598469e-29, 8.598482e-29, 
    8.59847e-29, 8.598518e-29, 8.598497e-29, 8.598556e-29, 8.598541e-29, 
    8.598548e-29, 8.598556e-29, 8.598533e-29, 8.598509e-29, 8.598508e-29, 
    8.598501e-29, 8.598479e-29, 8.598516e-29, 8.5984e-29, 8.598472e-29, 
    8.598578e-29, 8.598557e-29, 8.598554e-29, 8.598562e-29, 8.598504e-29, 
    8.598525e-29, 8.598469e-29, 8.598485e-29, 8.598459e-29, 8.598472e-29, 
    8.598474e-29, 8.598489e-29, 8.5985e-29, 8.598524e-29, 8.598545e-29, 
    8.598561e-29, 8.598557e-29, 8.598539e-29, 8.598507e-29, 8.598477e-29, 
    8.598483e-29, 8.598461e-29, 8.59852e-29, 8.598495e-29, 8.598505e-29, 
    8.59848e-29, 8.598535e-29, 8.598488e-29, 8.598547e-29, 8.598542e-29, 
    8.598525e-29, 8.598494e-29, 8.598487e-29, 8.598479e-29, 8.598484e-29, 
    8.598506e-29, 8.59851e-29, 8.598526e-29, 8.59853e-29, 8.598543e-29, 
    8.598553e-29, 8.598544e-29, 8.598534e-29, 8.598506e-29, 8.598482e-29, 
    8.598455e-29, 8.598448e-29, 8.598417e-29, 8.598442e-29, 8.5984e-29, 
    8.598436e-29, 8.598374e-29, 8.598486e-29, 8.598437e-29, 8.598525e-29, 
    8.598516e-29, 8.598498e-29, 8.598459e-29, 8.59848e-29, 8.598456e-29, 
    8.59851e-29, 8.598539e-29, 8.598546e-29, 8.59856e-29, 8.598546e-29, 
    8.598547e-29, 8.598533e-29, 8.598538e-29, 8.598506e-29, 8.598523e-29, 
    8.598474e-29, 8.598456e-29, 8.598405e-29, 8.598374e-29, 8.598342e-29, 
    8.598328e-29, 8.598324e-29, 8.598322e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.164952e-08, 1.170074e-08, 1.169078e-08, 1.173209e-08, 1.170917e-08, 
    1.173622e-08, 1.16599e-08, 1.170277e-08, 1.16754e-08, 1.165413e-08, 
    1.181225e-08, 1.173393e-08, 1.18936e-08, 1.184365e-08, 1.196912e-08, 
    1.188583e-08, 1.198592e-08, 1.196672e-08, 1.20245e-08, 1.200795e-08, 
    1.208186e-08, 1.203214e-08, 1.212017e-08, 1.206998e-08, 1.207783e-08, 
    1.20305e-08, 1.174969e-08, 1.18025e-08, 1.174656e-08, 1.175409e-08, 
    1.175071e-08, 1.170965e-08, 1.168895e-08, 1.16456e-08, 1.165347e-08, 
    1.168531e-08, 1.175748e-08, 1.173298e-08, 1.179472e-08, 1.179333e-08, 
    1.186206e-08, 1.183107e-08, 1.194659e-08, 1.191376e-08, 1.200864e-08, 
    1.198478e-08, 1.200752e-08, 1.200062e-08, 1.200761e-08, 1.197261e-08, 
    1.198761e-08, 1.195681e-08, 1.183687e-08, 1.187212e-08, 1.176699e-08, 
    1.170378e-08, 1.166178e-08, 1.163199e-08, 1.16362e-08, 1.164423e-08, 
    1.16855e-08, 1.172429e-08, 1.175386e-08, 1.177364e-08, 1.179313e-08, 
    1.185211e-08, 1.188333e-08, 1.195323e-08, 1.194062e-08, 1.196199e-08, 
    1.19824e-08, 1.201668e-08, 1.201104e-08, 1.202614e-08, 1.196142e-08, 
    1.200444e-08, 1.193343e-08, 1.195285e-08, 1.179843e-08, 1.173959e-08, 
    1.171458e-08, 1.169269e-08, 1.163944e-08, 1.167621e-08, 1.166172e-08, 
    1.169621e-08, 1.171812e-08, 1.170728e-08, 1.177418e-08, 1.174817e-08, 
    1.188518e-08, 1.182617e-08, 1.198002e-08, 1.194321e-08, 1.198885e-08, 
    1.196556e-08, 1.200546e-08, 1.196955e-08, 1.203176e-08, 1.204531e-08, 
    1.203605e-08, 1.207161e-08, 1.196756e-08, 1.200752e-08, 1.170698e-08, 
    1.170875e-08, 1.171698e-08, 1.168078e-08, 1.167857e-08, 1.164539e-08, 
    1.167491e-08, 1.168748e-08, 1.171939e-08, 1.173827e-08, 1.175621e-08, 
    1.179566e-08, 1.183972e-08, 1.190133e-08, 1.194559e-08, 1.197526e-08, 
    1.195707e-08, 1.197313e-08, 1.195518e-08, 1.194676e-08, 1.204023e-08, 
    1.198775e-08, 1.20665e-08, 1.206214e-08, 1.20265e-08, 1.206263e-08, 
    1.170999e-08, 1.169982e-08, 1.16645e-08, 1.169214e-08, 1.164178e-08, 
    1.166997e-08, 1.168618e-08, 1.174872e-08, 1.176246e-08, 1.17752e-08, 
    1.180036e-08, 1.183266e-08, 1.188931e-08, 1.19386e-08, 1.198359e-08, 
    1.198029e-08, 1.198146e-08, 1.199151e-08, 1.196661e-08, 1.19956e-08, 
    1.200046e-08, 1.198774e-08, 1.206155e-08, 1.204047e-08, 1.206205e-08, 
    1.204831e-08, 1.170312e-08, 1.172024e-08, 1.171099e-08, 1.172838e-08, 
    1.171613e-08, 1.177062e-08, 1.178695e-08, 1.186339e-08, 1.183202e-08, 
    1.188195e-08, 1.183709e-08, 1.184504e-08, 1.188358e-08, 1.183952e-08, 
    1.193588e-08, 1.187055e-08, 1.19919e-08, 1.192666e-08, 1.199599e-08, 
    1.19834e-08, 1.200424e-08, 1.202291e-08, 1.204639e-08, 1.208973e-08, 
    1.207969e-08, 1.211593e-08, 1.174576e-08, 1.176796e-08, 1.176601e-08, 
    1.178924e-08, 1.180642e-08, 1.184366e-08, 1.19034e-08, 1.188093e-08, 
    1.192217e-08, 1.193045e-08, 1.18678e-08, 1.190627e-08, 1.178282e-08, 
    1.180277e-08, 1.179089e-08, 1.174751e-08, 1.188611e-08, 1.181498e-08, 
    1.194632e-08, 1.190779e-08, 1.202025e-08, 1.196432e-08, 1.207417e-08, 
    1.212113e-08, 1.216532e-08, 1.221697e-08, 1.178008e-08, 1.176499e-08, 
    1.1792e-08, 1.182937e-08, 1.186405e-08, 1.191014e-08, 1.191486e-08, 
    1.19235e-08, 1.194586e-08, 1.196467e-08, 1.192623e-08, 1.196939e-08, 
    1.180739e-08, 1.189229e-08, 1.175929e-08, 1.179934e-08, 1.182717e-08, 
    1.181496e-08, 1.187837e-08, 1.189331e-08, 1.195404e-08, 1.192265e-08, 
    1.210954e-08, 1.202685e-08, 1.225629e-08, 1.219217e-08, 1.175972e-08, 
    1.178002e-08, 1.185069e-08, 1.181707e-08, 1.191322e-08, 1.193689e-08, 
    1.195613e-08, 1.198072e-08, 1.198338e-08, 1.199795e-08, 1.197407e-08, 
    1.199701e-08, 1.191024e-08, 1.194902e-08, 1.184261e-08, 1.186851e-08, 
    1.18566e-08, 1.184353e-08, 1.188386e-08, 1.192683e-08, 1.192775e-08, 
    1.194153e-08, 1.198036e-08, 1.191361e-08, 1.212021e-08, 1.199262e-08, 
    1.180217e-08, 1.184128e-08, 1.184686e-08, 1.183171e-08, 1.193452e-08, 
    1.189727e-08, 1.199759e-08, 1.197048e-08, 1.201491e-08, 1.199283e-08, 
    1.198958e-08, 1.196123e-08, 1.194357e-08, 1.189897e-08, 1.186269e-08, 
    1.183391e-08, 1.18406e-08, 1.187221e-08, 1.192946e-08, 1.198362e-08, 
    1.197176e-08, 1.201153e-08, 1.190625e-08, 1.19504e-08, 1.193333e-08, 
    1.197782e-08, 1.188034e-08, 1.196336e-08, 1.185912e-08, 1.186826e-08, 
    1.189653e-08, 1.195339e-08, 1.196597e-08, 1.19794e-08, 1.197111e-08, 
    1.193091e-08, 1.192433e-08, 1.189584e-08, 1.188797e-08, 1.186627e-08, 
    1.18483e-08, 1.186472e-08, 1.188196e-08, 1.193093e-08, 1.197506e-08, 
    1.202317e-08, 1.203495e-08, 1.209117e-08, 1.20454e-08, 1.212092e-08, 
    1.205672e-08, 1.216786e-08, 1.196817e-08, 1.205483e-08, 1.189781e-08, 
    1.191473e-08, 1.194533e-08, 1.20155e-08, 1.197761e-08, 1.202192e-08, 
    1.192407e-08, 1.18733e-08, 1.186016e-08, 1.183566e-08, 1.186072e-08, 
    1.185869e-08, 1.188267e-08, 1.187497e-08, 1.193256e-08, 1.190162e-08, 
    1.19895e-08, 1.202157e-08, 1.211213e-08, 1.216765e-08, 1.222416e-08, 
    1.224911e-08, 1.22567e-08, 1.225988e-08 ;

 SOIL1N_TO_SOIL3N =
  1.382178e-10, 1.388257e-10, 1.387075e-10, 1.391978e-10, 1.389258e-10, 
    1.392469e-10, 1.38341e-10, 1.388498e-10, 1.38525e-10, 1.382725e-10, 
    1.401493e-10, 1.392197e-10, 1.411149e-10, 1.40522e-10, 1.420113e-10, 
    1.410226e-10, 1.422107e-10, 1.419828e-10, 1.426686e-10, 1.424721e-10, 
    1.433494e-10, 1.427593e-10, 1.438042e-10, 1.432085e-10, 1.433017e-10, 
    1.427399e-10, 1.394067e-10, 1.400336e-10, 1.393696e-10, 1.39459e-10, 
    1.394189e-10, 1.389314e-10, 1.386858e-10, 1.381713e-10, 1.382647e-10, 
    1.386426e-10, 1.394992e-10, 1.392084e-10, 1.399412e-10, 1.399247e-10, 
    1.407405e-10, 1.403727e-10, 1.417439e-10, 1.413542e-10, 1.424803e-10, 
    1.421971e-10, 1.424671e-10, 1.423852e-10, 1.424681e-10, 1.420527e-10, 
    1.422307e-10, 1.418652e-10, 1.404415e-10, 1.4086e-10, 1.396121e-10, 
    1.388618e-10, 1.383633e-10, 1.380097e-10, 1.380597e-10, 1.38155e-10, 
    1.386448e-10, 1.391053e-10, 1.394562e-10, 1.39691e-10, 1.399223e-10, 
    1.406224e-10, 1.40993e-10, 1.418227e-10, 1.41673e-10, 1.419266e-10, 
    1.421689e-10, 1.425758e-10, 1.425088e-10, 1.426881e-10, 1.419199e-10, 
    1.424305e-10, 1.415877e-10, 1.418182e-10, 1.399852e-10, 1.392868e-10, 
    1.3899e-10, 1.387302e-10, 1.380981e-10, 1.385346e-10, 1.383626e-10, 
    1.387719e-10, 1.39032e-10, 1.389034e-10, 1.396974e-10, 1.393887e-10, 
    1.410149e-10, 1.403145e-10, 1.421407e-10, 1.417037e-10, 1.422454e-10, 
    1.41969e-10, 1.424427e-10, 1.420164e-10, 1.427548e-10, 1.429156e-10, 
    1.428057e-10, 1.432278e-10, 1.419927e-10, 1.424671e-10, 1.388998e-10, 
    1.389208e-10, 1.390185e-10, 1.385888e-10, 1.385626e-10, 1.381688e-10, 
    1.385192e-10, 1.386684e-10, 1.390471e-10, 1.392712e-10, 1.394841e-10, 
    1.399524e-10, 1.404754e-10, 1.412067e-10, 1.41732e-10, 1.420842e-10, 
    1.418682e-10, 1.420589e-10, 1.418458e-10, 1.417459e-10, 1.428554e-10, 
    1.422324e-10, 1.431671e-10, 1.431154e-10, 1.426924e-10, 1.431212e-10, 
    1.389355e-10, 1.388148e-10, 1.383955e-10, 1.387236e-10, 1.381259e-10, 
    1.384605e-10, 1.386529e-10, 1.393952e-10, 1.395583e-10, 1.397095e-10, 
    1.400082e-10, 1.403915e-10, 1.410639e-10, 1.41649e-10, 1.42183e-10, 
    1.421439e-10, 1.421577e-10, 1.42277e-10, 1.419815e-10, 1.423255e-10, 
    1.423833e-10, 1.422323e-10, 1.431085e-10, 1.428581e-10, 1.431143e-10, 
    1.429513e-10, 1.38854e-10, 1.390572e-10, 1.389474e-10, 1.391538e-10, 
    1.390084e-10, 1.396551e-10, 1.39849e-10, 1.407563e-10, 1.403839e-10, 
    1.409765e-10, 1.404441e-10, 1.405385e-10, 1.409959e-10, 1.404729e-10, 
    1.416167e-10, 1.408413e-10, 1.422816e-10, 1.415073e-10, 1.423302e-10, 
    1.421807e-10, 1.424281e-10, 1.426497e-10, 1.429285e-10, 1.434429e-10, 
    1.433238e-10, 1.437539e-10, 1.393601e-10, 1.396236e-10, 1.396004e-10, 
    1.398762e-10, 1.400801e-10, 1.405221e-10, 1.412311e-10, 1.409645e-10, 
    1.41454e-10, 1.415522e-10, 1.408086e-10, 1.412652e-10, 1.397999e-10, 
    1.400367e-10, 1.398957e-10, 1.393809e-10, 1.41026e-10, 1.401817e-10, 
    1.417407e-10, 1.412833e-10, 1.426181e-10, 1.419543e-10, 1.432582e-10, 
    1.438156e-10, 1.443402e-10, 1.449533e-10, 1.397674e-10, 1.395883e-10, 
    1.399089e-10, 1.403525e-10, 1.407641e-10, 1.413112e-10, 1.413672e-10, 
    1.414697e-10, 1.417352e-10, 1.419584e-10, 1.415021e-10, 1.420144e-10, 
    1.400916e-10, 1.410993e-10, 1.395207e-10, 1.39996e-10, 1.403264e-10, 
    1.401814e-10, 1.409341e-10, 1.411114e-10, 1.418323e-10, 1.414596e-10, 
    1.43678e-10, 1.426965e-10, 1.4542e-10, 1.446589e-10, 1.395258e-10, 
    1.397668e-10, 1.406056e-10, 1.402065e-10, 1.413478e-10, 1.416287e-10, 
    1.41857e-10, 1.42149e-10, 1.421805e-10, 1.423535e-10, 1.4207e-10, 
    1.423423e-10, 1.413124e-10, 1.417726e-10, 1.405097e-10, 1.408171e-10, 
    1.406756e-10, 1.405205e-10, 1.409993e-10, 1.415093e-10, 1.415202e-10, 
    1.416837e-10, 1.421447e-10, 1.413524e-10, 1.438048e-10, 1.422903e-10, 
    1.400296e-10, 1.404938e-10, 1.405601e-10, 1.403803e-10, 1.416005e-10, 
    1.411584e-10, 1.423492e-10, 1.420274e-10, 1.425547e-10, 1.422927e-10, 
    1.422541e-10, 1.419176e-10, 1.41708e-10, 1.411787e-10, 1.407479e-10, 
    1.404063e-10, 1.404858e-10, 1.40861e-10, 1.415405e-10, 1.421833e-10, 
    1.420425e-10, 1.425147e-10, 1.41265e-10, 1.41789e-10, 1.415865e-10, 
    1.421146e-10, 1.409574e-10, 1.419429e-10, 1.407056e-10, 1.408141e-10, 
    1.411496e-10, 1.418246e-10, 1.419739e-10, 1.421333e-10, 1.420349e-10, 
    1.415578e-10, 1.414796e-10, 1.411414e-10, 1.410481e-10, 1.407904e-10, 
    1.405771e-10, 1.40772e-10, 1.409767e-10, 1.41558e-10, 1.420818e-10, 
    1.426529e-10, 1.427926e-10, 1.4346e-10, 1.429168e-10, 1.438132e-10, 
    1.430511e-10, 1.443703e-10, 1.419999e-10, 1.430287e-10, 1.411649e-10, 
    1.413657e-10, 1.417288e-10, 1.425618e-10, 1.421121e-10, 1.42638e-10, 
    1.414765e-10, 1.408739e-10, 1.40718e-10, 1.404271e-10, 1.407247e-10, 
    1.407005e-10, 1.409852e-10, 1.408937e-10, 1.415773e-10, 1.412101e-10, 
    1.422532e-10, 1.426338e-10, 1.437088e-10, 1.443678e-10, 1.450386e-10, 
    1.453348e-10, 1.454249e-10, 1.454626e-10 ;

 SOIL1N_vr =
  2.497417, 2.49741, 2.497412, 2.497406, 2.497409, 2.497406, 2.497416, 
    2.49741, 2.497414, 2.497416, 2.497396, 2.497406, 2.497385, 2.497391, 
    2.497375, 2.497386, 2.497373, 2.497375, 2.497368, 2.49737, 2.49736, 
    2.497367, 2.497355, 2.497362, 2.497361, 2.497367, 2.497404, 2.497397, 
    2.497404, 2.497403, 2.497404, 2.497409, 2.497412, 2.497418, 2.497416, 
    2.497412, 2.497403, 2.497406, 2.497398, 2.497398, 2.497389, 2.497393, 
    2.497378, 2.497382, 2.49737, 2.497373, 2.49737, 2.497371, 2.49737, 
    2.497375, 2.497373, 2.497377, 2.497392, 2.497388, 2.497402, 2.49741, 
    2.497416, 2.497419, 2.497419, 2.497418, 2.497412, 2.497407, 2.497403, 
    2.497401, 2.497398, 2.497391, 2.497386, 2.497377, 2.497379, 2.497376, 
    2.497373, 2.497369, 2.49737, 2.497368, 2.497376, 2.49737, 2.49738, 
    2.497377, 2.497397, 2.497405, 2.497408, 2.497411, 2.497418, 2.497414, 
    2.497416, 2.497411, 2.497408, 2.49741, 2.497401, 2.497404, 2.497386, 
    2.497394, 2.497374, 2.497379, 2.497373, 2.497375, 2.49737, 2.497375, 
    2.497367, 2.497365, 2.497366, 2.497362, 2.497375, 2.49737, 2.49741, 
    2.497409, 2.497408, 2.497413, 2.497413, 2.497418, 2.497414, 2.497412, 
    2.497408, 2.497405, 2.497403, 2.497398, 2.497392, 2.497384, 2.497378, 
    2.497374, 2.497377, 2.497375, 2.497377, 2.497378, 2.497366, 2.497373, 
    2.497362, 2.497363, 2.497368, 2.497363, 2.497409, 2.497411, 2.497415, 
    2.497411, 2.497418, 2.497414, 2.497412, 2.497404, 2.497402, 2.497401, 
    2.497397, 2.497393, 2.497386, 2.497379, 2.497373, 2.497374, 2.497374, 
    2.497372, 2.497375, 2.497372, 2.497371, 2.497373, 2.497363, 2.497366, 
    2.497363, 2.497365, 2.49741, 2.497408, 2.497409, 2.497407, 2.497408, 
    2.497401, 2.497399, 2.497389, 2.497393, 2.497386, 2.497392, 2.497391, 
    2.497386, 2.497392, 2.49738, 2.497388, 2.497372, 2.497381, 2.497372, 
    2.497373, 2.49737, 2.497368, 2.497365, 2.497359, 2.497361, 2.497356, 
    2.497404, 2.497401, 2.497402, 2.497399, 2.497396, 2.497391, 2.497384, 
    2.497387, 2.497381, 2.49738, 2.497388, 2.497383, 2.4974, 2.497397, 
    2.497398, 2.497404, 2.497386, 2.497395, 2.497378, 2.497383, 2.497368, 
    2.497376, 2.497361, 2.497355, 2.49735, 2.497343, 2.4974, 2.497402, 
    2.497398, 2.497393, 2.497389, 2.497383, 2.497382, 2.497381, 2.497378, 
    2.497376, 2.497381, 2.497375, 2.497396, 2.497385, 2.497403, 2.497397, 
    2.497394, 2.497395, 2.497387, 2.497385, 2.497377, 2.497381, 2.497357, 
    2.497368, 2.497338, 2.497346, 2.497403, 2.4974, 2.497391, 2.497395, 
    2.497382, 2.497379, 2.497377, 2.497374, 2.497373, 2.497371, 2.497375, 
    2.497371, 2.497383, 2.497378, 2.497392, 2.497388, 2.49739, 2.497391, 
    2.497386, 2.497381, 2.49738, 2.497379, 2.497374, 2.497382, 2.497355, 
    2.497372, 2.497397, 2.497392, 2.497391, 2.497393, 2.49738, 2.497385, 
    2.497371, 2.497375, 2.497369, 2.497372, 2.497372, 2.497376, 2.497378, 
    2.497384, 2.497389, 2.497393, 2.497392, 2.497388, 2.49738, 2.497373, 
    2.497375, 2.49737, 2.497383, 2.497378, 2.49738, 2.497374, 2.497387, 
    2.497376, 2.49739, 2.497388, 2.497385, 2.497377, 2.497375, 2.497374, 
    2.497375, 2.49738, 2.497381, 2.497385, 2.497386, 2.497389, 2.497391, 
    2.497389, 2.497386, 2.49738, 2.497374, 2.497368, 2.497366, 2.497359, 
    2.497365, 2.497355, 2.497364, 2.497349, 2.497375, 2.497364, 2.497385, 
    2.497382, 2.497378, 2.497369, 2.497374, 2.497368, 2.497381, 2.497388, 
    2.497389, 2.497393, 2.497389, 2.49739, 2.497386, 2.497387, 2.49738, 
    2.497384, 2.497372, 2.497368, 2.497356, 2.497349, 2.497342, 2.497339, 
    2.497338, 2.497337,
  2.497626, 2.497617, 2.497618, 2.497611, 2.497615, 2.497611, 2.497624, 
    2.497617, 2.497621, 2.497625, 2.497597, 2.497611, 2.497583, 2.497592, 
    2.497571, 2.497585, 2.497567, 2.497571, 2.497561, 2.497564, 2.497551, 
    2.49756, 2.497545, 2.497553, 2.497552, 2.49756, 2.497608, 2.497599, 
    2.497609, 2.497607, 2.497608, 2.497615, 2.497619, 2.497626, 2.497625, 
    2.497619, 2.497607, 2.497611, 2.497601, 2.497601, 2.497589, 2.497594, 
    2.497574, 2.49758, 2.497564, 2.497568, 2.497564, 2.497565, 2.497564, 
    2.49757, 2.497567, 2.497572, 2.497593, 2.497587, 2.497605, 2.497616, 
    2.497623, 2.497629, 2.497628, 2.497627, 2.497619, 2.497613, 2.497608, 
    2.497604, 2.497601, 2.497591, 2.497585, 2.497573, 2.497575, 2.497572, 
    2.497568, 2.497562, 2.497563, 2.497561, 2.497572, 2.497564, 2.497576, 
    2.497573, 2.4976, 2.49761, 2.497614, 2.497618, 2.497627, 2.497621, 
    2.497624, 2.497617, 2.497614, 2.497616, 2.497604, 2.497609, 2.497585, 
    2.497595, 2.497569, 2.497575, 2.497567, 2.497571, 2.497564, 2.49757, 
    2.49756, 2.497557, 2.497559, 2.497553, 2.497571, 2.497564, 2.497616, 
    2.497615, 2.497614, 2.49762, 2.497621, 2.497626, 2.497621, 2.497619, 
    2.497614, 2.49761, 2.497607, 2.4976, 2.497593, 2.497582, 2.497575, 
    2.497569, 2.497572, 2.49757, 2.497573, 2.497574, 2.497558, 2.497567, 
    2.497554, 2.497554, 2.497561, 2.497554, 2.497615, 2.497617, 2.497623, 
    2.497618, 2.497627, 2.497622, 2.497619, 2.497608, 2.497606, 2.497604, 
    2.4976, 2.497594, 2.497584, 2.497576, 2.497568, 2.497569, 2.497568, 
    2.497566, 2.497571, 2.497566, 2.497565, 2.497567, 2.497555, 2.497558, 
    2.497554, 2.497557, 2.497616, 2.497613, 2.497615, 2.497612, 2.497614, 
    2.497605, 2.497602, 2.497589, 2.497594, 2.497586, 2.497593, 2.497592, 
    2.497585, 2.497593, 2.497576, 2.497587, 2.497566, 2.497578, 2.497566, 
    2.497568, 2.497564, 2.497561, 2.497557, 2.49755, 2.497551, 2.497545, 
    2.497609, 2.497605, 2.497606, 2.497602, 2.497598, 2.497592, 2.497582, 
    2.497586, 2.497579, 2.497577, 2.497588, 2.497581, 2.497603, 2.497599, 
    2.497601, 2.497609, 2.497585, 2.497597, 2.497574, 2.497581, 2.497562, 
    2.497571, 2.497552, 2.497544, 2.497537, 2.497528, 2.497603, 2.497606, 
    2.497601, 2.497595, 2.497589, 2.497581, 2.49758, 2.497578, 2.497574, 
    2.497571, 2.497578, 2.49757, 2.497598, 2.497584, 2.497607, 2.4976, 
    2.497595, 2.497597, 2.497586, 2.497583, 2.497573, 2.497578, 2.497546, 
    2.497561, 2.497521, 2.497532, 2.497607, 2.497603, 2.497591, 2.497597, 
    2.49758, 2.497576, 2.497573, 2.497568, 2.497568, 2.497566, 2.49757, 
    2.497566, 2.497581, 2.497574, 2.497592, 2.497588, 2.49759, 2.497592, 
    2.497585, 2.497578, 2.497578, 2.497575, 2.497568, 2.49758, 2.497545, 
    2.497566, 2.497599, 2.497592, 2.497591, 2.497594, 2.497576, 2.497583, 
    2.497566, 2.49757, 2.497562, 2.497566, 2.497567, 2.497572, 2.497575, 
    2.497582, 2.497589, 2.497594, 2.497593, 2.497587, 2.497577, 2.497568, 
    2.49757, 2.497563, 2.497581, 2.497574, 2.497576, 2.497569, 2.497586, 
    2.497571, 2.497589, 2.497588, 2.497583, 2.497573, 2.497571, 2.497569, 
    2.49757, 2.497577, 2.497578, 2.497583, 2.497584, 2.497588, 2.497591, 
    2.497588, 2.497586, 2.497577, 2.497569, 2.497561, 2.497559, 2.497549, 
    2.497557, 2.497544, 2.497555, 2.497536, 2.497571, 2.497556, 2.497583, 
    2.49758, 2.497575, 2.497562, 2.497569, 2.497561, 2.497578, 2.497587, 
    2.497589, 2.497593, 2.497589, 2.49759, 2.497585, 2.497587, 2.497577, 
    2.497582, 2.497567, 2.497561, 2.497546, 2.497536, 2.497527, 2.497522, 
    2.497521, 2.49752,
  2.497841, 2.497832, 2.497833, 2.497826, 2.49783, 2.497825, 2.497839, 
    2.497831, 2.497836, 2.49784, 2.497811, 2.497825, 2.497796, 2.497805, 
    2.497782, 2.497797, 2.497779, 2.497782, 2.497772, 2.497775, 2.497761, 
    2.49777, 2.497754, 2.497763, 2.497762, 2.497771, 2.497823, 2.497813, 
    2.497823, 2.497822, 2.497822, 2.49783, 2.497834, 2.497842, 2.49784, 
    2.497834, 2.497821, 2.497826, 2.497814, 2.497814, 2.497802, 2.497808, 
    2.497786, 2.497792, 2.497775, 2.497779, 2.497775, 2.497776, 2.497775, 
    2.497781, 2.497779, 2.497784, 2.497806, 2.4978, 2.497819, 2.497831, 
    2.497839, 2.497844, 2.497844, 2.497842, 2.497834, 2.497827, 2.497822, 
    2.497818, 2.497814, 2.497803, 2.497798, 2.497785, 2.497787, 2.497783, 
    2.49778, 2.497773, 2.497774, 2.497772, 2.497783, 2.497776, 2.497789, 
    2.497785, 2.497813, 2.497824, 2.497829, 2.497833, 2.497843, 2.497836, 
    2.497839, 2.497832, 2.497828, 2.49783, 2.497818, 2.497823, 2.497797, 
    2.497808, 2.49778, 2.497787, 2.497778, 2.497783, 2.497775, 2.497782, 
    2.497771, 2.497768, 2.49777, 2.497763, 2.497782, 2.497775, 2.49783, 
    2.49783, 2.497828, 2.497835, 2.497836, 2.497842, 2.497836, 2.497834, 
    2.497828, 2.497825, 2.497821, 2.497814, 2.497806, 2.497794, 2.497786, 
    2.497781, 2.497784, 2.497781, 2.497785, 2.497786, 2.497769, 2.497779, 
    2.497764, 2.497765, 2.497772, 2.497765, 2.49783, 2.497832, 2.497838, 
    2.497833, 2.497843, 2.497837, 2.497834, 2.497823, 2.49782, 2.497818, 
    2.497813, 2.497807, 2.497797, 2.497788, 2.497779, 2.49778, 2.49778, 
    2.497778, 2.497782, 2.497777, 2.497776, 2.497779, 2.497765, 2.497769, 
    2.497765, 2.497767, 2.497831, 2.497828, 2.49783, 2.497826, 2.497829, 
    2.497819, 2.497816, 2.497802, 2.497807, 2.497798, 2.497806, 2.497805, 
    2.497798, 2.497806, 2.497788, 2.4978, 2.497778, 2.49779, 2.497777, 
    2.497779, 2.497776, 2.497772, 2.497768, 2.49776, 2.497762, 2.497755, 
    2.497823, 2.497819, 2.497819, 2.497815, 2.497812, 2.497805, 2.497794, 
    2.497798, 2.497791, 2.497789, 2.497801, 2.497794, 2.497816, 2.497813, 
    2.497815, 2.497823, 2.497797, 2.49781, 2.497786, 2.497793, 2.497773, 
    2.497783, 2.497763, 2.497754, 2.497746, 2.497736, 2.497817, 2.49782, 
    2.497815, 2.497808, 2.497801, 2.497793, 2.497792, 2.49779, 2.497786, 
    2.497783, 2.49779, 2.497782, 2.497812, 2.497796, 2.497821, 2.497813, 
    2.497808, 2.49781, 2.497799, 2.497796, 2.497785, 2.497791, 2.497756, 
    2.497771, 2.497729, 2.497741, 2.497821, 2.497817, 2.497804, 2.49781, 
    2.497792, 2.497788, 2.497784, 2.49778, 2.497779, 2.497777, 2.497781, 
    2.497777, 2.497793, 2.497786, 2.497805, 2.497801, 2.497803, 2.497805, 
    2.497798, 2.49779, 2.49779, 2.497787, 2.49778, 2.497792, 2.497754, 
    2.497778, 2.497813, 2.497806, 2.497805, 2.497807, 2.497788, 2.497795, 
    2.497777, 2.497782, 2.497774, 2.497778, 2.497778, 2.497783, 2.497787, 
    2.497795, 2.497802, 2.497807, 2.497806, 2.4978, 2.497789, 2.497779, 
    2.497782, 2.497774, 2.497794, 2.497785, 2.497789, 2.49778, 2.497798, 
    2.497783, 2.497802, 2.497801, 2.497795, 2.497785, 2.497782, 2.49778, 
    2.497782, 2.497789, 2.49779, 2.497796, 2.497797, 2.497801, 2.497804, 
    2.497801, 2.497798, 2.497789, 2.497781, 2.497772, 2.49777, 2.49776, 
    2.497768, 2.497754, 2.497766, 2.497746, 2.497782, 2.497766, 2.497795, 
    2.497792, 2.497786, 2.497773, 2.49778, 2.497772, 2.49779, 2.4978, 
    2.497802, 2.497807, 2.497802, 2.497802, 2.497798, 2.497799, 2.497789, 
    2.497794, 2.497778, 2.497772, 2.497756, 2.497746, 2.497735, 2.49773, 
    2.497729, 2.497729,
  2.498013, 2.498003, 2.498005, 2.497998, 2.498002, 2.497997, 2.498011, 
    2.498003, 2.498008, 2.498012, 2.497983, 2.497997, 2.497968, 2.497977, 
    2.497954, 2.49797, 2.497951, 2.497955, 2.497944, 2.497947, 2.497934, 
    2.497943, 2.497927, 2.497936, 2.497934, 2.497943, 2.497994, 2.497985, 
    2.497995, 2.497994, 2.497994, 2.498002, 2.498006, 2.498013, 2.498012, 
    2.498006, 2.497993, 2.497998, 2.497986, 2.497987, 2.497974, 2.49798, 
    2.497958, 2.497964, 2.497947, 2.497952, 2.497947, 2.497948, 2.497947, 
    2.497954, 2.497951, 2.497957, 2.497978, 2.497972, 2.497991, 2.498003, 
    2.498011, 2.498016, 2.498015, 2.498014, 2.498006, 2.497999, 2.497994, 
    2.49799, 2.497987, 2.497976, 2.49797, 2.497957, 2.49796, 2.497956, 
    2.497952, 2.497946, 2.497947, 2.497944, 2.497956, 2.497948, 2.497961, 
    2.497957, 2.497986, 2.497996, 2.498001, 2.498005, 2.498015, 2.498008, 
    2.498011, 2.498004, 2.498, 2.498002, 2.49799, 2.497995, 2.49797, 2.49798, 
    2.497952, 2.497959, 2.497951, 2.497955, 2.497948, 2.497954, 2.497943, 
    2.49794, 2.497942, 2.497936, 2.497955, 2.497947, 2.498002, 2.498002, 
    2.498, 2.498007, 2.498008, 2.498013, 2.498008, 2.498006, 2.498, 2.497997, 
    2.497993, 2.497986, 2.497978, 2.497967, 2.497959, 2.497953, 2.497957, 
    2.497954, 2.497957, 2.497958, 2.497941, 2.497951, 2.497936, 2.497937, 
    2.497944, 2.497937, 2.498002, 2.498003, 2.49801, 2.498005, 2.498014, 
    2.498009, 2.498006, 2.497995, 2.497992, 2.49799, 2.497985, 2.497979, 
    2.497969, 2.49796, 2.497952, 2.497952, 2.497952, 2.49795, 2.497955, 
    2.497949, 2.497949, 2.497951, 2.497937, 2.497941, 2.497937, 2.49794, 
    2.498003, 2.498, 2.498002, 2.497998, 2.498001, 2.497991, 2.497988, 
    2.497974, 2.497979, 2.49797, 2.497978, 2.497977, 2.49797, 2.497978, 
    2.49796, 2.497972, 2.49795, 2.497962, 2.497949, 2.497952, 2.497948, 
    2.497944, 2.49794, 2.497932, 2.497934, 2.497927, 2.497995, 2.497991, 
    2.497992, 2.497987, 2.497984, 2.497977, 2.497966, 2.49797, 2.497963, 
    2.497961, 2.497973, 2.497966, 2.497988, 2.497985, 2.497987, 2.497995, 
    2.497969, 2.497983, 2.497958, 2.497966, 2.497945, 2.497955, 2.497935, 
    2.497926, 2.497918, 2.497909, 2.497989, 2.497992, 2.497987, 2.49798, 
    2.497973, 2.497965, 2.497964, 2.497963, 2.497959, 2.497955, 2.497962, 
    2.497954, 2.497984, 2.497968, 2.497993, 2.497985, 2.49798, 2.497983, 
    2.497971, 2.497968, 2.497957, 2.497963, 2.497929, 2.497944, 2.497902, 
    2.497914, 2.497993, 2.497989, 2.497976, 2.497982, 2.497965, 2.49796, 
    2.497957, 2.497952, 2.497952, 2.497949, 2.497953, 2.497949, 2.497965, 
    2.497958, 2.497977, 2.497973, 2.497975, 2.497977, 2.49797, 2.497962, 
    2.497962, 2.497959, 2.497952, 2.497964, 2.497927, 2.49795, 2.497985, 
    2.497978, 2.497977, 2.497979, 2.497961, 2.497967, 2.497949, 2.497954, 
    2.497946, 2.49795, 2.497951, 2.497956, 2.497959, 2.497967, 2.497974, 
    2.497979, 2.497978, 2.497972, 2.497962, 2.497952, 2.497954, 2.497947, 
    2.497966, 2.497958, 2.497961, 2.497953, 2.497971, 2.497955, 2.497974, 
    2.497973, 2.497967, 2.497957, 2.497955, 2.497952, 2.497954, 2.497961, 
    2.497962, 2.497968, 2.497969, 2.497973, 2.497976, 2.497973, 2.49797, 
    2.497961, 2.497953, 2.497944, 2.497942, 2.497932, 2.49794, 2.497926, 
    2.497938, 2.497918, 2.497954, 2.497939, 2.497967, 2.497964, 2.497959, 
    2.497946, 2.497953, 2.497945, 2.497962, 2.497972, 2.497974, 2.497979, 
    2.497974, 2.497974, 2.49797, 2.497972, 2.497961, 2.497967, 2.497951, 
    2.497945, 2.497928, 2.497918, 2.497908, 2.497903, 2.497902, 2.497901,
  2.498213, 2.498205, 2.498207, 2.4982, 2.498204, 2.498199, 2.498212, 
    2.498205, 2.498209, 2.498213, 2.498187, 2.498199, 2.498174, 2.498182, 
    2.498161, 2.498175, 2.498159, 2.498162, 2.498152, 2.498155, 2.498143, 
    2.498151, 2.498137, 2.498145, 2.498144, 2.498151, 2.498197, 2.498188, 
    2.498198, 2.498196, 2.498197, 2.498204, 2.498207, 2.498214, 2.498213, 
    2.498207, 2.498196, 2.4982, 2.49819, 2.49819, 2.498179, 2.498184, 
    2.498165, 2.49817, 2.498155, 2.498159, 2.498155, 2.498156, 2.498155, 
    2.498161, 2.498158, 2.498163, 2.498183, 2.498177, 2.498194, 2.498204, 
    2.498211, 2.498216, 2.498215, 2.498214, 2.498207, 2.498201, 2.498196, 
    2.498193, 2.49819, 2.49818, 2.498175, 2.498164, 2.498166, 2.498163, 
    2.498159, 2.498154, 2.498154, 2.498152, 2.498163, 2.498156, 2.498167, 
    2.498164, 2.498189, 2.498199, 2.498203, 2.498206, 2.498215, 2.498209, 
    2.498211, 2.498206, 2.498202, 2.498204, 2.498193, 2.498197, 2.498175, 
    2.498185, 2.49816, 2.498166, 2.498158, 2.498162, 2.498155, 2.498161, 
    2.498151, 2.498149, 2.49815, 2.498145, 2.498162, 2.498155, 2.498204, 
    2.498204, 2.498202, 2.498208, 2.498209, 2.498214, 2.498209, 2.498207, 
    2.498202, 2.498199, 2.498196, 2.498189, 2.498182, 2.498172, 2.498165, 
    2.49816, 2.498163, 2.498161, 2.498164, 2.498165, 2.49815, 2.498158, 
    2.498145, 2.498146, 2.498152, 2.498146, 2.498204, 2.498205, 2.498211, 
    2.498206, 2.498214, 2.49821, 2.498207, 2.498197, 2.498195, 2.498193, 
    2.498189, 2.498183, 2.498174, 2.498166, 2.498159, 2.498159, 2.498159, 
    2.498158, 2.498162, 2.498157, 2.498156, 2.498158, 2.498146, 2.49815, 
    2.498146, 2.498148, 2.498204, 2.498202, 2.498203, 2.4982, 2.498202, 
    2.498194, 2.498191, 2.498178, 2.498184, 2.498175, 2.498183, 2.498182, 
    2.498175, 2.498182, 2.498167, 2.498177, 2.498158, 2.498168, 2.498157, 
    2.498159, 2.498156, 2.498152, 2.498149, 2.498142, 2.498143, 2.498137, 
    2.498198, 2.498194, 2.498194, 2.498191, 2.498188, 2.498182, 2.498172, 
    2.498176, 2.498169, 2.498168, 2.498178, 2.498172, 2.498192, 2.498188, 
    2.49819, 2.498197, 2.498175, 2.498186, 2.498165, 2.498171, 2.498153, 
    2.498162, 2.498144, 2.498137, 2.498129, 2.498121, 2.498192, 2.498194, 
    2.49819, 2.498184, 2.498178, 2.498171, 2.49817, 2.498169, 2.498165, 
    2.498162, 2.498168, 2.498161, 2.498188, 2.498174, 2.498195, 2.498189, 
    2.498184, 2.498186, 2.498176, 2.498174, 2.498164, 2.498169, 2.498138, 
    2.498152, 2.498115, 2.498125, 2.498195, 2.498192, 2.498181, 2.498186, 
    2.49817, 2.498167, 2.498163, 2.498159, 2.498159, 2.498157, 2.498161, 
    2.498157, 2.498171, 2.498165, 2.498182, 2.498178, 2.49818, 2.498182, 
    2.498175, 2.498168, 2.498168, 2.498166, 2.498159, 2.49817, 2.498137, 
    2.498158, 2.498188, 2.498182, 2.498181, 2.498184, 2.498167, 2.498173, 
    2.498157, 2.498161, 2.498154, 2.498158, 2.498158, 2.498163, 2.498165, 
    2.498173, 2.498179, 2.498183, 2.498182, 2.498177, 2.498168, 2.498159, 
    2.498161, 2.498154, 2.498172, 2.498164, 2.498167, 2.49816, 2.498176, 
    2.498162, 2.498179, 2.498178, 2.498173, 2.498164, 2.498162, 2.49816, 
    2.498161, 2.498168, 2.498169, 2.498173, 2.498174, 2.498178, 2.498181, 
    2.498178, 2.498175, 2.498168, 2.49816, 2.498152, 2.498151, 2.498142, 
    2.498149, 2.498137, 2.498147, 2.498129, 2.498162, 2.498147, 2.498173, 
    2.49817, 2.498165, 2.498154, 2.49816, 2.498153, 2.498169, 2.498177, 
    2.498179, 2.498183, 2.498179, 2.498179, 2.498175, 2.498177, 2.498167, 
    2.498172, 2.498158, 2.498153, 2.498138, 2.498129, 2.49812, 2.498116, 
    2.498114, 2.498114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.139198e-08, 6.166193e-08, 6.160945e-08, 6.182718e-08, 6.170639e-08, 
    6.184897e-08, 6.144671e-08, 6.167265e-08, 6.152841e-08, 6.141628e-08, 
    6.224973e-08, 6.183689e-08, 6.267852e-08, 6.241524e-08, 6.307661e-08, 
    6.263755e-08, 6.316512e-08, 6.306393e-08, 6.33685e-08, 6.328124e-08, 
    6.367082e-08, 6.340877e-08, 6.387275e-08, 6.360823e-08, 6.364962e-08, 
    6.340012e-08, 6.191997e-08, 6.219834e-08, 6.190348e-08, 6.194317e-08, 
    6.192536e-08, 6.17089e-08, 6.159981e-08, 6.137134e-08, 6.141282e-08, 
    6.158062e-08, 6.196102e-08, 6.183189e-08, 6.215732e-08, 6.214997e-08, 
    6.251226e-08, 6.234892e-08, 6.295784e-08, 6.278477e-08, 6.328489e-08, 
    6.315911e-08, 6.327897e-08, 6.324263e-08, 6.327945e-08, 6.309499e-08, 
    6.317403e-08, 6.301171e-08, 6.237951e-08, 6.256531e-08, 6.201116e-08, 
    6.167795e-08, 6.145662e-08, 6.129956e-08, 6.132176e-08, 6.136409e-08, 
    6.15816e-08, 6.17861e-08, 6.194195e-08, 6.20462e-08, 6.214891e-08, 
    6.245984e-08, 6.262439e-08, 6.299284e-08, 6.292634e-08, 6.303899e-08, 
    6.31466e-08, 6.332728e-08, 6.329753e-08, 6.337714e-08, 6.303601e-08, 
    6.326273e-08, 6.288847e-08, 6.299083e-08, 6.217687e-08, 6.186672e-08, 
    6.173492e-08, 6.161954e-08, 6.133883e-08, 6.153268e-08, 6.145627e-08, 
    6.163806e-08, 6.175357e-08, 6.169644e-08, 6.204905e-08, 6.191197e-08, 
    6.263414e-08, 6.232308e-08, 6.313405e-08, 6.293999e-08, 6.318056e-08, 
    6.30578e-08, 6.326815e-08, 6.307884e-08, 6.340677e-08, 6.347817e-08, 
    6.342938e-08, 6.361681e-08, 6.306834e-08, 6.327898e-08, 6.169484e-08, 
    6.170416e-08, 6.174757e-08, 6.155675e-08, 6.154508e-08, 6.137021e-08, 
    6.152581e-08, 6.159207e-08, 6.176027e-08, 6.185977e-08, 6.195435e-08, 
    6.216229e-08, 6.239453e-08, 6.271927e-08, 6.295257e-08, 6.310896e-08, 
    6.301306e-08, 6.309772e-08, 6.300308e-08, 6.295872e-08, 6.345142e-08, 
    6.317477e-08, 6.358985e-08, 6.356689e-08, 6.337903e-08, 6.356947e-08, 
    6.171071e-08, 6.165708e-08, 6.147091e-08, 6.161661e-08, 6.135116e-08, 
    6.149975e-08, 6.158519e-08, 6.191484e-08, 6.198726e-08, 6.205442e-08, 
    6.218706e-08, 6.235727e-08, 6.265589e-08, 6.291569e-08, 6.315286e-08, 
    6.313548e-08, 6.31416e-08, 6.319458e-08, 6.306334e-08, 6.321613e-08, 
    6.324178e-08, 6.317472e-08, 6.356381e-08, 6.345265e-08, 6.35664e-08, 
    6.349402e-08, 6.167451e-08, 6.176474e-08, 6.171599e-08, 6.180766e-08, 
    6.174308e-08, 6.203027e-08, 6.211638e-08, 6.251928e-08, 6.235393e-08, 
    6.261709e-08, 6.238066e-08, 6.242255e-08, 6.262568e-08, 6.239343e-08, 
    6.290137e-08, 6.255701e-08, 6.319664e-08, 6.285278e-08, 6.32182e-08, 
    6.315184e-08, 6.32617e-08, 6.33601e-08, 6.348389e-08, 6.371231e-08, 
    6.365941e-08, 6.385043e-08, 6.189924e-08, 6.201627e-08, 6.200596e-08, 
    6.212843e-08, 6.2219e-08, 6.24153e-08, 6.273014e-08, 6.261175e-08, 
    6.28291e-08, 6.287274e-08, 6.254253e-08, 6.274527e-08, 6.209459e-08, 
    6.219972e-08, 6.213713e-08, 6.190847e-08, 6.263904e-08, 6.226412e-08, 
    6.295642e-08, 6.275332e-08, 6.334607e-08, 6.30513e-08, 6.36303e-08, 
    6.387783e-08, 6.411076e-08, 6.438301e-08, 6.208013e-08, 6.200062e-08, 
    6.214299e-08, 6.233998e-08, 6.252274e-08, 6.276571e-08, 6.279057e-08, 
    6.283609e-08, 6.295399e-08, 6.305312e-08, 6.285049e-08, 6.307798e-08, 
    6.222412e-08, 6.267158e-08, 6.197056e-08, 6.218166e-08, 6.232837e-08, 
    6.226401e-08, 6.259822e-08, 6.267699e-08, 6.299708e-08, 6.283161e-08, 
    6.381674e-08, 6.33809e-08, 6.459028e-08, 6.425232e-08, 6.197283e-08, 
    6.207986e-08, 6.245234e-08, 6.227511e-08, 6.278193e-08, 6.290668e-08, 
    6.300809e-08, 6.313773e-08, 6.315172e-08, 6.322854e-08, 6.310267e-08, 
    6.322357e-08, 6.276623e-08, 6.29706e-08, 6.240975e-08, 6.254626e-08, 
    6.248347e-08, 6.241458e-08, 6.262718e-08, 6.285368e-08, 6.285851e-08, 
    6.293114e-08, 6.313581e-08, 6.278398e-08, 6.387301e-08, 6.320047e-08, 
    6.219656e-08, 6.240271e-08, 6.243214e-08, 6.235229e-08, 6.289417e-08, 
    6.269784e-08, 6.322666e-08, 6.308374e-08, 6.331792e-08, 6.320155e-08, 
    6.318443e-08, 6.303497e-08, 6.294192e-08, 6.270684e-08, 6.251556e-08, 
    6.236387e-08, 6.239914e-08, 6.256577e-08, 6.286754e-08, 6.3153e-08, 
    6.309047e-08, 6.330012e-08, 6.274518e-08, 6.297788e-08, 6.288795e-08, 
    6.312245e-08, 6.260861e-08, 6.30462e-08, 6.249675e-08, 6.254493e-08, 
    6.269394e-08, 6.299367e-08, 6.305997e-08, 6.313078e-08, 6.308709e-08, 
    6.287519e-08, 6.284047e-08, 6.269031e-08, 6.264886e-08, 6.253444e-08, 
    6.243971e-08, 6.252626e-08, 6.261715e-08, 6.287528e-08, 6.310789e-08, 
    6.33615e-08, 6.342356e-08, 6.37199e-08, 6.347868e-08, 6.387675e-08, 
    6.353834e-08, 6.412414e-08, 6.307155e-08, 6.352837e-08, 6.270071e-08, 
    6.278988e-08, 6.295116e-08, 6.332105e-08, 6.312135e-08, 6.335489e-08, 
    6.283911e-08, 6.257152e-08, 6.250227e-08, 6.23731e-08, 6.250522e-08, 
    6.249448e-08, 6.262091e-08, 6.258028e-08, 6.288385e-08, 6.272079e-08, 
    6.3184e-08, 6.335304e-08, 6.383041e-08, 6.412306e-08, 6.442093e-08, 
    6.455244e-08, 6.459247e-08, 6.46092e-08 ;

 SOIL1_HR_S3 =
  7.285347e-10, 7.317394e-10, 7.311164e-10, 7.337012e-10, 7.322673e-10, 
    7.339599e-10, 7.291844e-10, 7.318667e-10, 7.301543e-10, 7.288232e-10, 
    7.387176e-10, 7.338165e-10, 7.438081e-10, 7.406825e-10, 7.485342e-10, 
    7.433218e-10, 7.495852e-10, 7.483837e-10, 7.519997e-10, 7.509637e-10, 
    7.55589e-10, 7.524777e-10, 7.579865e-10, 7.548459e-10, 7.553372e-10, 
    7.523752e-10, 7.348028e-10, 7.381075e-10, 7.34607e-10, 7.350782e-10, 
    7.348667e-10, 7.32297e-10, 7.31002e-10, 7.282897e-10, 7.287821e-10, 
    7.307742e-10, 7.352901e-10, 7.337571e-10, 7.376205e-10, 7.375333e-10, 
    7.418344e-10, 7.398951e-10, 7.471243e-10, 7.450696e-10, 7.51007e-10, 
    7.495138e-10, 7.509369e-10, 7.505053e-10, 7.509425e-10, 7.487526e-10, 
    7.496908e-10, 7.477638e-10, 7.402583e-10, 7.424641e-10, 7.358853e-10, 
    7.319297e-10, 7.293021e-10, 7.274376e-10, 7.277012e-10, 7.282037e-10, 
    7.307859e-10, 7.332136e-10, 7.350637e-10, 7.363013e-10, 7.375207e-10, 
    7.41212e-10, 7.431655e-10, 7.475398e-10, 7.467503e-10, 7.480877e-10, 
    7.493652e-10, 7.515103e-10, 7.511572e-10, 7.521023e-10, 7.480523e-10, 
    7.50744e-10, 7.463006e-10, 7.475159e-10, 7.378526e-10, 7.341707e-10, 
    7.32606e-10, 7.312362e-10, 7.279038e-10, 7.302051e-10, 7.292979e-10, 
    7.314561e-10, 7.328274e-10, 7.321492e-10, 7.363352e-10, 7.347077e-10, 
    7.432813e-10, 7.395884e-10, 7.492162e-10, 7.469123e-10, 7.497685e-10, 
    7.48311e-10, 7.508082e-10, 7.485608e-10, 7.52454e-10, 7.533018e-10, 
    7.527224e-10, 7.549478e-10, 7.484361e-10, 7.509369e-10, 7.321302e-10, 
    7.322408e-10, 7.327561e-10, 7.304908e-10, 7.303523e-10, 7.282763e-10, 
    7.301235e-10, 7.309101e-10, 7.329069e-10, 7.340881e-10, 7.352108e-10, 
    7.376795e-10, 7.404367e-10, 7.44292e-10, 7.470616e-10, 7.489183e-10, 
    7.477798e-10, 7.487849e-10, 7.476613e-10, 7.471347e-10, 7.529841e-10, 
    7.496996e-10, 7.546277e-10, 7.54355e-10, 7.521248e-10, 7.543857e-10, 
    7.323185e-10, 7.316819e-10, 7.294718e-10, 7.312014e-10, 7.280502e-10, 
    7.298141e-10, 7.308284e-10, 7.347418e-10, 7.356016e-10, 7.363989e-10, 
    7.379735e-10, 7.399943e-10, 7.435394e-10, 7.466238e-10, 7.494396e-10, 
    7.492332e-10, 7.493059e-10, 7.499349e-10, 7.483768e-10, 7.501907e-10, 
    7.504952e-10, 7.496992e-10, 7.543184e-10, 7.529988e-10, 7.543492e-10, 
    7.534899e-10, 7.318888e-10, 7.329599e-10, 7.323812e-10, 7.334695e-10, 
    7.327028e-10, 7.361123e-10, 7.371345e-10, 7.419177e-10, 7.399546e-10, 
    7.430788e-10, 7.402719e-10, 7.407693e-10, 7.431809e-10, 7.404236e-10, 
    7.464538e-10, 7.423656e-10, 7.499594e-10, 7.45877e-10, 7.502152e-10, 
    7.494274e-10, 7.507318e-10, 7.519e-10, 7.533696e-10, 7.560815e-10, 
    7.554535e-10, 7.577213e-10, 7.345567e-10, 7.35946e-10, 7.358236e-10, 
    7.372775e-10, 7.383528e-10, 7.406832e-10, 7.44421e-10, 7.430154e-10, 
    7.455959e-10, 7.461139e-10, 7.421936e-10, 7.446007e-10, 7.368758e-10, 
    7.381239e-10, 7.373807e-10, 7.346663e-10, 7.433394e-10, 7.388884e-10, 
    7.471074e-10, 7.446962e-10, 7.517335e-10, 7.482337e-10, 7.551078e-10, 
    7.580467e-10, 7.608122e-10, 7.640446e-10, 7.367042e-10, 7.357602e-10, 
    7.374504e-10, 7.39789e-10, 7.419587e-10, 7.448433e-10, 7.451384e-10, 
    7.456788e-10, 7.470786e-10, 7.482555e-10, 7.458498e-10, 7.485505e-10, 
    7.384135e-10, 7.437257e-10, 7.354033e-10, 7.379095e-10, 7.396511e-10, 
    7.388871e-10, 7.428548e-10, 7.4379e-10, 7.475902e-10, 7.456256e-10, 
    7.573214e-10, 7.521468e-10, 7.665055e-10, 7.624929e-10, 7.354304e-10, 
    7.367009e-10, 7.411229e-10, 7.390189e-10, 7.450358e-10, 7.465168e-10, 
    7.477208e-10, 7.4926e-10, 7.494261e-10, 7.50338e-10, 7.488437e-10, 
    7.50279e-10, 7.448494e-10, 7.472757e-10, 7.406174e-10, 7.42238e-10, 
    7.414924e-10, 7.406747e-10, 7.431986e-10, 7.458876e-10, 7.45945e-10, 
    7.468072e-10, 7.492372e-10, 7.450602e-10, 7.579894e-10, 7.500048e-10, 
    7.380864e-10, 7.405337e-10, 7.408832e-10, 7.399352e-10, 7.463684e-10, 
    7.440374e-10, 7.503158e-10, 7.486189e-10, 7.513992e-10, 7.500176e-10, 
    7.498144e-10, 7.4804e-10, 7.469353e-10, 7.441444e-10, 7.418735e-10, 
    7.400727e-10, 7.404914e-10, 7.424695e-10, 7.460521e-10, 7.494412e-10, 
    7.486988e-10, 7.511879e-10, 7.445995e-10, 7.473622e-10, 7.462945e-10, 
    7.490785e-10, 7.429781e-10, 7.481733e-10, 7.416502e-10, 7.422221e-10, 
    7.439911e-10, 7.475496e-10, 7.483368e-10, 7.491774e-10, 7.486587e-10, 
    7.46143e-10, 7.457309e-10, 7.439481e-10, 7.43456e-10, 7.420976e-10, 
    7.409731e-10, 7.420005e-10, 7.430796e-10, 7.46144e-10, 7.489057e-10, 
    7.519166e-10, 7.526534e-10, 7.561717e-10, 7.533078e-10, 7.58034e-10, 
    7.540161e-10, 7.609711e-10, 7.484742e-10, 7.538977e-10, 7.440716e-10, 
    7.451302e-10, 7.470449e-10, 7.514363e-10, 7.490654e-10, 7.518381e-10, 
    7.457147e-10, 7.425378e-10, 7.417157e-10, 7.401821e-10, 7.417508e-10, 
    7.416232e-10, 7.431242e-10, 7.426419e-10, 7.462458e-10, 7.443099e-10, 
    7.498093e-10, 7.518162e-10, 7.574837e-10, 7.609582e-10, 7.644948e-10, 
    7.660562e-10, 7.665314e-10, 7.667301e-10 ;

 SOIL2C =
  5.784045, 5.784051, 5.78405, 5.784055, 5.784052, 5.784055, 5.784046, 
    5.784051, 5.784048, 5.784045, 5.784065, 5.784055, 5.784075, 5.784069, 
    5.784084, 5.784074, 5.784086, 5.784084, 5.784091, 5.784089, 5.784098, 
    5.784092, 5.784103, 5.784097, 5.784098, 5.784091, 5.784057, 5.784063, 
    5.784057, 5.784058, 5.784057, 5.784052, 5.78405, 5.784044, 5.784045, 
    5.784049, 5.784058, 5.784055, 5.784062, 5.784062, 5.784071, 5.784067, 
    5.784081, 5.784077, 5.784089, 5.784086, 5.784089, 5.784088, 5.784089, 
    5.784084, 5.784086, 5.784082, 5.784068, 5.784072, 5.784059, 5.784051, 
    5.784046, 5.784042, 5.784043, 5.784044, 5.784049, 5.784054, 5.784058, 
    5.78406, 5.784062, 5.78407, 5.784073, 5.784082, 5.784081, 5.784083, 
    5.784086, 5.78409, 5.784089, 5.784091, 5.784083, 5.784089, 5.78408, 
    5.784082, 5.784063, 5.784056, 5.784052, 5.78405, 5.784043, 5.784048, 
    5.784046, 5.78405, 5.784053, 5.784052, 5.78406, 5.784057, 5.784074, 
    5.784066, 5.784085, 5.784081, 5.784087, 5.784084, 5.784089, 5.784084, 
    5.784092, 5.784093, 5.784092, 5.784097, 5.784084, 5.784089, 5.784051, 
    5.784052, 5.784053, 5.784049, 5.784048, 5.784044, 5.784048, 5.784049, 
    5.784053, 5.784056, 5.784058, 5.784062, 5.784068, 5.784076, 5.784081, 
    5.784085, 5.784082, 5.784084, 5.784082, 5.784081, 5.784093, 5.784086, 
    5.784096, 5.784096, 5.784091, 5.784096, 5.784052, 5.784051, 5.784046, 
    5.78405, 5.784044, 5.784047, 5.784049, 5.784057, 5.784059, 5.78406, 
    5.784063, 5.784067, 5.784074, 5.784081, 5.784086, 5.784085, 5.784086, 
    5.784087, 5.784084, 5.784087, 5.784088, 5.784086, 5.784095, 5.784093, 
    5.784096, 5.784094, 5.784051, 5.784053, 5.784052, 5.784054, 5.784053, 
    5.78406, 5.784061, 5.784071, 5.784067, 5.784073, 5.784068, 5.784069, 
    5.784073, 5.784068, 5.78408, 5.784072, 5.784087, 5.784079, 5.784087, 
    5.784086, 5.784089, 5.784091, 5.784093, 5.784099, 5.784098, 5.784102, 
    5.784057, 5.784059, 5.784059, 5.784062, 5.784064, 5.784069, 5.784076, 
    5.784073, 5.784078, 5.784079, 5.784071, 5.784076, 5.784061, 5.784063, 
    5.784062, 5.784057, 5.784074, 5.784065, 5.784081, 5.784077, 5.784091, 
    5.784083, 5.784097, 5.784103, 5.784108, 5.784115, 5.78406, 5.784059, 
    5.784062, 5.784067, 5.784071, 5.784077, 5.784077, 5.784079, 5.784081, 
    5.784083, 5.784079, 5.784084, 5.784064, 5.784075, 5.784058, 5.784063, 
    5.784067, 5.784065, 5.784073, 5.784075, 5.784082, 5.784078, 5.784101, 
    5.784091, 5.78412, 5.784111, 5.784058, 5.78406, 5.78407, 5.784065, 
    5.784077, 5.78408, 5.784082, 5.784085, 5.784086, 5.784088, 5.784085, 
    5.784088, 5.784077, 5.784081, 5.784069, 5.784071, 5.78407, 5.784069, 
    5.784073, 5.784079, 5.784079, 5.784081, 5.784085, 5.784077, 5.784103, 
    5.784087, 5.784063, 5.784068, 5.784069, 5.784067, 5.78408, 5.784075, 
    5.784088, 5.784084, 5.78409, 5.784087, 5.784087, 5.784083, 5.784081, 
    5.784075, 5.784071, 5.784067, 5.784068, 5.784072, 5.784079, 5.784086, 
    5.784084, 5.784089, 5.784076, 5.784082, 5.78408, 5.784085, 5.784073, 
    5.784083, 5.78407, 5.784071, 5.784075, 5.784082, 5.784084, 5.784085, 
    5.784084, 5.78408, 5.784079, 5.784075, 5.784074, 5.784071, 5.784069, 
    5.784071, 5.784073, 5.78408, 5.784085, 5.784091, 5.784092, 5.784099, 
    5.784093, 5.784103, 5.784095, 5.784109, 5.784084, 5.784095, 5.784075, 
    5.784077, 5.784081, 5.78409, 5.784085, 5.784091, 5.784079, 5.784072, 
    5.78407, 5.784068, 5.78407, 5.78407, 5.784073, 5.784072, 5.78408, 
    5.784076, 5.784087, 5.784091, 5.784101, 5.784109, 5.784116, 5.784119, 
    5.78412, 5.78412 ;

 SOIL2C_TO_SOIL1C =
  1.086144e-09, 1.090923e-09, 1.089994e-09, 1.093849e-09, 1.091711e-09, 
    1.094235e-09, 1.087113e-09, 1.091113e-09, 1.088559e-09, 1.086574e-09, 
    1.101331e-09, 1.094021e-09, 1.108923e-09, 1.104261e-09, 1.115971e-09, 
    1.108197e-09, 1.117538e-09, 1.115746e-09, 1.121139e-09, 1.119594e-09, 
    1.126492e-09, 1.121852e-09, 1.130067e-09, 1.125384e-09, 1.126116e-09, 
    1.121699e-09, 1.095492e-09, 1.100421e-09, 1.0952e-09, 1.095903e-09, 
    1.095588e-09, 1.091755e-09, 1.089824e-09, 1.085778e-09, 1.086513e-09, 
    1.089484e-09, 1.096219e-09, 1.093933e-09, 1.099694e-09, 1.099564e-09, 
    1.105979e-09, 1.103087e-09, 1.113868e-09, 1.110804e-09, 1.119659e-09, 
    1.117432e-09, 1.119554e-09, 1.11891e-09, 1.119562e-09, 1.116296e-09, 
    1.117696e-09, 1.114822e-09, 1.103628e-09, 1.106918e-09, 1.097107e-09, 
    1.091207e-09, 1.087288e-09, 1.084508e-09, 1.084901e-09, 1.08565e-09, 
    1.089501e-09, 1.093122e-09, 1.095881e-09, 1.097727e-09, 1.099546e-09, 
    1.105051e-09, 1.107964e-09, 1.114488e-09, 1.11331e-09, 1.115305e-09, 
    1.11721e-09, 1.120409e-09, 1.119883e-09, 1.121292e-09, 1.115252e-09, 
    1.119266e-09, 1.11264e-09, 1.114452e-09, 1.100041e-09, 1.094549e-09, 
    1.092216e-09, 1.090173e-09, 1.085203e-09, 1.088635e-09, 1.087282e-09, 
    1.090501e-09, 1.092546e-09, 1.091535e-09, 1.097778e-09, 1.09535e-09, 
    1.108137e-09, 1.102629e-09, 1.116988e-09, 1.113552e-09, 1.117812e-09, 
    1.115638e-09, 1.119362e-09, 1.11601e-09, 1.121817e-09, 1.123081e-09, 
    1.122217e-09, 1.125536e-09, 1.115825e-09, 1.119554e-09, 1.091506e-09, 
    1.091671e-09, 1.09244e-09, 1.089061e-09, 1.088855e-09, 1.085758e-09, 
    1.088513e-09, 1.089687e-09, 1.092665e-09, 1.094426e-09, 1.096101e-09, 
    1.099782e-09, 1.103894e-09, 1.109644e-09, 1.113775e-09, 1.116544e-09, 
    1.114846e-09, 1.116345e-09, 1.114669e-09, 1.113884e-09, 1.122607e-09, 
    1.117709e-09, 1.125058e-09, 1.124651e-09, 1.121325e-09, 1.124697e-09, 
    1.091787e-09, 1.090838e-09, 1.087542e-09, 1.090121e-09, 1.085421e-09, 
    1.088052e-09, 1.089565e-09, 1.095401e-09, 1.096683e-09, 1.097873e-09, 
    1.100221e-09, 1.103235e-09, 1.108522e-09, 1.113122e-09, 1.117321e-09, 
    1.117013e-09, 1.117122e-09, 1.11806e-09, 1.115736e-09, 1.118441e-09, 
    1.118895e-09, 1.117708e-09, 1.124597e-09, 1.122629e-09, 1.124643e-09, 
    1.123361e-09, 1.091146e-09, 1.092744e-09, 1.09188e-09, 1.093504e-09, 
    1.09236e-09, 1.097445e-09, 1.09897e-09, 1.106103e-09, 1.103175e-09, 
    1.107835e-09, 1.103649e-09, 1.10439e-09, 1.107987e-09, 1.103875e-09, 
    1.112868e-09, 1.106771e-09, 1.118096e-09, 1.112008e-09, 1.118478e-09, 
    1.117303e-09, 1.119248e-09, 1.12099e-09, 1.123182e-09, 1.127226e-09, 
    1.12629e-09, 1.129672e-09, 1.095125e-09, 1.097197e-09, 1.097015e-09, 
    1.099183e-09, 1.100787e-09, 1.104262e-09, 1.109837e-09, 1.10774e-09, 
    1.111589e-09, 1.112361e-09, 1.106515e-09, 1.110104e-09, 1.098584e-09, 
    1.100445e-09, 1.099337e-09, 1.095289e-09, 1.108224e-09, 1.101585e-09, 
    1.113843e-09, 1.110247e-09, 1.120742e-09, 1.115523e-09, 1.125774e-09, 
    1.130157e-09, 1.134281e-09, 1.139102e-09, 1.098328e-09, 1.09692e-09, 
    1.099441e-09, 1.102929e-09, 1.106164e-09, 1.110466e-09, 1.110906e-09, 
    1.111712e-09, 1.1138e-09, 1.115555e-09, 1.111967e-09, 1.115995e-09, 
    1.100877e-09, 1.1088e-09, 1.096388e-09, 1.100125e-09, 1.102723e-09, 
    1.101583e-09, 1.107501e-09, 1.108895e-09, 1.114563e-09, 1.111633e-09, 
    1.129075e-09, 1.121358e-09, 1.142772e-09, 1.136788e-09, 1.096428e-09, 
    1.098323e-09, 1.104918e-09, 1.10178e-09, 1.110753e-09, 1.112962e-09, 
    1.114758e-09, 1.117053e-09, 1.117301e-09, 1.118661e-09, 1.116432e-09, 
    1.118573e-09, 1.110475e-09, 1.114094e-09, 1.104164e-09, 1.106581e-09, 
    1.105469e-09, 1.104249e-09, 1.108013e-09, 1.112024e-09, 1.112109e-09, 
    1.113395e-09, 1.117019e-09, 1.11079e-09, 1.130072e-09, 1.118164e-09, 
    1.100389e-09, 1.104039e-09, 1.10456e-09, 1.103147e-09, 1.112741e-09, 
    1.109265e-09, 1.118628e-09, 1.116097e-09, 1.120243e-09, 1.118183e-09, 
    1.11788e-09, 1.115234e-09, 1.113586e-09, 1.109424e-09, 1.106037e-09, 
    1.103352e-09, 1.103976e-09, 1.106926e-09, 1.112269e-09, 1.117323e-09, 
    1.116216e-09, 1.119928e-09, 1.110103e-09, 1.114223e-09, 1.112631e-09, 
    1.116783e-09, 1.107685e-09, 1.115433e-09, 1.105704e-09, 1.106557e-09, 
    1.109196e-09, 1.114502e-09, 1.115676e-09, 1.11693e-09, 1.116156e-09, 
    1.112405e-09, 1.11179e-09, 1.109131e-09, 1.108397e-09, 1.106372e-09, 
    1.104694e-09, 1.106227e-09, 1.107836e-09, 1.112406e-09, 1.116525e-09, 
    1.121015e-09, 1.122114e-09, 1.127361e-09, 1.12309e-09, 1.130138e-09, 
    1.124146e-09, 1.134518e-09, 1.115881e-09, 1.12397e-09, 1.109316e-09, 
    1.110894e-09, 1.11375e-09, 1.120299e-09, 1.116763e-09, 1.120898e-09, 
    1.111766e-09, 1.107028e-09, 1.105802e-09, 1.103515e-09, 1.105854e-09, 
    1.105664e-09, 1.107903e-09, 1.107183e-09, 1.112558e-09, 1.109671e-09, 
    1.117872e-09, 1.120865e-09, 1.129317e-09, 1.134499e-09, 1.139773e-09, 
    1.142101e-09, 1.14281e-09, 1.143106e-09 ;

 SOIL2C_TO_SOIL3C =
  7.75817e-11, 7.79231e-11, 7.785673e-11, 7.813209e-11, 7.797934e-11, 
    7.815965e-11, 7.765092e-11, 7.793666e-11, 7.775425e-11, 7.761244e-11, 
    7.866648e-11, 7.814437e-11, 7.920876e-11, 7.887579e-11, 7.97122e-11, 
    7.915694e-11, 7.982415e-11, 7.969617e-11, 8.008135e-11, 7.9971e-11, 
    8.04637e-11, 8.013228e-11, 8.071908e-11, 8.038455e-11, 8.043689e-11, 
    8.012135e-11, 7.824943e-11, 7.860148e-11, 7.822858e-11, 7.827878e-11, 
    7.825626e-11, 7.79825e-11, 7.784455e-11, 7.755561e-11, 7.760807e-11, 
    7.782028e-11, 7.830135e-11, 7.813804e-11, 7.85496e-11, 7.854031e-11, 
    7.89985e-11, 7.879191e-11, 7.9562e-11, 7.934313e-11, 7.997561e-11, 
    7.981655e-11, 7.996814e-11, 7.992217e-11, 7.996874e-11, 7.973546e-11, 
    7.983541e-11, 7.963013e-11, 7.88306e-11, 7.906558e-11, 7.836476e-11, 
    7.794337e-11, 7.766345e-11, 7.746483e-11, 7.749291e-11, 7.754644e-11, 
    7.782152e-11, 7.808014e-11, 7.827723e-11, 7.840907e-11, 7.853897e-11, 
    7.893219e-11, 7.91403e-11, 7.960627e-11, 7.952217e-11, 7.966464e-11, 
    7.980073e-11, 8.002923e-11, 7.999161e-11, 8.009229e-11, 7.966087e-11, 
    7.994759e-11, 7.947427e-11, 7.960373e-11, 7.857432e-11, 7.81821e-11, 
    7.801541e-11, 7.786949e-11, 7.751449e-11, 7.775965e-11, 7.766301e-11, 
    7.789291e-11, 7.803901e-11, 7.796675e-11, 7.841268e-11, 7.823932e-11, 
    7.915263e-11, 7.875924e-11, 7.978485e-11, 7.953943e-11, 7.984367e-11, 
    7.968842e-11, 7.995445e-11, 7.971503e-11, 8.012975e-11, 8.022006e-11, 
    8.015835e-11, 8.039539e-11, 7.970176e-11, 7.996814e-11, 7.796473e-11, 
    7.797651e-11, 7.803141e-11, 7.779009e-11, 7.777533e-11, 7.755417e-11, 
    7.775095e-11, 7.783475e-11, 7.804747e-11, 7.81733e-11, 7.829291e-11, 
    7.85559e-11, 7.88496e-11, 7.926029e-11, 7.955533e-11, 7.975311e-11, 
    7.963184e-11, 7.973891e-11, 7.961921e-11, 7.956311e-11, 8.018622e-11, 
    7.983634e-11, 8.03613e-11, 8.033225e-11, 8.009468e-11, 8.033552e-11, 
    7.798479e-11, 7.791697e-11, 7.768153e-11, 7.786579e-11, 7.753009e-11, 
    7.7718e-11, 7.782605e-11, 7.824295e-11, 7.833453e-11, 7.841947e-11, 
    7.858721e-11, 7.880249e-11, 7.918013e-11, 7.95087e-11, 7.980864e-11, 
    7.978666e-11, 7.97944e-11, 7.986141e-11, 7.969543e-11, 7.988866e-11, 
    7.992109e-11, 7.98363e-11, 8.032836e-11, 8.018778e-11, 8.033163e-11, 
    8.02401e-11, 7.793902e-11, 7.805312e-11, 7.799146e-11, 7.810741e-11, 
    7.802572e-11, 7.838894e-11, 7.849783e-11, 7.900737e-11, 7.879825e-11, 
    7.913106e-11, 7.883205e-11, 7.888504e-11, 7.914193e-11, 7.884821e-11, 
    7.949059e-11, 7.905509e-11, 7.986402e-11, 7.942914e-11, 7.989127e-11, 
    7.980734e-11, 7.994629e-11, 8.007073e-11, 8.022729e-11, 8.051616e-11, 
    8.044927e-11, 8.069084e-11, 7.822322e-11, 7.837123e-11, 7.835819e-11, 
    7.851307e-11, 7.862761e-11, 7.887587e-11, 7.927405e-11, 7.912431e-11, 
    7.939919e-11, 7.945437e-11, 7.903676e-11, 7.929318e-11, 7.847027e-11, 
    7.860324e-11, 7.852406e-11, 7.82349e-11, 7.915883e-11, 7.868467e-11, 
    7.956021e-11, 7.930336e-11, 8.005299e-11, 7.968019e-11, 8.041245e-11, 
    8.07255e-11, 8.102009e-11, 8.13644e-11, 7.845199e-11, 7.835143e-11, 
    7.853149e-11, 7.878061e-11, 7.901174e-11, 7.931902e-11, 7.935046e-11, 
    7.940803e-11, 7.955714e-11, 7.968251e-11, 7.942624e-11, 7.971394e-11, 
    7.863408e-11, 7.919998e-11, 7.831342e-11, 7.858039e-11, 7.876592e-11, 
    7.868453e-11, 7.910719e-11, 7.920681e-11, 7.961163e-11, 7.940237e-11, 
    8.064824e-11, 8.009703e-11, 8.162654e-11, 8.119911e-11, 7.831629e-11, 
    7.845164e-11, 7.892271e-11, 7.869858e-11, 7.933953e-11, 7.94973e-11, 
    7.962556e-11, 7.978952e-11, 7.980721e-11, 7.990435e-11, 7.974517e-11, 
    7.989806e-11, 7.931968e-11, 7.957814e-11, 7.886886e-11, 7.90415e-11, 
    7.896207e-11, 7.887496e-11, 7.914382e-11, 7.943027e-11, 7.943638e-11, 
    7.952823e-11, 7.978709e-11, 7.934213e-11, 8.07194e-11, 7.986885e-11, 
    7.859923e-11, 7.885995e-11, 7.889717e-11, 7.879618e-11, 7.948149e-11, 
    7.923318e-11, 7.990198e-11, 7.972122e-11, 8.001739e-11, 7.987022e-11, 
    7.984857e-11, 7.965955e-11, 7.954187e-11, 7.924457e-11, 7.900266e-11, 
    7.881083e-11, 7.885543e-11, 7.906616e-11, 7.94478e-11, 7.980882e-11, 
    7.972973e-11, 7.999488e-11, 7.929306e-11, 7.958735e-11, 7.947362e-11, 
    7.977018e-11, 7.912034e-11, 7.967375e-11, 7.897888e-11, 7.90398e-11, 
    7.922825e-11, 7.960732e-11, 7.969117e-11, 7.978072e-11, 7.972546e-11, 
    7.945748e-11, 7.941357e-11, 7.922367e-11, 7.917124e-11, 7.902654e-11, 
    7.890674e-11, 7.90162e-11, 7.913115e-11, 7.945759e-11, 7.975177e-11, 
    8.007251e-11, 8.0151e-11, 8.052577e-11, 8.022071e-11, 8.072414e-11, 
    8.029614e-11, 8.103701e-11, 7.97058e-11, 8.028354e-11, 7.923683e-11, 
    7.934958e-11, 7.955355e-11, 8.002134e-11, 7.976879e-11, 8.006415e-11, 
    7.941185e-11, 7.907343e-11, 7.898586e-11, 7.882249e-11, 7.898959e-11, 
    7.8976e-11, 7.91359e-11, 7.908452e-11, 7.946842e-11, 7.926221e-11, 
    7.984803e-11, 8.006181e-11, 8.066553e-11, 8.103563e-11, 8.141236e-11, 
    8.157867e-11, 8.16293e-11, 8.165046e-11 ;

 SOIL2C_vr =
  20.00646, 20.00648, 20.00648, 20.00649, 20.00648, 20.00649, 20.00646, 
    20.00648, 20.00647, 20.00646, 20.00652, 20.00649, 20.00654, 20.00653, 
    20.00657, 20.00654, 20.00657, 20.00657, 20.00658, 20.00658, 20.0066, 
    20.00659, 20.00661, 20.0066, 20.0066, 20.00659, 20.00649, 20.00651, 
    20.00649, 20.0065, 20.00649, 20.00648, 20.00647, 20.00646, 20.00646, 
    20.00647, 20.0065, 20.00649, 20.00651, 20.00651, 20.00653, 20.00652, 
    20.00656, 20.00655, 20.00658, 20.00657, 20.00658, 20.00658, 20.00658, 
    20.00657, 20.00657, 20.00656, 20.00652, 20.00653, 20.0065, 20.00648, 
    20.00647, 20.00646, 20.00646, 20.00646, 20.00647, 20.00649, 20.0065, 
    20.0065, 20.00651, 20.00653, 20.00654, 20.00656, 20.00656, 20.00656, 
    20.00657, 20.00658, 20.00658, 20.00658, 20.00656, 20.00658, 20.00656, 
    20.00656, 20.00651, 20.00649, 20.00648, 20.00648, 20.00646, 20.00647, 
    20.00647, 20.00648, 20.00648, 20.00648, 20.0065, 20.00649, 20.00654, 
    20.00652, 20.00657, 20.00656, 20.00657, 20.00657, 20.00658, 20.00657, 
    20.00659, 20.00659, 20.00659, 20.0066, 20.00657, 20.00658, 20.00648, 
    20.00648, 20.00648, 20.00647, 20.00647, 20.00646, 20.00647, 20.00647, 
    20.00648, 20.00649, 20.0065, 20.00651, 20.00652, 20.00654, 20.00656, 
    20.00657, 20.00656, 20.00657, 20.00656, 20.00656, 20.00659, 20.00657, 
    20.0066, 20.0066, 20.00658, 20.0066, 20.00648, 20.00648, 20.00647, 
    20.00648, 20.00646, 20.00647, 20.00647, 20.00649, 20.0065, 20.0065, 
    20.00651, 20.00652, 20.00654, 20.00656, 20.00657, 20.00657, 20.00657, 
    20.00657, 20.00657, 20.00657, 20.00658, 20.00657, 20.0066, 20.00659, 
    20.0066, 20.00659, 20.00648, 20.00648, 20.00648, 20.00649, 20.00648, 
    20.0065, 20.00651, 20.00653, 20.00652, 20.00654, 20.00652, 20.00653, 
    20.00654, 20.00652, 20.00656, 20.00653, 20.00657, 20.00655, 20.00657, 
    20.00657, 20.00658, 20.00658, 20.00659, 20.00661, 20.0066, 20.00661, 
    20.00649, 20.0065, 20.0065, 20.00651, 20.00651, 20.00653, 20.00654, 
    20.00654, 20.00655, 20.00655, 20.00653, 20.00655, 20.00651, 20.00651, 
    20.00651, 20.00649, 20.00654, 20.00652, 20.00656, 20.00655, 20.00658, 
    20.00657, 20.0066, 20.00662, 20.00663, 20.00665, 20.0065, 20.0065, 
    20.00651, 20.00652, 20.00653, 20.00655, 20.00655, 20.00655, 20.00656, 
    20.00657, 20.00655, 20.00657, 20.00651, 20.00654, 20.0065, 20.00651, 
    20.00652, 20.00652, 20.00654, 20.00654, 20.00656, 20.00655, 20.00661, 
    20.00659, 20.00666, 20.00664, 20.0065, 20.0065, 20.00653, 20.00652, 
    20.00655, 20.00656, 20.00656, 20.00657, 20.00657, 20.00658, 20.00657, 
    20.00657, 20.00655, 20.00656, 20.00653, 20.00653, 20.00653, 20.00653, 
    20.00654, 20.00655, 20.00655, 20.00656, 20.00657, 20.00655, 20.00662, 
    20.00657, 20.00651, 20.00653, 20.00653, 20.00652, 20.00656, 20.00654, 
    20.00658, 20.00657, 20.00658, 20.00657, 20.00657, 20.00656, 20.00656, 
    20.00654, 20.00653, 20.00652, 20.00653, 20.00653, 20.00655, 20.00657, 
    20.00657, 20.00658, 20.00655, 20.00656, 20.00655, 20.00657, 20.00654, 
    20.00657, 20.00653, 20.00653, 20.00654, 20.00656, 20.00657, 20.00657, 
    20.00657, 20.00655, 20.00655, 20.00654, 20.00654, 20.00653, 20.00653, 
    20.00653, 20.00654, 20.00655, 20.00657, 20.00658, 20.00659, 20.00661, 
    20.00659, 20.00662, 20.0066, 20.00663, 20.00657, 20.00659, 20.00654, 
    20.00655, 20.00656, 20.00658, 20.00657, 20.00658, 20.00655, 20.00653, 
    20.00653, 20.00652, 20.00653, 20.00653, 20.00654, 20.00653, 20.00655, 
    20.00654, 20.00657, 20.00658, 20.00661, 20.00663, 20.00665, 20.00666, 
    20.00666, 20.00666,
  20.00607, 20.00609, 20.00609, 20.00611, 20.0061, 20.00611, 20.00607, 
    20.00609, 20.00608, 20.00607, 20.00614, 20.00611, 20.00618, 20.00616, 
    20.00621, 20.00617, 20.00622, 20.00621, 20.00624, 20.00623, 20.00626, 
    20.00624, 20.00628, 20.00626, 20.00626, 20.00624, 20.00611, 20.00614, 
    20.00611, 20.00612, 20.00611, 20.0061, 20.00609, 20.00607, 20.00607, 
    20.00609, 20.00612, 20.00611, 20.00613, 20.00613, 20.00616, 20.00615, 
    20.0062, 20.00619, 20.00623, 20.00622, 20.00623, 20.00623, 20.00623, 
    20.00621, 20.00622, 20.00621, 20.00615, 20.00617, 20.00612, 20.00609, 
    20.00607, 20.00606, 20.00606, 20.00607, 20.00609, 20.0061, 20.00612, 
    20.00612, 20.00613, 20.00616, 20.00617, 20.0062, 20.0062, 20.00621, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00621, 20.00623, 20.0062, 
    20.0062, 20.00614, 20.00611, 20.0061, 20.00609, 20.00607, 20.00608, 
    20.00607, 20.00609, 20.0061, 20.0061, 20.00612, 20.00611, 20.00617, 
    20.00615, 20.00622, 20.0062, 20.00622, 20.00621, 20.00623, 20.00621, 
    20.00624, 20.00624, 20.00624, 20.00626, 20.00621, 20.00623, 20.0061, 
    20.0061, 20.0061, 20.00608, 20.00608, 20.00607, 20.00608, 20.00609, 
    20.0061, 20.00611, 20.00612, 20.00613, 20.00615, 20.00618, 20.0062, 
    20.00621, 20.00621, 20.00621, 20.0062, 20.0062, 20.00624, 20.00622, 
    20.00625, 20.00625, 20.00624, 20.00625, 20.0061, 20.00609, 20.00608, 
    20.00609, 20.00607, 20.00608, 20.00609, 20.00611, 20.00612, 20.00612, 
    20.00614, 20.00615, 20.00618, 20.0062, 20.00622, 20.00622, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00623, 20.00622, 20.00625, 20.00624, 
    20.00625, 20.00625, 20.00609, 20.0061, 20.0061, 20.00611, 20.0061, 
    20.00612, 20.00613, 20.00616, 20.00615, 20.00617, 20.00615, 20.00616, 
    20.00617, 20.00615, 20.0062, 20.00617, 20.00622, 20.00619, 20.00622, 
    20.00622, 20.00623, 20.00624, 20.00624, 20.00626, 20.00626, 20.00628, 
    20.00611, 20.00612, 20.00612, 20.00613, 20.00614, 20.00616, 20.00618, 
    20.00617, 20.00619, 20.00619, 20.00617, 20.00618, 20.00613, 20.00614, 
    20.00613, 20.00611, 20.00617, 20.00614, 20.0062, 20.00618, 20.00623, 
    20.00621, 20.00626, 20.00628, 20.0063, 20.00632, 20.00613, 20.00612, 
    20.00613, 20.00615, 20.00616, 20.00619, 20.00619, 20.00619, 20.0062, 
    20.00621, 20.00619, 20.00621, 20.00614, 20.00618, 20.00612, 20.00614, 
    20.00615, 20.00614, 20.00617, 20.00618, 20.0062, 20.00619, 20.00627, 
    20.00624, 20.00634, 20.00631, 20.00612, 20.00613, 20.00616, 20.00614, 
    20.00619, 20.0062, 20.0062, 20.00622, 20.00622, 20.00622, 20.00621, 
    20.00622, 20.00619, 20.0062, 20.00616, 20.00617, 20.00616, 20.00616, 
    20.00617, 20.00619, 20.00619, 20.0062, 20.00622, 20.00619, 20.00628, 
    20.00622, 20.00614, 20.00616, 20.00616, 20.00615, 20.0062, 20.00618, 
    20.00622, 20.00621, 20.00623, 20.00622, 20.00622, 20.00621, 20.0062, 
    20.00618, 20.00616, 20.00615, 20.00616, 20.00617, 20.00619, 20.00622, 
    20.00621, 20.00623, 20.00618, 20.0062, 20.0062, 20.00621, 20.00617, 
    20.00621, 20.00616, 20.00617, 20.00618, 20.0062, 20.00621, 20.00622, 
    20.00621, 20.0062, 20.00619, 20.00618, 20.00618, 20.00617, 20.00616, 
    20.00616, 20.00617, 20.0062, 20.00621, 20.00624, 20.00624, 20.00627, 
    20.00624, 20.00628, 20.00625, 20.0063, 20.00621, 20.00625, 20.00618, 
    20.00619, 20.0062, 20.00623, 20.00621, 20.00624, 20.00619, 20.00617, 
    20.00616, 20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.0062, 
    20.00618, 20.00622, 20.00623, 20.00627, 20.0063, 20.00632, 20.00633, 
    20.00634, 20.00634,
  20.00552, 20.00554, 20.00554, 20.00556, 20.00555, 20.00556, 20.00552, 
    20.00554, 20.00553, 20.00552, 20.0056, 20.00556, 20.00563, 20.00561, 
    20.00567, 20.00563, 20.00568, 20.00567, 20.0057, 20.00569, 20.00572, 
    20.0057, 20.00574, 20.00572, 20.00572, 20.0057, 20.00557, 20.00559, 
    20.00557, 20.00557, 20.00557, 20.00555, 20.00554, 20.00552, 20.00552, 
    20.00554, 20.00557, 20.00556, 20.00559, 20.00559, 20.00562, 20.00561, 
    20.00566, 20.00564, 20.00569, 20.00568, 20.00569, 20.00569, 20.00569, 
    20.00567, 20.00568, 20.00566, 20.00561, 20.00562, 20.00558, 20.00554, 
    20.00553, 20.00551, 20.00551, 20.00552, 20.00554, 20.00555, 20.00557, 
    20.00558, 20.00559, 20.00562, 20.00563, 20.00566, 20.00566, 20.00567, 
    20.00568, 20.00569, 20.00569, 20.0057, 20.00567, 20.00569, 20.00565, 
    20.00566, 20.00559, 20.00556, 20.00555, 20.00554, 20.00551, 20.00553, 
    20.00553, 20.00554, 20.00555, 20.00555, 20.00558, 20.00557, 20.00563, 
    20.0056, 20.00567, 20.00566, 20.00568, 20.00567, 20.00569, 20.00567, 
    20.0057, 20.00571, 20.0057, 20.00572, 20.00567, 20.00569, 20.00555, 
    20.00555, 20.00555, 20.00553, 20.00553, 20.00552, 20.00553, 20.00554, 
    20.00555, 20.00556, 20.00557, 20.00559, 20.00561, 20.00564, 20.00566, 
    20.00567, 20.00566, 20.00567, 20.00566, 20.00566, 20.0057, 20.00568, 
    20.00572, 20.00571, 20.0057, 20.00571, 20.00555, 20.00554, 20.00553, 
    20.00554, 20.00552, 20.00553, 20.00554, 20.00557, 20.00557, 20.00558, 
    20.00559, 20.00561, 20.00563, 20.00566, 20.00568, 20.00568, 20.00568, 
    20.00568, 20.00567, 20.00568, 20.00569, 20.00568, 20.00571, 20.0057, 
    20.00571, 20.00571, 20.00554, 20.00555, 20.00555, 20.00556, 20.00555, 
    20.00558, 20.00558, 20.00562, 20.00561, 20.00563, 20.00561, 20.00561, 
    20.00563, 20.00561, 20.00566, 20.00562, 20.00568, 20.00565, 20.00568, 
    20.00568, 20.00569, 20.0057, 20.00571, 20.00573, 20.00572, 20.00574, 
    20.00557, 20.00558, 20.00558, 20.00558, 20.00559, 20.00561, 20.00564, 
    20.00563, 20.00565, 20.00565, 20.00562, 20.00564, 20.00558, 20.00559, 
    20.00559, 20.00557, 20.00563, 20.0056, 20.00566, 20.00564, 20.00569, 
    20.00567, 20.00572, 20.00574, 20.00576, 20.00579, 20.00558, 20.00557, 
    20.00559, 20.0056, 20.00562, 20.00564, 20.00564, 20.00565, 20.00566, 
    20.00567, 20.00565, 20.00567, 20.00559, 20.00563, 20.00557, 20.00559, 
    20.0056, 20.0056, 20.00563, 20.00563, 20.00566, 20.00565, 20.00574, 
    20.0057, 20.00581, 20.00578, 20.00557, 20.00558, 20.00562, 20.0056, 
    20.00564, 20.00566, 20.00566, 20.00568, 20.00568, 20.00568, 20.00567, 
    20.00568, 20.00564, 20.00566, 20.00561, 20.00562, 20.00562, 20.00561, 
    20.00563, 20.00565, 20.00565, 20.00566, 20.00568, 20.00564, 20.00574, 
    20.00568, 20.00559, 20.00561, 20.00561, 20.00561, 20.00565, 20.00564, 
    20.00568, 20.00567, 20.00569, 20.00568, 20.00568, 20.00567, 20.00566, 
    20.00564, 20.00562, 20.00561, 20.00561, 20.00562, 20.00565, 20.00568, 
    20.00567, 20.00569, 20.00564, 20.00566, 20.00565, 20.00567, 20.00563, 
    20.00567, 20.00562, 20.00562, 20.00564, 20.00566, 20.00567, 20.00567, 
    20.00567, 20.00565, 20.00565, 20.00564, 20.00563, 20.00562, 20.00561, 
    20.00562, 20.00563, 20.00565, 20.00567, 20.0057, 20.0057, 20.00573, 
    20.00571, 20.00574, 20.00571, 20.00576, 20.00567, 20.00571, 20.00564, 
    20.00564, 20.00566, 20.00569, 20.00567, 20.0057, 20.00565, 20.00562, 
    20.00562, 20.00561, 20.00562, 20.00562, 20.00563, 20.00563, 20.00565, 
    20.00564, 20.00568, 20.0057, 20.00574, 20.00576, 20.00579, 20.0058, 
    20.00581, 20.00581,
  20.00508, 20.0051, 20.0051, 20.00512, 20.00511, 20.00512, 20.00508, 
    20.00511, 20.00509, 20.00508, 20.00516, 20.00512, 20.00519, 20.00517, 
    20.00523, 20.00519, 20.00524, 20.00523, 20.00525, 20.00525, 20.00528, 
    20.00526, 20.0053, 20.00528, 20.00528, 20.00526, 20.00513, 20.00515, 
    20.00513, 20.00513, 20.00513, 20.00511, 20.0051, 20.00508, 20.00508, 
    20.0051, 20.00513, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 
    20.00522, 20.0052, 20.00525, 20.00524, 20.00525, 20.00525, 20.00525, 
    20.00523, 20.00524, 20.00522, 20.00517, 20.00518, 20.00513, 20.00511, 
    20.00508, 20.00507, 20.00507, 20.00508, 20.0051, 20.00512, 20.00513, 
    20.00514, 20.00515, 20.00517, 20.00519, 20.00522, 20.00522, 20.00523, 
    20.00524, 20.00525, 20.00525, 20.00526, 20.00523, 20.00525, 20.00521, 
    20.00522, 20.00515, 20.00512, 20.00511, 20.0051, 20.00508, 20.00509, 
    20.00508, 20.0051, 20.00511, 20.00511, 20.00514, 20.00513, 20.00519, 
    20.00516, 20.00524, 20.00522, 20.00524, 20.00523, 20.00525, 20.00523, 
    20.00526, 20.00527, 20.00526, 20.00528, 20.00523, 20.00525, 20.00511, 
    20.00511, 20.00511, 20.00509, 20.00509, 20.00508, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00513, 20.00515, 20.00517, 20.0052, 20.00522, 
    20.00523, 20.00522, 20.00523, 20.00522, 20.00522, 20.00526, 20.00524, 
    20.00528, 20.00527, 20.00526, 20.00527, 20.00511, 20.0051, 20.00509, 
    20.0051, 20.00508, 20.00509, 20.0051, 20.00513, 20.00513, 20.00514, 
    20.00515, 20.00517, 20.00519, 20.00521, 20.00524, 20.00524, 20.00524, 
    20.00524, 20.00523, 20.00524, 20.00525, 20.00524, 20.00527, 20.00526, 
    20.00527, 20.00527, 20.00511, 20.00511, 20.00511, 20.00512, 20.00511, 
    20.00514, 20.00514, 20.00518, 20.00517, 20.00519, 20.00517, 20.00517, 
    20.00519, 20.00517, 20.00521, 20.00518, 20.00524, 20.00521, 20.00524, 
    20.00524, 20.00525, 20.00525, 20.00527, 20.00529, 20.00528, 20.0053, 
    20.00513, 20.00514, 20.00513, 20.00515, 20.00515, 20.00517, 20.0052, 
    20.00519, 20.00521, 20.00521, 20.00518, 20.0052, 20.00514, 20.00515, 
    20.00515, 20.00513, 20.00519, 20.00516, 20.00522, 20.0052, 20.00525, 
    20.00523, 20.00528, 20.0053, 20.00532, 20.00535, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00518, 20.0052, 20.00521, 20.00521, 20.00522, 
    20.00523, 20.00521, 20.00523, 20.00515, 20.00519, 20.00513, 20.00515, 
    20.00516, 20.00516, 20.00519, 20.00519, 20.00522, 20.00521, 20.00529, 
    20.00526, 20.00536, 20.00533, 20.00513, 20.00514, 20.00517, 20.00516, 
    20.0052, 20.00521, 20.00522, 20.00524, 20.00524, 20.00524, 20.00523, 
    20.00524, 20.0052, 20.00522, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00519, 20.00521, 20.00521, 20.00522, 20.00524, 20.0052, 20.0053, 
    20.00524, 20.00515, 20.00517, 20.00517, 20.00517, 20.00521, 20.0052, 
    20.00524, 20.00523, 20.00525, 20.00524, 20.00524, 20.00523, 20.00522, 
    20.0052, 20.00518, 20.00517, 20.00517, 20.00518, 20.00521, 20.00524, 
    20.00523, 20.00525, 20.0052, 20.00522, 20.00521, 20.00523, 20.00519, 
    20.00523, 20.00518, 20.00518, 20.0052, 20.00522, 20.00523, 20.00523, 
    20.00523, 20.00521, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00518, 20.00519, 20.00521, 20.00523, 20.00525, 20.00526, 20.00529, 
    20.00527, 20.0053, 20.00527, 20.00532, 20.00523, 20.00527, 20.0052, 
    20.00521, 20.00522, 20.00525, 20.00523, 20.00525, 20.00521, 20.00518, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00519, 20.00519, 20.00521, 
    20.0052, 20.00524, 20.00525, 20.0053, 20.00532, 20.00535, 20.00536, 
    20.00536, 20.00537,
  20.00437, 20.00439, 20.00439, 20.0044, 20.00439, 20.00441, 20.00438, 
    20.00439, 20.00438, 20.00437, 20.00444, 20.0044, 20.00447, 20.00445, 
    20.0045, 20.00447, 20.00451, 20.0045, 20.00452, 20.00451, 20.00454, 
    20.00452, 20.00456, 20.00454, 20.00454, 20.00452, 20.00441, 20.00443, 
    20.00441, 20.00441, 20.00441, 20.00439, 20.00439, 20.00437, 20.00437, 
    20.00438, 20.00441, 20.0044, 20.00443, 20.00443, 20.00446, 20.00444, 
    20.00449, 20.00448, 20.00451, 20.00451, 20.00451, 20.00451, 20.00451, 
    20.0045, 20.00451, 20.00449, 20.00445, 20.00446, 20.00442, 20.00439, 
    20.00438, 20.00436, 20.00437, 20.00437, 20.00438, 20.0044, 20.00441, 
    20.00442, 20.00443, 20.00445, 20.00446, 20.00449, 20.00449, 20.0045, 
    20.0045, 20.00452, 20.00451, 20.00452, 20.0045, 20.00451, 20.00448, 
    20.00449, 20.00443, 20.00441, 20.0044, 20.00439, 20.00437, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.00439, 20.00442, 20.00441, 20.00447, 
    20.00444, 20.0045, 20.00449, 20.00451, 20.0045, 20.00451, 20.0045, 
    20.00452, 20.00453, 20.00452, 20.00454, 20.0045, 20.00451, 20.00439, 
    20.00439, 20.0044, 20.00438, 20.00438, 20.00437, 20.00438, 20.00439, 
    20.0044, 20.00441, 20.00441, 20.00443, 20.00445, 20.00447, 20.00449, 
    20.0045, 20.00449, 20.0045, 20.00449, 20.00449, 20.00453, 20.00451, 
    20.00454, 20.00454, 20.00452, 20.00454, 20.00439, 20.00439, 20.00438, 
    20.00439, 20.00437, 20.00438, 20.00438, 20.00441, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00447, 20.00449, 20.0045, 20.0045, 20.0045, 
    20.00451, 20.0045, 20.00451, 20.00451, 20.00451, 20.00454, 20.00453, 
    20.00454, 20.00453, 20.00439, 20.0044, 20.00439, 20.0044, 20.0044, 
    20.00442, 20.00443, 20.00446, 20.00444, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00445, 20.00448, 20.00446, 20.00451, 20.00448, 20.00451, 
    20.0045, 20.00451, 20.00452, 20.00453, 20.00455, 20.00454, 20.00456, 
    20.00441, 20.00442, 20.00442, 20.00443, 20.00443, 20.00445, 20.00447, 
    20.00446, 20.00448, 20.00448, 20.00446, 20.00447, 20.00442, 20.00443, 
    20.00443, 20.00441, 20.00447, 20.00444, 20.00449, 20.00447, 20.00452, 
    20.0045, 20.00454, 20.00456, 20.00458, 20.0046, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00446, 20.00447, 20.00448, 20.00448, 20.00449, 
    20.0045, 20.00448, 20.0045, 20.00443, 20.00447, 20.00442, 20.00443, 
    20.00444, 20.00444, 20.00446, 20.00447, 20.00449, 20.00448, 20.00455, 
    20.00452, 20.00461, 20.00459, 20.00442, 20.00442, 20.00445, 20.00444, 
    20.00448, 20.00449, 20.00449, 20.0045, 20.0045, 20.00451, 20.0045, 
    20.00451, 20.00447, 20.00449, 20.00445, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00448, 20.00448, 20.00449, 20.0045, 20.00448, 20.00456, 
    20.00451, 20.00443, 20.00445, 20.00445, 20.00444, 20.00448, 20.00447, 
    20.00451, 20.0045, 20.00452, 20.00451, 20.00451, 20.0045, 20.00449, 
    20.00447, 20.00446, 20.00444, 20.00445, 20.00446, 20.00448, 20.0045, 
    20.0045, 20.00451, 20.00447, 20.00449, 20.00448, 20.0045, 20.00446, 
    20.0045, 20.00445, 20.00446, 20.00447, 20.00449, 20.0045, 20.0045, 
    20.0045, 20.00448, 20.00448, 20.00447, 20.00447, 20.00446, 20.00445, 
    20.00446, 20.00446, 20.00448, 20.0045, 20.00452, 20.00452, 20.00455, 
    20.00453, 20.00456, 20.00453, 20.00458, 20.0045, 20.00453, 20.00447, 
    20.00448, 20.00449, 20.00452, 20.0045, 20.00452, 20.00448, 20.00446, 
    20.00446, 20.00444, 20.00446, 20.00445, 20.00446, 20.00446, 20.00448, 
    20.00447, 20.00451, 20.00452, 20.00455, 20.00458, 20.0046, 20.00461, 
    20.00461, 20.00461,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258222, 0.5258228, 0.5258227, 0.5258232, 0.5258229, 0.5258232, 
    0.5258223, 0.5258228, 0.5258225, 0.5258223, 0.5258241, 0.5258232, 
    0.525825, 0.5258244, 0.5258258, 0.5258249, 0.525826, 0.5258258, 
    0.5258265, 0.5258263, 0.5258271, 0.5258265, 0.5258275, 0.5258269, 
    0.5258271, 0.5258265, 0.5258234, 0.525824, 0.5258233, 0.5258234, 
    0.5258234, 0.5258229, 0.5258227, 0.5258222, 0.5258223, 0.5258226, 
    0.5258235, 0.5258232, 0.5258239, 0.5258238, 0.5258246, 0.5258242, 
    0.5258256, 0.5258252, 0.5258263, 0.525826, 0.5258263, 0.5258262, 
    0.5258263, 0.5258259, 0.525826, 0.5258257, 0.5258243, 0.5258247, 
    0.5258235, 0.5258228, 0.5258223, 0.525822, 0.5258221, 0.5258222, 
    0.5258226, 0.5258231, 0.5258234, 0.5258237, 0.5258238, 0.5258245, 
    0.5258248, 0.5258256, 0.5258255, 0.5258257, 0.525826, 0.5258263, 
    0.5258263, 0.5258265, 0.5258257, 0.5258262, 0.5258254, 0.5258256, 
    0.5258239, 0.5258232, 0.5258229, 0.5258227, 0.5258221, 0.5258225, 
    0.5258223, 0.5258228, 0.525823, 0.5258229, 0.5258237, 0.5258234, 
    0.5258249, 0.5258242, 0.5258259, 0.5258256, 0.525826, 0.5258258, 
    0.5258262, 0.5258258, 0.5258265, 0.5258267, 0.5258266, 0.525827, 
    0.5258258, 0.5258263, 0.5258229, 0.5258229, 0.525823, 0.5258226, 
    0.5258226, 0.5258222, 0.5258225, 0.5258226, 0.525823, 0.5258232, 
    0.5258234, 0.5258239, 0.5258244, 0.5258251, 0.5258256, 0.5258259, 
    0.5258257, 0.5258259, 0.5258257, 0.5258256, 0.5258266, 0.525826, 
    0.5258269, 0.5258269, 0.5258265, 0.5258269, 0.5258229, 0.5258228, 
    0.5258224, 0.5258227, 0.5258222, 0.5258225, 0.5258226, 0.5258234, 
    0.5258235, 0.5258237, 0.525824, 0.5258243, 0.5258249, 0.5258255, 
    0.525826, 0.525826, 0.525826, 0.5258261, 0.5258258, 0.5258261, 0.5258262, 
    0.525826, 0.5258269, 0.5258266, 0.5258269, 0.5258267, 0.5258228, 
    0.525823, 0.5258229, 0.5258231, 0.525823, 0.5258236, 0.5258238, 
    0.5258246, 0.5258243, 0.5258248, 0.5258244, 0.5258244, 0.5258248, 
    0.5258244, 0.5258254, 0.5258247, 0.5258261, 0.5258253, 0.5258261, 
    0.525826, 0.5258262, 0.5258265, 0.5258267, 0.5258272, 0.5258271, 
    0.5258275, 0.5258233, 0.5258235, 0.5258235, 0.5258238, 0.525824, 
    0.5258244, 0.5258251, 0.5258248, 0.5258253, 0.5258254, 0.5258247, 
    0.5258251, 0.5258237, 0.525824, 0.5258238, 0.5258234, 0.5258249, 
    0.5258241, 0.5258256, 0.5258251, 0.5258264, 0.5258258, 0.525827, 
    0.5258275, 0.525828, 0.5258286, 0.5258237, 0.5258235, 0.5258238, 
    0.5258242, 0.5258247, 0.5258251, 0.5258252, 0.5258253, 0.5258256, 
    0.5258258, 0.5258253, 0.5258258, 0.525824, 0.525825, 0.5258235, 
    0.5258239, 0.5258242, 0.5258241, 0.5258248, 0.525825, 0.5258257, 
    0.5258253, 0.5258274, 0.5258265, 0.5258291, 0.5258283, 0.5258235, 
    0.5258237, 0.5258245, 0.5258241, 0.5258252, 0.5258254, 0.5258257, 
    0.525826, 0.525826, 0.5258262, 0.5258259, 0.5258262, 0.5258251, 
    0.5258256, 0.5258244, 0.5258247, 0.5258245, 0.5258244, 0.5258248, 
    0.5258253, 0.5258254, 0.5258255, 0.525826, 0.5258252, 0.5258275, 
    0.5258261, 0.525824, 0.5258244, 0.5258244, 0.5258243, 0.5258254, 
    0.525825, 0.5258262, 0.5258259, 0.5258263, 0.5258261, 0.525826, 
    0.5258257, 0.5258256, 0.525825, 0.5258246, 0.5258243, 0.5258244, 
    0.5258247, 0.5258254, 0.525826, 0.5258259, 0.5258263, 0.5258251, 
    0.5258256, 0.5258254, 0.5258259, 0.5258248, 0.5258257, 0.5258246, 
    0.5258247, 0.525825, 0.5258256, 0.5258258, 0.5258259, 0.5258259, 
    0.5258254, 0.5258253, 0.525825, 0.5258249, 0.5258247, 0.5258245, 
    0.5258247, 0.5258248, 0.5258254, 0.5258259, 0.5258265, 0.5258266, 
    0.5258272, 0.5258267, 0.5258275, 0.5258268, 0.5258281, 0.5258258, 
    0.5258268, 0.525825, 0.5258252, 0.5258256, 0.5258263, 0.5258259, 
    0.5258264, 0.5258253, 0.5258247, 0.5258246, 0.5258243, 0.5258246, 
    0.5258246, 0.5258248, 0.5258248, 0.5258254, 0.5258251, 0.525826, 
    0.5258264, 0.5258274, 0.5258281, 0.5258287, 0.525829, 0.5258291, 0.5258291 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -2.569961e-21, -7.709882e-21, 1.28498e-20, 2.055969e-20, -7.709882e-21, 
    1.28498e-20, 2.055969e-20, -1.541976e-20, 2.055969e-20, 0, 7.709882e-21, 
    1.027984e-20, -5.139921e-21, -7.709882e-21, -1.28498e-20, 7.709882e-21, 
    -1.027984e-20, 1.027984e-20, -7.709882e-21, 1.003089e-36, 5.139921e-21, 
    2.569961e-20, 5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, 2.312965e-20, 1.027984e-20, 
    7.709882e-21, -2.312965e-20, -5.139921e-21, 3.340949e-20, 0, 
    -5.139921e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, -2.569961e-21, -1.541976e-20, 1.541976e-20, 
    -7.709882e-21, -7.709882e-21, 7.709882e-21, 1.027984e-20, -1.28498e-20, 
    -5.139921e-21, 1.027984e-20, 7.709882e-21, 7.709882e-21, 2.569961e-20, 
    -5.139921e-21, 1.28498e-20, 1.027984e-20, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, -1.003089e-36, 1.027984e-20, -1.003089e-36, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, -1.28498e-20, 
    -1.541976e-20, 7.709882e-21, 1.798972e-20, -5.139921e-21, -2.569961e-21, 
    2.055969e-20, -7.709882e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    2.569961e-20, 1.798972e-20, -7.709882e-21, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 1.798972e-20, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -7.709882e-21, 7.709882e-21, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, 7.709882e-21, 2.569961e-20, -1.027984e-20, 
    -1.003089e-36, -1.541976e-20, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    1.003089e-36, -5.139921e-21, 1.027984e-20, -1.541976e-20, 2.569961e-21, 
    -2.569961e-21, -1.28498e-20, -5.139921e-21, 1.541976e-20, 0, 
    1.541976e-20, -5.139921e-21, 2.569961e-21, -7.709882e-21, 1.003089e-36, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 0, -1.027984e-20, 
    -1.28498e-20, 1.027984e-20, -1.003089e-36, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, 1.003089e-36, 7.709882e-21, 
    1.027984e-20, 5.139921e-21, -7.709882e-21, -2.569961e-21, -1.027984e-20, 
    -1.28498e-20, -2.569961e-21, 1.798972e-20, 5.139921e-21, -1.28498e-20, 
    1.28498e-20, -2.569961e-21, 0, -1.027984e-20, -1.798972e-20, 
    -5.139921e-21, 0, -2.569961e-21, -1.798972e-20, 2.569961e-21, 
    -1.798972e-20, 2.569961e-21, 7.709882e-21, -2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 1.541976e-20, 1.28498e-20, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 1.541976e-20, 0, 7.709882e-21, 
    -1.541976e-20, -1.28498e-20, 2.569961e-21, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, 1.003089e-36, 1.28498e-20, 1.541976e-20, 
    -1.28498e-20, 2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.541976e-20, 1.28498e-20, -2.569961e-21, -1.28498e-20, 1.003089e-36, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -7.709882e-21, 1.28498e-20, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    1.28498e-20, 5.139921e-21, 0, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -2.569961e-21, -1.003089e-36, 2.312965e-20, -1.28498e-20, -7.709882e-21, 
    -1.798972e-20, 1.541976e-20, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 1.798972e-20, -1.28498e-20, -5.139921e-21, 
    -1.541976e-20, -2.569961e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 1.28498e-20, -1.798972e-20, 
    -1.28498e-20, 1.798972e-20, 2.569961e-21, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, -5.139921e-21, -2.312965e-20, -1.541976e-20, 5.139921e-21, 
    -1.027984e-20, 7.709882e-21, -1.28498e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, 0, -1.798972e-20, 2.569961e-21, 5.139921e-21, 1.798972e-20, 
    1.003089e-36, -5.139921e-21, 1.541976e-20, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, -1.027984e-20, 1.541976e-20, 1.798972e-20, 
    1.541976e-20, 2.569961e-21, -1.027984e-20, 7.709882e-21, 2.569961e-21, 
    -1.003089e-36, -1.541976e-20, -2.312965e-20, 2.569961e-21, -5.139921e-21, 
    -1.003089e-36, -1.798972e-20, 7.709882e-21, -1.003089e-36, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, -1.798972e-20, 7.709882e-21, 
    0, -5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, -5.139921e-21, 1.541976e-20, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.798972e-20, 5.139921e-21, -1.28498e-20, 
    -1.027984e-20, -1.28498e-20, 1.027984e-20, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -2.055969e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, 1.798972e-20,
  -2.569961e-21, -5.139921e-21, 7.709882e-21, -1.541976e-20, 5.139921e-21, 
    -1.28498e-20, 1.027984e-20, 2.569961e-21, -1.003089e-36, 1.027984e-20, 
    -2.569961e-21, -1.541976e-20, 1.28498e-20, -1.027984e-20, -1.027984e-20, 
    -1.28498e-20, -7.709882e-21, 0, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 0, 2.569961e-21, 1.003089e-36, -7.709882e-21, 
    1.003089e-36, -7.709882e-21, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, -1.027984e-20, 2.569961e-21, 0, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 2.569961e-21, 
    0, 0, 1.027984e-20, 1.003089e-36, 0, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -1.28498e-20, -1.003089e-36, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 1.798972e-20, 
    -2.569961e-21, -5.139921e-21, 0, -1.027984e-20, 1.027984e-20, 
    -7.709882e-21, 0, -1.003089e-36, 7.709882e-21, 1.027984e-20, 0, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 1.003089e-36, -1.28498e-20, 
    0, 7.709882e-21, -5.139921e-21, 0, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, -1.027984e-20, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, 
    -1.541976e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    1.003089e-36, -5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 1.28498e-20, -2.569961e-21, -5.139921e-21, -3.083953e-20, 
    1.027984e-20, -2.569961e-21, -1.027984e-20, 0, 5.139921e-21, 0, 
    -1.027984e-20, -2.569961e-21, 2.569961e-21, -1.28498e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, 2.055969e-20, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 1.003089e-36, 1.003089e-36, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 
    1.027984e-20, -7.709882e-21, 1.027984e-20, 7.709882e-21, -2.569961e-21, 
    7.709882e-21, 0, 1.28498e-20, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    0, 0, 5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    2.569961e-21, -1.28498e-20, -1.027984e-20, 5.139921e-21, 0, 7.709882e-21, 
    -1.003089e-36, -1.003089e-36, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 1.28498e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    0, 1.027984e-20, -1.027984e-20, 0, -2.569961e-21, 0, -1.003089e-36, 0, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, 0, 0, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, 1.541976e-20, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -1.027984e-20, 1.003089e-36, 1.003089e-36, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, 0, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 1.003089e-36, 
    1.003089e-36, -1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, 0, 
    -1.28498e-20, 1.28498e-20, 1.027984e-20, -1.027984e-20, 0, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -1.003089e-36, -1.003089e-36, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 7.709882e-21, -1.28498e-20, -1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, 0, 2.569961e-21, 
    7.709882e-21, 1.28498e-20, 0, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    -2.569961e-21, 1.28498e-20, -1.027984e-20, -5.139921e-21, 1.003089e-36, 
    2.055969e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 0, 2.569961e-21, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -2.569961e-21, 0, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 1.541976e-20, 7.709882e-21, 7.709882e-21,
  5.139921e-21, -2.569961e-21, 7.709882e-21, 1.003089e-36, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, 0, 0, -2.569961e-21, 1.027984e-20, 
    1.798972e-20, -2.569961e-21, 1.027984e-20, 0, -1.28498e-20, 
    -1.798972e-20, 7.709882e-21, 0, -2.569961e-21, 1.28498e-20, -1.28498e-20, 
    5.139921e-21, -1.28498e-20, -1.541976e-20, 1.003089e-36, -7.709882e-21, 
    2.569961e-21, 1.027984e-20, 7.709882e-21, 5.139921e-21, 0, -2.569961e-21, 
    7.709882e-21, -1.003089e-36, -2.569961e-21, -5.139921e-21, 0, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, -1.003089e-36, 
    -1.027984e-20, 0, -1.003089e-36, 0, 5.139921e-21, -2.569961e-21, 
    1.798972e-20, 0, 7.709882e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    1.541976e-20, 2.569961e-21, 1.003089e-36, 0, 1.003089e-36, -7.709882e-21, 
    0, -1.28498e-20, 7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, 
    -1.003089e-36, 0, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -1.28498e-20, 2.569961e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, -7.709882e-21, 0, 5.139921e-21, 
    1.28498e-20, 1.027984e-20, -1.798972e-20, 5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, -2.569961e-21, 1.28498e-20, 1.027984e-20, -2.569961e-21, 
    1.003089e-36, 1.28498e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 0, 2.569961e-21, -1.28498e-20, 7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, -7.709882e-21, 
    7.709882e-21, 0, 0, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, 2.569961e-21, 1.027984e-20, 0, -7.709882e-21, 7.709882e-21, 
    -5.139921e-21, 7.709882e-21, 1.003089e-36, 2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 1.541976e-20, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, 1.027984e-20, 0, 0, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -1.003089e-36, -5.139921e-21, 1.003089e-36, -1.28498e-20, 
    5.139921e-21, 0, 0, -2.569961e-21, -1.541976e-20, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -1.003089e-36, -1.027984e-20, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 0, 7.709882e-21, -1.003089e-36, 1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    2.055969e-20, 1.003089e-36, -5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, -1.541976e-20, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, -1.798972e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -2.569961e-21, 1.28498e-20, 1.28498e-20, -7.709882e-21, 
    -2.569961e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 0, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    -7.709882e-21, 1.027984e-20, -1.003089e-36, 2.569961e-21, -1.798972e-20, 
    7.709882e-21, 7.709882e-21, 1.003089e-36, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 1.28498e-20, -5.139921e-21, -1.28498e-20, 
    -7.709882e-21, -5.139921e-21, 0, 1.798972e-20, 7.709882e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    0, -2.569961e-21, 0, 1.28498e-20, 1.28498e-20, 5.139921e-21, 
    -1.027984e-20, -2.569961e-21, 1.027984e-20, 1.027984e-20, 1.798972e-20, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, 1.027984e-20, 
    1.003089e-36, 7.709882e-21, 5.139921e-21, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, -1.003089e-36, 2.312965e-20, 2.312965e-20, 
    1.798972e-20, 5.139921e-21, 7.709882e-21, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.003089e-36, -5.139921e-21, -1.28498e-20, -1.28498e-20, 
    1.28498e-20, 7.709882e-21, -1.28498e-20, 5.139921e-21, 1.003089e-36, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -2.055969e-20, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, -2.569961e-21, 0, 2.569961e-21, 
    -1.28498e-20, 7.709882e-21, -1.541976e-20, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, -7.709882e-21, 
    7.709882e-21, 1.28498e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, -1.28498e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, 7.709882e-21, 1.027984e-20, 
    -1.28498e-20,
  -1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, -2.312965e-20, -7.709882e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 5.139921e-21, -2.055969e-20, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, 1.027984e-20, -1.28498e-20, -7.709882e-21, 
    -1.798972e-20, 1.28498e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, 1.003089e-36, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.569961e-21, -1.003089e-36, 2.569961e-21, 
    2.569961e-21, -1.003089e-36, 1.28498e-20, -1.003089e-36, -2.312965e-20, 
    -1.027984e-20, -7.709882e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, 
    -1.003089e-36, -5.139921e-21, 0, -2.569961e-21, 1.798972e-20, 
    -1.541976e-20, -1.28498e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, 1.798972e-20, 1.027984e-20, 1.003089e-36, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 0, 
    1.541976e-20, -2.569961e-21, -1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, 1.003089e-36, 2.569961e-21, 
    -1.003089e-36, -2.569961e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 7.709882e-21, -7.709882e-21, 
    -1.541976e-20, -2.055969e-20, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -1.541976e-20, 2.569961e-21, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    2.569961e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 0, -7.709882e-21, 
    -1.28498e-20, -7.709882e-21, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    1.798972e-20, 0, -5.139921e-21, 1.28498e-20, 1.28498e-20, 1.027984e-20, 
    0, -1.28498e-20, -2.569961e-21, -7.709882e-21, -1.28498e-20, 
    -1.28498e-20, -2.569961e-21, -1.28498e-20, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, -1.541976e-20, 
    1.027984e-20, -7.709882e-21, -1.541976e-20, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, 0, 5.139921e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, 
    0, 0, 5.139921e-21, -1.003089e-36, -1.28498e-20, -1.003089e-36, 
    -5.139921e-21, -2.055969e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, 1.28498e-20, 
    1.798972e-20, -1.541976e-20, 1.541976e-20, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -1.541976e-20, 1.003089e-36, -1.798972e-20, 
    -2.569961e-21, 5.139921e-21, 0, 1.003089e-36, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, 1.003089e-36, -2.569961e-21, 2.569961e-21, 
    2.055969e-20, 0, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, -2.055969e-20, 
    1.003089e-36, 1.541976e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, -1.027984e-20, 
    -1.541976e-20, 2.055969e-20, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -7.709882e-21, 1.28498e-20, -1.28498e-20, -1.28498e-20, 7.709882e-21, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, -1.28498e-20, 
    1.027984e-20, 2.569961e-21, -1.541976e-20, -5.139921e-21, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -1.541976e-20, -2.569961e-21, -1.798972e-20, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, -1.003089e-36, 1.027984e-20, 
    1.003089e-36, -7.709882e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    1.798972e-20, 5.139921e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 2.055969e-20, 7.709882e-21, 1.027984e-20, 
    2.569961e-21, 1.541976e-20, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.003089e-36, 0, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -1.003089e-36, 0, 1.027984e-20, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 1.541976e-20, -2.569961e-21, 7.709882e-21, -1.28498e-20, 
    -1.027984e-20, -7.709882e-21, -2.826957e-20, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 1.027984e-20, 1.28498e-20, 5.139921e-21, 
    1.541976e-20, -7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 7.709882e-21, 7.709882e-21, -5.139921e-21, 
    1.798972e-20, -1.798972e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -1.003089e-36,
  2.569961e-21, 5.139921e-21, -1.003089e-36, 1.541976e-20, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    1.541976e-20, 2.569961e-21, 1.28498e-20, 5.139921e-21, 1.027984e-20, 
    -1.28498e-20, -7.709882e-21, -3.083953e-20, -1.003089e-36, -1.003089e-36, 
    1.027984e-20, -2.569961e-21, 1.798972e-20, -2.569961e-21, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, -2.006177e-36, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, 7.709882e-21, -5.139921e-21, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 0, -1.28498e-20, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, 1.541976e-20, 7.709882e-21, -1.28498e-20, 1.003089e-36, 
    7.709882e-21, 0, 2.569961e-21, 5.139921e-21, 1.027984e-20, 2.055969e-20, 
    -7.709882e-21, 1.28498e-20, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -1.28498e-20, -1.798972e-20, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    0, 1.541976e-20, -1.798972e-20, -2.055969e-20, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -1.003089e-36, 0, 1.027984e-20, 
    1.003089e-36, 2.569961e-21, 2.569961e-21, 1.798972e-20, -2.055969e-20, 
    -7.709882e-21, -2.055969e-20, 7.709882e-21, -1.027984e-20, -5.139921e-21, 
    7.709882e-21, 1.28498e-20, -2.569961e-20, 2.055969e-20, 2.826957e-20, 
    -5.139921e-21, 1.027984e-20, 2.569961e-21, -1.541976e-20, 2.055969e-20, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, -1.28498e-20, 2.569961e-21, 
    -1.28498e-20, 2.569961e-21, -1.798972e-20, 7.709882e-21, 2.569961e-21, 
    2.055969e-20, 7.709882e-21, 1.003089e-36, -2.569961e-21, 1.798972e-20, 
    1.027984e-20, 1.027984e-20, -2.569961e-20, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, -1.798972e-20, -1.798972e-20, 
    -5.139921e-21, -1.027984e-20, -2.312965e-20, 1.541976e-20, 5.139921e-21, 
    1.798972e-20, 5.139921e-21, 1.541976e-20, 1.28498e-20, -2.569961e-21, 
    1.003089e-36, -5.139921e-21, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    -1.28498e-20, -1.28498e-20, -2.569961e-21, 2.312965e-20, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, 2.312965e-20, 1.541976e-20, 5.139921e-21, 
    1.003089e-36, 1.541976e-20, -1.027984e-20, -1.027984e-20, 7.709882e-21, 
    7.709882e-21, 1.003089e-36, -1.28498e-20, 2.569961e-21, -2.312965e-20, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 1.28498e-20, 7.709882e-21, 
    -1.027984e-20, 1.027984e-20, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    1.28498e-20, -1.027984e-20, 1.027984e-20, -1.003089e-36, 2.569961e-21, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, 1.28498e-20, 
    -1.798972e-20, 5.139921e-21, 0, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    0, 0, 2.569961e-21, 1.027984e-20, 5.139921e-21, 2.055969e-20, 
    -1.003089e-36, -2.055969e-20, -1.798972e-20, -5.139921e-21, 0, 
    -2.569961e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -1.541976e-20, -7.709882e-21, -3.083953e-20, 
    -1.798972e-20, -2.569961e-21, -1.28498e-20, -1.027984e-20, -2.569961e-21, 
    1.027984e-20, 0, 7.709882e-21, -1.027984e-20, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, 2.055969e-20, -7.709882e-21, 
    1.28498e-20, 1.541976e-20, -1.28498e-20, -1.28498e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.027984e-20, 1.28498e-20, -1.027984e-20, 
    1.28498e-20, 5.139921e-21, -1.027984e-20, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -1.003089e-36, -1.003089e-36, -7.709882e-21, -5.139921e-21, 
    -1.003089e-36, 1.541976e-20, -1.027984e-20, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 2.826957e-20, -5.139921e-21, 2.055969e-20, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -2.312965e-20, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 2.569961e-21, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, -2.569961e-21, 1.003089e-36, 7.709882e-21, 
    1.003089e-36, 2.569961e-21, -1.798972e-20, 1.027984e-20, -2.569961e-21, 
    1.027984e-20, 2.569961e-21, 1.027984e-20, 7.709882e-21, 1.798972e-20, 
    5.139921e-21, 2.569961e-21, 0, 7.709882e-21, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, 1.28498e-20, 
    5.139921e-21, -2.569961e-21, -1.541976e-20, 1.027984e-20, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, -1.28498e-20, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 5.139921e-21, 
    1.798972e-20, -5.139921e-21, 7.709882e-21, 5.139921e-21, 2.826957e-20, 
    2.569961e-21, 1.003089e-36, -1.28498e-20, -5.139921e-21, 1.28498e-20, 
    1.541976e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -2.569961e-21, 7.709882e-21, 1.28498e-20, -1.003089e-36, -7.709882e-21,
  6.259414e-29, 6.25942e-29, 6.259419e-29, 6.259424e-29, 6.259422e-29, 
    6.259425e-29, 6.259416e-29, 6.25942e-29, 6.259417e-29, 6.259414e-29, 
    6.259434e-29, 6.259425e-29, 6.259444e-29, 6.259438e-29, 6.259453e-29, 
    6.259443e-29, 6.259456e-29, 6.259453e-29, 6.259461e-29, 6.259459e-29, 
    6.259468e-29, 6.259462e-29, 6.259473e-29, 6.259466e-29, 6.259467e-29, 
    6.259461e-29, 6.259426e-29, 6.259433e-29, 6.259426e-29, 6.259427e-29, 
    6.259426e-29, 6.259422e-29, 6.259419e-29, 6.259414e-29, 6.259414e-29, 
    6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259432e-29, 6.259432e-29, 
    6.25944e-29, 6.259437e-29, 6.259451e-29, 6.259447e-29, 6.259459e-29, 
    6.259456e-29, 6.259458e-29, 6.259458e-29, 6.259458e-29, 6.259454e-29, 
    6.259456e-29, 6.259452e-29, 6.259437e-29, 6.259441e-29, 6.259429e-29, 
    6.259421e-29, 6.259416e-29, 6.259412e-29, 6.259413e-29, 6.259413e-29, 
    6.259419e-29, 6.259423e-29, 6.259427e-29, 6.259429e-29, 6.259432e-29, 
    6.259439e-29, 6.259443e-29, 6.259452e-29, 6.25945e-29, 6.259453e-29, 
    6.259455e-29, 6.259459e-29, 6.259459e-29, 6.259461e-29, 6.259453e-29, 
    6.259458e-29, 6.259449e-29, 6.259452e-29, 6.259432e-29, 6.259425e-29, 
    6.259422e-29, 6.259419e-29, 6.259413e-29, 6.259417e-29, 6.259416e-29, 
    6.25942e-29, 6.259423e-29, 6.259421e-29, 6.259429e-29, 6.259426e-29, 
    6.259443e-29, 6.259436e-29, 6.259455e-29, 6.25945e-29, 6.259456e-29, 
    6.259453e-29, 6.259458e-29, 6.259454e-29, 6.259461e-29, 6.259463e-29, 
    6.259462e-29, 6.259467e-29, 6.259453e-29, 6.259458e-29, 6.259421e-29, 
    6.259422e-29, 6.259422e-29, 6.259418e-29, 6.259417e-29, 6.259414e-29, 
    6.259417e-29, 6.259419e-29, 6.259423e-29, 6.259425e-29, 6.259427e-29, 
    6.259432e-29, 6.259438e-29, 6.259445e-29, 6.259451e-29, 6.259455e-29, 
    6.259452e-29, 6.259454e-29, 6.259452e-29, 6.259451e-29, 6.259463e-29, 
    6.259456e-29, 6.259466e-29, 6.259466e-29, 6.259461e-29, 6.259466e-29, 
    6.259422e-29, 6.25942e-29, 6.259416e-29, 6.259419e-29, 6.259413e-29, 
    6.259417e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 6.259429e-29, 
    6.259433e-29, 6.259437e-29, 6.259444e-29, 6.25945e-29, 6.259455e-29, 
    6.259455e-29, 6.259455e-29, 6.259456e-29, 6.259453e-29, 6.259457e-29, 
    6.259458e-29, 6.259456e-29, 6.259466e-29, 6.259463e-29, 6.259466e-29, 
    6.259464e-29, 6.259421e-29, 6.259423e-29, 6.259422e-29, 6.259424e-29, 
    6.259422e-29, 6.259429e-29, 6.259431e-29, 6.259441e-29, 6.259437e-29, 
    6.259443e-29, 6.259437e-29, 6.259438e-29, 6.259443e-29, 6.259438e-29, 
    6.25945e-29, 6.259441e-29, 6.259456e-29, 6.259449e-29, 6.259457e-29, 
    6.259455e-29, 6.259458e-29, 6.259461e-29, 6.259463e-29, 6.259469e-29, 
    6.259467e-29, 6.259472e-29, 6.259426e-29, 6.259429e-29, 6.259428e-29, 
    6.259431e-29, 6.259434e-29, 6.259438e-29, 6.259446e-29, 6.259443e-29, 
    6.259448e-29, 6.259449e-29, 6.259441e-29, 6.259446e-29, 6.259431e-29, 
    6.259433e-29, 6.259432e-29, 6.259426e-29, 6.259443e-29, 6.259435e-29, 
    6.259451e-29, 6.259446e-29, 6.25946e-29, 6.259453e-29, 6.259467e-29, 
    6.259473e-29, 6.259478e-29, 6.259485e-29, 6.25943e-29, 6.259428e-29, 
    6.259432e-29, 6.259437e-29, 6.259441e-29, 6.259446e-29, 6.259447e-29, 
    6.259448e-29, 6.259451e-29, 6.259453e-29, 6.259449e-29, 6.259454e-29, 
    6.259434e-29, 6.259444e-29, 6.259428e-29, 6.259432e-29, 6.259436e-29, 
    6.259435e-29, 6.259443e-29, 6.259444e-29, 6.259452e-29, 6.259448e-29, 
    6.259472e-29, 6.259461e-29, 6.25949e-29, 6.259482e-29, 6.259428e-29, 
    6.25943e-29, 6.259439e-29, 6.259435e-29, 6.259447e-29, 6.25945e-29, 
    6.259452e-29, 6.259455e-29, 6.259455e-29, 6.259457e-29, 6.259455e-29, 
    6.259457e-29, 6.259446e-29, 6.259451e-29, 6.259438e-29, 6.259441e-29, 
    6.25944e-29, 6.259438e-29, 6.259443e-29, 6.259449e-29, 6.259449e-29, 
    6.25945e-29, 6.259455e-29, 6.259447e-29, 6.259473e-29, 6.259456e-29, 
    6.259433e-29, 6.259438e-29, 6.259438e-29, 6.259437e-29, 6.259449e-29, 
    6.259445e-29, 6.259457e-29, 6.259454e-29, 6.259459e-29, 6.259456e-29, 
    6.259456e-29, 6.259453e-29, 6.25945e-29, 6.259445e-29, 6.25944e-29, 
    6.259437e-29, 6.259438e-29, 6.259441e-29, 6.259449e-29, 6.259455e-29, 
    6.259454e-29, 6.259459e-29, 6.259446e-29, 6.259452e-29, 6.259449e-29, 
    6.259455e-29, 6.259443e-29, 6.259453e-29, 6.25944e-29, 6.259441e-29, 
    6.259444e-29, 6.259452e-29, 6.259453e-29, 6.259455e-29, 6.259454e-29, 
    6.259449e-29, 6.259448e-29, 6.259444e-29, 6.259444e-29, 6.259441e-29, 
    6.259438e-29, 6.259441e-29, 6.259443e-29, 6.259449e-29, 6.259455e-29, 
    6.259461e-29, 6.259462e-29, 6.259469e-29, 6.259463e-29, 6.259473e-29, 
    6.259465e-29, 6.259479e-29, 6.259453e-29, 6.259464e-29, 6.259445e-29, 
    6.259447e-29, 6.259451e-29, 6.259459e-29, 6.259455e-29, 6.25946e-29, 
    6.259448e-29, 6.259442e-29, 6.25944e-29, 6.259437e-29, 6.25944e-29, 
    6.25944e-29, 6.259443e-29, 6.259442e-29, 6.259449e-29, 6.259446e-29, 
    6.259456e-29, 6.25946e-29, 6.259472e-29, 6.259479e-29, 6.259485e-29, 
    6.259489e-29, 6.25949e-29, 6.25949e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.19423e-10, 2.203886e-10, 2.202009e-10, 2.209797e-10, 2.205476e-10, 
    2.210576e-10, 2.196188e-10, 2.204269e-10, 2.19911e-10, 2.195099e-10, 
    2.22491e-10, 2.210144e-10, 2.240248e-10, 2.23083e-10, 2.254486e-10, 
    2.238782e-10, 2.257653e-10, 2.254033e-10, 2.264927e-10, 2.261806e-10, 
    2.275741e-10, 2.266368e-10, 2.282964e-10, 2.273502e-10, 2.274983e-10, 
    2.266058e-10, 2.213115e-10, 2.223072e-10, 2.212525e-10, 2.213945e-10, 
    2.213308e-10, 2.205566e-10, 2.201664e-10, 2.193492e-10, 2.194975e-10, 
    2.200978e-10, 2.214584e-10, 2.209965e-10, 2.221605e-10, 2.221342e-10, 
    2.234301e-10, 2.228458e-10, 2.250238e-10, 2.244048e-10, 2.261936e-10, 
    2.257438e-10, 2.261725e-10, 2.260425e-10, 2.261742e-10, 2.255144e-10, 
    2.257971e-10, 2.252165e-10, 2.229552e-10, 2.236198e-10, 2.216377e-10, 
    2.204459e-10, 2.196542e-10, 2.190924e-10, 2.191719e-10, 2.193233e-10, 
    2.201013e-10, 2.208327e-10, 2.213902e-10, 2.21763e-10, 2.221304e-10, 
    2.232426e-10, 2.238311e-10, 2.25149e-10, 2.249112e-10, 2.253141e-10, 
    2.25699e-10, 2.263453e-10, 2.262389e-10, 2.265236e-10, 2.253035e-10, 
    2.261144e-10, 2.247757e-10, 2.251418e-10, 2.222304e-10, 2.211211e-10, 
    2.206497e-10, 2.202369e-10, 2.192329e-10, 2.199263e-10, 2.19653e-10, 
    2.203032e-10, 2.207164e-10, 2.20512e-10, 2.217732e-10, 2.212829e-10, 
    2.23866e-10, 2.227534e-10, 2.256541e-10, 2.2496e-10, 2.258205e-10, 
    2.253814e-10, 2.261338e-10, 2.254566e-10, 2.266296e-10, 2.26885e-10, 
    2.267105e-10, 2.273809e-10, 2.254191e-10, 2.261725e-10, 2.205063e-10, 
    2.205396e-10, 2.206949e-10, 2.200124e-10, 2.199706e-10, 2.193451e-10, 
    2.199017e-10, 2.201387e-10, 2.207403e-10, 2.210962e-10, 2.214345e-10, 
    2.221783e-10, 2.23009e-10, 2.241705e-10, 2.25005e-10, 2.255644e-10, 
    2.252214e-10, 2.255242e-10, 2.251857e-10, 2.25027e-10, 2.267893e-10, 
    2.257998e-10, 2.272845e-10, 2.272023e-10, 2.265304e-10, 2.272116e-10, 
    2.20563e-10, 2.203712e-10, 2.197054e-10, 2.202265e-10, 2.19277e-10, 
    2.198085e-10, 2.201141e-10, 2.212932e-10, 2.215522e-10, 2.217924e-10, 
    2.222669e-10, 2.228757e-10, 2.239438e-10, 2.248731e-10, 2.257214e-10, 
    2.256593e-10, 2.256811e-10, 2.258707e-10, 2.254012e-10, 2.259477e-10, 
    2.260395e-10, 2.257996e-10, 2.271913e-10, 2.267937e-10, 2.272006e-10, 
    2.269417e-10, 2.204336e-10, 2.207563e-10, 2.205819e-10, 2.209098e-10, 
    2.206788e-10, 2.217061e-10, 2.220141e-10, 2.234552e-10, 2.228637e-10, 
    2.23805e-10, 2.229593e-10, 2.231092e-10, 2.238358e-10, 2.23005e-10, 
    2.248219e-10, 2.235901e-10, 2.25878e-10, 2.246481e-10, 2.259551e-10, 
    2.257177e-10, 2.261107e-10, 2.264627e-10, 2.269055e-10, 2.277225e-10, 
    2.275333e-10, 2.282165e-10, 2.212374e-10, 2.21656e-10, 2.216191e-10, 
    2.220572e-10, 2.223811e-10, 2.230833e-10, 2.242094e-10, 2.237859e-10, 
    2.245634e-10, 2.247195e-10, 2.235383e-10, 2.242635e-10, 2.219361e-10, 
    2.223122e-10, 2.220883e-10, 2.212704e-10, 2.238836e-10, 2.225425e-10, 
    2.250188e-10, 2.242923e-10, 2.264125e-10, 2.253581e-10, 2.274291e-10, 
    2.283145e-10, 2.291477e-10, 2.301215e-10, 2.218844e-10, 2.216e-10, 
    2.221092e-10, 2.228139e-10, 2.234676e-10, 2.243366e-10, 2.244255e-10, 
    2.245884e-10, 2.250101e-10, 2.253647e-10, 2.246399e-10, 2.254536e-10, 
    2.223994e-10, 2.239999e-10, 2.214925e-10, 2.222476e-10, 2.227723e-10, 
    2.225421e-10, 2.237375e-10, 2.240193e-10, 2.251642e-10, 2.245723e-10, 
    2.28096e-10, 2.265371e-10, 2.308629e-10, 2.29654e-10, 2.215006e-10, 
    2.218834e-10, 2.232157e-10, 2.225818e-10, 2.243946e-10, 2.248409e-10, 
    2.252036e-10, 2.256673e-10, 2.257174e-10, 2.259921e-10, 2.255419e-10, 
    2.259743e-10, 2.243385e-10, 2.250695e-10, 2.230634e-10, 2.235517e-10, 
    2.233271e-10, 2.230807e-10, 2.238411e-10, 2.246513e-10, 2.246686e-10, 
    2.249283e-10, 2.256604e-10, 2.24402e-10, 2.282973e-10, 2.258917e-10, 
    2.223009e-10, 2.230382e-10, 2.231435e-10, 2.228579e-10, 2.247961e-10, 
    2.240938e-10, 2.259854e-10, 2.254742e-10, 2.263118e-10, 2.258956e-10, 
    2.258343e-10, 2.252997e-10, 2.249669e-10, 2.241261e-10, 2.234419e-10, 
    2.228993e-10, 2.230255e-10, 2.236215e-10, 2.247008e-10, 2.257219e-10, 
    2.254982e-10, 2.262481e-10, 2.242632e-10, 2.250955e-10, 2.247739e-10, 
    2.256126e-10, 2.237747e-10, 2.253399e-10, 2.233746e-10, 2.235469e-10, 
    2.240799e-10, 2.25152e-10, 2.253892e-10, 2.256424e-10, 2.254861e-10, 
    2.247282e-10, 2.24604e-10, 2.240669e-10, 2.239187e-10, 2.235094e-10, 
    2.231706e-10, 2.234802e-10, 2.238053e-10, 2.247285e-10, 2.255606e-10, 
    2.264677e-10, 2.266897e-10, 2.277497e-10, 2.268868e-10, 2.283107e-10, 
    2.271002e-10, 2.291956e-10, 2.254305e-10, 2.270645e-10, 2.241041e-10, 
    2.244231e-10, 2.249999e-10, 2.26323e-10, 2.256087e-10, 2.26444e-10, 
    2.245992e-10, 2.23642e-10, 2.233943e-10, 2.229323e-10, 2.234049e-10, 
    2.233665e-10, 2.238187e-10, 2.236734e-10, 2.247592e-10, 2.241759e-10, 
    2.258328e-10, 2.264375e-10, 2.281449e-10, 2.291917e-10, 2.302572e-10, 
    2.307276e-10, 2.308707e-10, 2.309306e-10 ;

 SOIL2N_TO_SOIL3N =
  1.567307e-11, 1.574204e-11, 1.572863e-11, 1.578426e-11, 1.57534e-11, 
    1.578983e-11, 1.568705e-11, 1.574478e-11, 1.570793e-11, 1.567928e-11, 
    1.589222e-11, 1.578674e-11, 1.600177e-11, 1.59345e-11, 1.610347e-11, 
    1.59913e-11, 1.612609e-11, 1.610024e-11, 1.617805e-11, 1.615576e-11, 
    1.625529e-11, 1.618834e-11, 1.630688e-11, 1.62393e-11, 1.624987e-11, 
    1.618613e-11, 1.580797e-11, 1.587909e-11, 1.580375e-11, 1.58139e-11, 
    1.580934e-11, 1.575404e-11, 1.572617e-11, 1.56678e-11, 1.56784e-11, 
    1.572127e-11, 1.581846e-11, 1.578546e-11, 1.586861e-11, 1.586673e-11, 
    1.595929e-11, 1.591756e-11, 1.607313e-11, 1.602892e-11, 1.615669e-11, 
    1.612455e-11, 1.615518e-11, 1.614589e-11, 1.61553e-11, 1.610817e-11, 
    1.612837e-11, 1.60869e-11, 1.592537e-11, 1.597284e-11, 1.583127e-11, 
    1.574614e-11, 1.568959e-11, 1.564946e-11, 1.565513e-11, 1.566595e-11, 
    1.572152e-11, 1.577377e-11, 1.581358e-11, 1.584022e-11, 1.586646e-11, 
    1.59459e-11, 1.598794e-11, 1.608207e-11, 1.606508e-11, 1.609387e-11, 
    1.612136e-11, 1.616752e-11, 1.615992e-11, 1.618026e-11, 1.60931e-11, 
    1.615103e-11, 1.605541e-11, 1.608156e-11, 1.58736e-11, 1.579436e-11, 
    1.576069e-11, 1.573121e-11, 1.565949e-11, 1.570902e-11, 1.56895e-11, 
    1.573594e-11, 1.576546e-11, 1.575086e-11, 1.584094e-11, 1.580592e-11, 
    1.599043e-11, 1.591096e-11, 1.611815e-11, 1.606857e-11, 1.613003e-11, 
    1.609867e-11, 1.615241e-11, 1.610405e-11, 1.618783e-11, 1.620607e-11, 
    1.619361e-11, 1.624149e-11, 1.610137e-11, 1.615518e-11, 1.575045e-11, 
    1.575283e-11, 1.576392e-11, 1.571517e-11, 1.571219e-11, 1.566751e-11, 
    1.570726e-11, 1.572419e-11, 1.576717e-11, 1.579259e-11, 1.581675e-11, 
    1.586988e-11, 1.592921e-11, 1.601218e-11, 1.607178e-11, 1.611174e-11, 
    1.608724e-11, 1.610887e-11, 1.608469e-11, 1.607336e-11, 1.619924e-11, 
    1.612855e-11, 1.623461e-11, 1.622874e-11, 1.618074e-11, 1.62294e-11, 
    1.57545e-11, 1.57408e-11, 1.569324e-11, 1.573046e-11, 1.566264e-11, 
    1.570061e-11, 1.572243e-11, 1.580666e-11, 1.582516e-11, 1.584232e-11, 
    1.58762e-11, 1.591969e-11, 1.599599e-11, 1.606236e-11, 1.612296e-11, 
    1.611852e-11, 1.612008e-11, 1.613362e-11, 1.610009e-11, 1.613912e-11, 
    1.614568e-11, 1.612854e-11, 1.622795e-11, 1.619955e-11, 1.622861e-11, 
    1.621012e-11, 1.574526e-11, 1.576831e-11, 1.575585e-11, 1.577927e-11, 
    1.576277e-11, 1.583615e-11, 1.585815e-11, 1.596108e-11, 1.591884e-11, 
    1.598607e-11, 1.592567e-11, 1.593637e-11, 1.598827e-11, 1.592893e-11, 
    1.60587e-11, 1.597072e-11, 1.613414e-11, 1.604629e-11, 1.613965e-11, 
    1.61227e-11, 1.615077e-11, 1.617591e-11, 1.620753e-11, 1.626589e-11, 
    1.625238e-11, 1.630118e-11, 1.580267e-11, 1.583257e-11, 1.582994e-11, 
    1.586123e-11, 1.588437e-11, 1.593452e-11, 1.601496e-11, 1.598471e-11, 
    1.604024e-11, 1.605139e-11, 1.596702e-11, 1.601882e-11, 1.585258e-11, 
    1.587944e-11, 1.586345e-11, 1.580503e-11, 1.599168e-11, 1.589589e-11, 
    1.607277e-11, 1.602088e-11, 1.617232e-11, 1.609701e-11, 1.624494e-11, 
    1.630818e-11, 1.63677e-11, 1.643725e-11, 1.584889e-11, 1.582857e-11, 
    1.586495e-11, 1.591527e-11, 1.596197e-11, 1.602404e-11, 1.60304e-11, 
    1.604203e-11, 1.607215e-11, 1.609748e-11, 1.60457e-11, 1.610382e-11, 
    1.588567e-11, 1.6e-11, 1.582089e-11, 1.587483e-11, 1.591231e-11, 
    1.589586e-11, 1.598125e-11, 1.600138e-11, 1.608316e-11, 1.604088e-11, 
    1.629257e-11, 1.618122e-11, 1.649021e-11, 1.640386e-11, 1.582147e-11, 
    1.584882e-11, 1.594398e-11, 1.58987e-11, 1.602819e-11, 1.606006e-11, 
    1.608597e-11, 1.611909e-11, 1.612267e-11, 1.614229e-11, 1.611013e-11, 
    1.614102e-11, 1.602418e-11, 1.607639e-11, 1.59331e-11, 1.596798e-11, 
    1.595193e-11, 1.593434e-11, 1.598865e-11, 1.604652e-11, 1.604775e-11, 
    1.606631e-11, 1.61186e-11, 1.602871e-11, 1.630695e-11, 1.613512e-11, 
    1.587863e-11, 1.59313e-11, 1.593882e-11, 1.591842e-11, 1.605687e-11, 
    1.60067e-11, 1.614181e-11, 1.61053e-11, 1.616513e-11, 1.61354e-11, 
    1.613102e-11, 1.609284e-11, 1.606906e-11, 1.6009e-11, 1.596013e-11, 
    1.592138e-11, 1.593039e-11, 1.597296e-11, 1.605006e-11, 1.612299e-11, 
    1.610702e-11, 1.616058e-11, 1.60188e-11, 1.607825e-11, 1.605528e-11, 
    1.611519e-11, 1.598391e-11, 1.609571e-11, 1.595533e-11, 1.596764e-11, 
    1.600571e-11, 1.608229e-11, 1.609923e-11, 1.611732e-11, 1.610615e-11, 
    1.605202e-11, 1.604315e-11, 1.600478e-11, 1.599419e-11, 1.596496e-11, 
    1.594076e-11, 1.596287e-11, 1.598609e-11, 1.605204e-11, 1.611147e-11, 
    1.617627e-11, 1.619212e-11, 1.626783e-11, 1.62062e-11, 1.630791e-11, 
    1.622144e-11, 1.637111e-11, 1.610218e-11, 1.62189e-11, 1.600744e-11, 
    1.603022e-11, 1.607143e-11, 1.616593e-11, 1.611491e-11, 1.617458e-11, 
    1.60428e-11, 1.597443e-11, 1.595674e-11, 1.592374e-11, 1.595749e-11, 
    1.595475e-11, 1.598705e-11, 1.597667e-11, 1.605423e-11, 1.601257e-11, 
    1.613091e-11, 1.61741e-11, 1.629607e-11, 1.637084e-11, 1.644694e-11, 
    1.648054e-11, 1.649077e-11, 1.649504e-11 ;

 SOIL2N_vr =
  1.818769, 1.818771, 1.81877, 1.818772, 1.818771, 1.818772, 1.81877, 
    1.818771, 1.81877, 1.818769, 1.818774, 1.818772, 1.818776, 1.818775, 
    1.818779, 1.818776, 1.818779, 1.818779, 1.81878, 1.81878, 1.818782, 
    1.818781, 1.818783, 1.818782, 1.818782, 1.818781, 1.818772, 1.818774, 
    1.818772, 1.818772, 1.818772, 1.818771, 1.81877, 1.818769, 1.818769, 
    1.81877, 1.818772, 1.818772, 1.818774, 1.818774, 1.818776, 1.818775, 
    1.818778, 1.818777, 1.81878, 1.818779, 1.81878, 1.81878, 1.81878, 
    1.818779, 1.818779, 1.818778, 1.818775, 1.818776, 1.818773, 1.818771, 
    1.81877, 1.818769, 1.818769, 1.818769, 1.81877, 1.818771, 1.818772, 
    1.818773, 1.818774, 1.818775, 1.818776, 1.818778, 1.818778, 1.818779, 
    1.818779, 1.81878, 1.81878, 1.81878, 1.818779, 1.81878, 1.818778, 
    1.818778, 1.818774, 1.818772, 1.818771, 1.818771, 1.818769, 1.81877, 
    1.81877, 1.818771, 1.818771, 1.818771, 1.818773, 1.818772, 1.818776, 
    1.818774, 1.818779, 1.818778, 1.818779, 1.818779, 1.81878, 1.818779, 
    1.818781, 1.818781, 1.818781, 1.818782, 1.818779, 1.81878, 1.818771, 
    1.818771, 1.818771, 1.81877, 1.81877, 1.818769, 1.81877, 1.81877, 
    1.818771, 1.818772, 1.818772, 1.818774, 1.818775, 1.818777, 1.818778, 
    1.818779, 1.818778, 1.818779, 1.818778, 1.818778, 1.818781, 1.818779, 
    1.818782, 1.818781, 1.81878, 1.818781, 1.818771, 1.818771, 1.81877, 
    1.818771, 1.818769, 1.81877, 1.81877, 1.818772, 1.818773, 1.818773, 
    1.818774, 1.818775, 1.818776, 1.818778, 1.818779, 1.818779, 1.818779, 
    1.818779, 1.818779, 1.81878, 1.81878, 1.818779, 1.818781, 1.818781, 
    1.818781, 1.818781, 1.818771, 1.818771, 1.818771, 1.818772, 1.818771, 
    1.818773, 1.818773, 1.818776, 1.818775, 1.818776, 1.818775, 1.818775, 
    1.818776, 1.818775, 1.818778, 1.818776, 1.818779, 1.818777, 1.81878, 
    1.818779, 1.81878, 1.81878, 1.818781, 1.818782, 1.818782, 1.818783, 
    1.818772, 1.818773, 1.818773, 1.818773, 1.818774, 1.818775, 1.818777, 
    1.818776, 1.818777, 1.818778, 1.818776, 1.818777, 1.818773, 1.818774, 
    1.818773, 1.818772, 1.818776, 1.818774, 1.818778, 1.818777, 1.81878, 
    1.818779, 1.818782, 1.818783, 1.818785, 1.818786, 1.818773, 1.818773, 
    1.818774, 1.818775, 1.818776, 1.818777, 1.818777, 1.818777, 1.818778, 
    1.818779, 1.818777, 1.818779, 1.818774, 1.818776, 1.818773, 1.818774, 
    1.818775, 1.818774, 1.818776, 1.818776, 1.818778, 1.818777, 1.818783, 
    1.81878, 1.818787, 1.818785, 1.818773, 1.818773, 1.818775, 1.818774, 
    1.818777, 1.818778, 1.818778, 1.818779, 1.818779, 1.81878, 1.818779, 
    1.81878, 1.818777, 1.818778, 1.818775, 1.818776, 1.818775, 1.818775, 
    1.818776, 1.818777, 1.818778, 1.818778, 1.818779, 1.818777, 1.818783, 
    1.818779, 1.818774, 1.818775, 1.818775, 1.818775, 1.818778, 1.818777, 
    1.81878, 1.818779, 1.81878, 1.818779, 1.818779, 1.818779, 1.818778, 
    1.818777, 1.818776, 1.818775, 1.818775, 1.818776, 1.818778, 1.818779, 
    1.818779, 1.81878, 1.818777, 1.818778, 1.818778, 1.818779, 1.818776, 
    1.818779, 1.818776, 1.818776, 1.818777, 1.818778, 1.818779, 1.818779, 
    1.818779, 1.818778, 1.818777, 1.818777, 1.818776, 1.818776, 1.818775, 
    1.818776, 1.818776, 1.818778, 1.818779, 1.81878, 1.818781, 1.818782, 
    1.818781, 1.818783, 1.818781, 1.818785, 1.818779, 1.818781, 1.818777, 
    1.818777, 1.818778, 1.81878, 1.818779, 1.81878, 1.818777, 1.818776, 
    1.818776, 1.818775, 1.818776, 1.818775, 1.818776, 1.818776, 1.818778, 
    1.818777, 1.818779, 1.81878, 1.818783, 1.818785, 1.818786, 1.818787, 
    1.818787, 1.818787,
  1.818734, 1.818736, 1.818735, 1.818737, 1.818736, 1.818737, 1.818734, 
    1.818736, 1.818735, 1.818734, 1.81874, 1.818737, 1.818743, 1.818741, 
    1.818746, 1.818743, 1.818747, 1.818746, 1.818749, 1.818748, 1.818751, 
    1.818749, 1.818753, 1.818751, 1.818751, 1.818749, 1.818738, 1.81874, 
    1.818738, 1.818738, 1.818738, 1.818736, 1.818735, 1.818733, 1.818734, 
    1.818735, 1.818738, 1.818737, 1.818739, 1.818739, 1.818742, 1.818741, 
    1.818745, 1.818744, 1.818748, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818747, 1.818746, 1.818741, 1.818743, 1.818738, 1.818736, 
    1.818734, 1.818733, 1.818733, 1.818733, 1.818735, 1.818737, 1.818738, 
    1.818739, 1.818739, 1.818742, 1.818743, 1.818746, 1.818745, 1.818746, 
    1.818747, 1.818748, 1.818748, 1.818749, 1.818746, 1.818748, 1.818745, 
    1.818746, 1.81874, 1.818737, 1.818736, 1.818735, 1.818733, 1.818735, 
    1.818734, 1.818735, 1.818736, 1.818736, 1.818739, 1.818738, 1.818743, 
    1.818741, 1.818747, 1.818745, 1.818747, 1.818746, 1.818748, 1.818746, 
    1.818749, 1.81875, 1.818749, 1.818751, 1.818746, 1.818748, 1.818736, 
    1.818736, 1.818736, 1.818735, 1.818735, 1.818733, 1.818735, 1.818735, 
    1.818736, 1.818737, 1.818738, 1.81874, 1.818741, 1.818744, 1.818745, 
    1.818747, 1.818746, 1.818747, 1.818746, 1.818746, 1.818749, 1.818747, 
    1.81875, 1.81875, 1.818749, 1.81875, 1.818736, 1.818736, 1.818734, 
    1.818735, 1.818733, 1.818734, 1.818735, 1.818738, 1.818738, 1.818739, 
    1.81874, 1.818741, 1.818743, 1.818745, 1.818747, 1.818747, 1.818747, 
    1.818747, 1.818746, 1.818748, 1.818748, 1.818747, 1.81875, 1.818749, 
    1.81875, 1.81875, 1.818736, 1.818736, 1.818736, 1.818737, 1.818736, 
    1.818738, 1.818739, 1.818742, 1.818741, 1.818743, 1.818741, 1.818741, 
    1.818743, 1.818741, 1.818745, 1.818743, 1.818747, 1.818745, 1.818748, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818751, 1.818751, 1.818752, 
    1.818738, 1.818738, 1.818738, 1.818739, 1.81874, 1.818741, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818742, 1.818744, 1.818739, 1.81874, 
    1.818739, 1.818738, 1.818743, 1.81874, 1.818745, 1.818744, 1.818748, 
    1.818746, 1.818751, 1.818753, 1.818754, 1.818756, 1.818739, 1.818738, 
    1.818739, 1.818741, 1.818742, 1.818744, 1.818744, 1.818745, 1.818745, 
    1.818746, 1.818745, 1.818746, 1.81874, 1.818743, 1.818738, 1.81874, 
    1.818741, 1.81874, 1.818743, 1.818743, 1.818746, 1.818745, 1.818752, 
    1.818749, 1.818758, 1.818755, 1.818738, 1.818739, 1.818742, 1.81874, 
    1.818744, 1.818745, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 
    1.818748, 1.818744, 1.818746, 1.818741, 1.818742, 1.818742, 1.818741, 
    1.818743, 1.818745, 1.818745, 1.818745, 1.818747, 1.818744, 1.818753, 
    1.818747, 1.81874, 1.818741, 1.818742, 1.818741, 1.818745, 1.818744, 
    1.818748, 1.818747, 1.818748, 1.818747, 1.818747, 1.818746, 1.818745, 
    1.818744, 1.818742, 1.818741, 1.818741, 1.818743, 1.818745, 1.818747, 
    1.818747, 1.818748, 1.818744, 1.818746, 1.818745, 1.818747, 1.818743, 
    1.818746, 1.818742, 1.818742, 1.818744, 1.818746, 1.818746, 1.818747, 
    1.818747, 1.818745, 1.818745, 1.818743, 1.818743, 1.818742, 1.818742, 
    1.818742, 1.818743, 1.818745, 1.818747, 1.818749, 1.818749, 1.818751, 
    1.81875, 1.818753, 1.81875, 1.818754, 1.818746, 1.81875, 1.818744, 
    1.818744, 1.818745, 1.818748, 1.818747, 1.818749, 1.818745, 1.818743, 
    1.818742, 1.818741, 1.818742, 1.818742, 1.818743, 1.818743, 1.818745, 
    1.818744, 1.818747, 1.818749, 1.818752, 1.818754, 1.818757, 1.818758, 
    1.818758, 1.818758,
  1.818684, 1.818686, 1.818685, 1.818687, 1.818686, 1.818687, 1.818684, 
    1.818686, 1.818685, 1.818684, 1.818691, 1.818687, 1.818694, 1.818692, 
    1.818697, 1.818694, 1.818698, 1.818697, 1.8187, 1.818699, 1.818702, 
    1.8187, 1.818704, 1.818702, 1.818702, 1.8187, 1.818688, 1.81869, 
    1.818688, 1.818688, 1.818688, 1.818686, 1.818685, 1.818683, 1.818684, 
    1.818685, 1.818688, 1.818687, 1.81869, 1.81869, 1.818693, 1.818691, 
    1.818696, 1.818695, 1.818699, 1.818698, 1.818699, 1.818699, 1.818699, 
    1.818697, 1.818698, 1.818697, 1.818692, 1.818693, 1.818689, 1.818686, 
    1.818684, 1.818683, 1.818683, 1.818683, 1.818685, 1.818687, 1.818688, 
    1.818689, 1.81869, 1.818692, 1.818694, 1.818697, 1.818696, 1.818697, 
    1.818698, 1.818699, 1.818699, 1.8187, 1.818697, 1.818699, 1.818696, 
    1.818697, 1.81869, 1.818687, 1.818686, 1.818685, 1.818683, 1.818685, 
    1.818684, 1.818686, 1.818686, 1.818686, 1.818689, 1.818688, 1.818694, 
    1.818691, 1.818698, 1.818696, 1.818698, 1.818697, 1.818699, 1.818697, 
    1.8187, 1.818701, 1.8187, 1.818702, 1.818697, 1.818699, 1.818686, 
    1.818686, 1.818686, 1.818685, 1.818685, 1.818683, 1.818685, 1.818685, 
    1.818687, 1.818687, 1.818688, 1.81869, 1.818692, 1.818694, 1.818696, 
    1.818698, 1.818697, 1.818697, 1.818697, 1.818696, 1.8187, 1.818698, 
    1.818702, 1.818701, 1.8187, 1.818701, 1.818686, 1.818686, 1.818684, 
    1.818685, 1.818683, 1.818684, 1.818685, 1.818688, 1.818688, 1.818689, 
    1.81869, 1.818691, 1.818694, 1.818696, 1.818698, 1.818698, 1.818698, 
    1.818698, 1.818697, 1.818698, 1.818699, 1.818698, 1.818701, 1.8187, 
    1.818701, 1.818701, 1.818686, 1.818687, 1.818686, 1.818687, 1.818686, 
    1.818689, 1.818689, 1.818693, 1.818691, 1.818694, 1.818692, 1.818692, 
    1.818694, 1.818692, 1.818696, 1.818693, 1.818698, 1.818695, 1.818698, 
    1.818698, 1.818699, 1.8187, 1.818701, 1.818702, 1.818702, 1.818704, 
    1.818688, 1.818689, 1.818689, 1.81869, 1.81869, 1.818692, 1.818694, 
    1.818694, 1.818695, 1.818696, 1.818693, 1.818695, 1.818689, 1.81869, 
    1.81869, 1.818688, 1.818694, 1.818691, 1.818696, 1.818695, 1.818699, 
    1.818697, 1.818702, 1.818704, 1.818706, 1.818708, 1.818689, 1.818689, 
    1.81869, 1.818691, 1.818693, 1.818695, 1.818695, 1.818695, 1.818696, 
    1.818697, 1.818695, 1.818697, 1.81869, 1.818694, 1.818688, 1.81869, 
    1.818691, 1.818691, 1.818693, 1.818694, 1.818697, 1.818695, 1.818703, 
    1.8187, 1.818709, 1.818707, 1.818688, 1.818689, 1.818692, 1.818691, 
    1.818695, 1.818696, 1.818697, 1.818698, 1.818698, 1.818699, 1.818697, 
    1.818699, 1.818695, 1.818696, 1.818692, 1.818693, 1.818692, 1.818692, 
    1.818694, 1.818695, 1.818696, 1.818696, 1.818698, 1.818695, 1.818704, 
    1.818698, 1.81869, 1.818692, 1.818692, 1.818691, 1.818696, 1.818694, 
    1.818699, 1.818697, 1.818699, 1.818698, 1.818698, 1.818697, 1.818696, 
    1.818694, 1.818693, 1.818691, 1.818692, 1.818693, 1.818696, 1.818698, 
    1.818697, 1.818699, 1.818695, 1.818696, 1.818696, 1.818698, 1.818694, 
    1.818697, 1.818693, 1.818693, 1.818694, 1.818697, 1.818697, 1.818698, 
    1.818697, 1.818696, 1.818695, 1.818694, 1.818694, 1.818693, 1.818692, 
    1.818693, 1.818694, 1.818696, 1.818698, 1.8187, 1.8187, 1.818702, 
    1.818701, 1.818704, 1.818701, 1.818706, 1.818697, 1.818701, 1.818694, 
    1.818695, 1.818696, 1.818699, 1.818698, 1.8187, 1.818695, 1.818693, 
    1.818693, 1.818692, 1.818693, 1.818693, 1.818694, 1.818693, 1.818696, 
    1.818694, 1.818698, 1.818699, 1.818703, 1.818706, 1.818708, 1.818709, 
    1.81871, 1.81871,
  1.818644, 1.818646, 1.818645, 1.818647, 1.818646, 1.818647, 1.818644, 
    1.818646, 1.818645, 1.818644, 1.818651, 1.818647, 1.818654, 1.818652, 
    1.818657, 1.818654, 1.818658, 1.818657, 1.81866, 1.818659, 1.818662, 
    1.81866, 1.818664, 1.818662, 1.818662, 1.81866, 1.818648, 1.81865, 
    1.818648, 1.818648, 1.818648, 1.818646, 1.818645, 1.818643, 1.818644, 
    1.818645, 1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 
    1.818656, 1.818655, 1.818659, 1.818658, 1.818659, 1.818659, 1.818659, 
    1.818657, 1.818658, 1.818657, 1.818652, 1.818653, 1.818649, 1.818646, 
    1.818644, 1.818643, 1.818643, 1.818643, 1.818645, 1.818647, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818654, 1.818657, 1.818656, 1.818657, 
    1.818658, 1.818659, 1.818659, 1.81866, 1.818657, 1.818659, 1.818656, 
    1.818657, 1.81865, 1.818648, 1.818646, 1.818645, 1.818643, 1.818645, 
    1.818644, 1.818646, 1.818647, 1.818646, 1.818649, 1.818648, 1.818654, 
    1.818651, 1.818658, 1.818656, 1.818658, 1.818657, 1.818659, 1.818657, 
    1.81866, 1.81866, 1.81866, 1.818662, 1.818657, 1.818659, 1.818646, 
    1.818646, 1.818647, 1.818645, 1.818645, 1.818643, 1.818645, 1.818645, 
    1.818647, 1.818647, 1.818648, 1.81865, 1.818652, 1.818654, 1.818656, 
    1.818658, 1.818657, 1.818657, 1.818657, 1.818656, 1.81866, 1.818658, 
    1.818661, 1.818661, 1.81866, 1.818661, 1.818646, 1.818646, 1.818644, 
    1.818645, 1.818643, 1.818645, 1.818645, 1.818648, 1.818648, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818656, 1.818658, 1.818658, 1.818658, 
    1.818658, 1.818657, 1.818658, 1.818659, 1.818658, 1.818661, 1.81866, 
    1.818661, 1.818661, 1.818646, 1.818647, 1.818646, 1.818647, 1.818646, 
    1.818649, 1.81865, 1.818653, 1.818651, 1.818654, 1.818652, 1.818652, 
    1.818654, 1.818652, 1.818656, 1.818653, 1.818658, 1.818655, 1.818658, 
    1.818658, 1.818659, 1.81866, 1.81866, 1.818662, 1.818662, 1.818663, 
    1.818648, 1.818649, 1.818649, 1.81865, 1.81865, 1.818652, 1.818654, 
    1.818653, 1.818655, 1.818656, 1.818653, 1.818655, 1.818649, 1.81865, 
    1.81865, 1.818648, 1.818654, 1.818651, 1.818656, 1.818655, 1.818659, 
    1.818657, 1.818662, 1.818664, 1.818666, 1.818668, 1.818649, 1.818649, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 1.818656, 
    1.818657, 1.818655, 1.818657, 1.81865, 1.818654, 1.818648, 1.81865, 
    1.818651, 1.818651, 1.818653, 1.818654, 1.818657, 1.818655, 1.818663, 
    1.81866, 1.818669, 1.818667, 1.818648, 1.818649, 1.818652, 1.818651, 
    1.818655, 1.818656, 1.818657, 1.818658, 1.818658, 1.818658, 1.818657, 
    1.818658, 1.818655, 1.818656, 1.818652, 1.818653, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818655, 1.818656, 1.818658, 1.818655, 1.818664, 
    1.818658, 1.81865, 1.818652, 1.818652, 1.818651, 1.818656, 1.818654, 
    1.818658, 1.818657, 1.818659, 1.818658, 1.818658, 1.818657, 1.818656, 
    1.818654, 1.818653, 1.818651, 1.818652, 1.818653, 1.818656, 1.818658, 
    1.818657, 1.818659, 1.818655, 1.818656, 1.818656, 1.818658, 1.818653, 
    1.818657, 1.818653, 1.818653, 1.818654, 1.818657, 1.818657, 1.818658, 
    1.818657, 1.818656, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.818653, 1.818654, 1.818656, 1.818658, 1.81866, 1.81866, 1.818662, 
    1.81866, 1.818664, 1.818661, 1.818666, 1.818657, 1.818661, 1.818654, 
    1.818655, 1.818656, 1.818659, 1.818658, 1.81866, 1.818655, 1.818653, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818659, 1.818663, 1.818666, 1.818668, 1.818669, 
    1.818669, 1.81867,
  1.818579, 1.818581, 1.818581, 1.818582, 1.818581, 1.818582, 1.81858, 
    1.818581, 1.81858, 1.818579, 1.818585, 1.818582, 1.818588, 1.818586, 
    1.818591, 1.818588, 1.818591, 1.818591, 1.818593, 1.818592, 1.818595, 
    1.818593, 1.818596, 1.818594, 1.818595, 1.818593, 1.818583, 1.818585, 
    1.818583, 1.818583, 1.818583, 1.818581, 1.818581, 1.818579, 1.818579, 
    1.818581, 1.818583, 1.818582, 1.818584, 1.818584, 1.818587, 1.818586, 
    1.81859, 1.818589, 1.818592, 1.818591, 1.818592, 1.818592, 1.818592, 
    1.818591, 1.818591, 1.81859, 1.818586, 1.818587, 1.818583, 1.818581, 
    1.81858, 1.818579, 1.818579, 1.818579, 1.818581, 1.818582, 1.818583, 
    1.818584, 1.818584, 1.818586, 1.818588, 1.81859, 1.81859, 1.818591, 
    1.818591, 1.818592, 1.818592, 1.818593, 1.81859, 1.818592, 1.818589, 
    1.81859, 1.818585, 1.818582, 1.818582, 1.818581, 1.818579, 1.81858, 
    1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 1.818588, 
    1.818586, 1.818591, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818593, 1.818594, 1.818593, 1.818594, 1.818591, 1.818592, 1.818581, 
    1.818581, 1.818582, 1.81858, 1.81858, 1.818579, 1.81858, 1.818581, 
    1.818582, 1.818582, 1.818583, 1.818584, 1.818586, 1.818588, 1.81859, 
    1.818591, 1.81859, 1.818591, 1.81859, 1.81859, 1.818593, 1.818591, 
    1.818594, 1.818594, 1.818593, 1.818594, 1.818581, 1.818581, 1.81858, 
    1.818581, 1.818579, 1.81858, 1.818581, 1.818583, 1.818583, 1.818584, 
    1.818585, 1.818586, 1.818588, 1.81859, 1.818591, 1.818591, 1.818591, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818594, 1.818593, 
    1.818594, 1.818594, 1.818581, 1.818582, 1.818581, 1.818582, 1.818582, 
    1.818584, 1.818584, 1.818587, 1.818586, 1.818588, 1.818586, 1.818586, 
    1.818588, 1.818586, 1.81859, 1.818587, 1.818592, 1.818589, 1.818592, 
    1.818591, 1.818592, 1.818593, 1.818594, 1.818595, 1.818595, 1.818596, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.818585, 1.818586, 1.818588, 
    1.818588, 1.818589, 1.818589, 1.818587, 1.818588, 1.818584, 1.818585, 
    1.818584, 1.818583, 1.818588, 1.818585, 1.81859, 1.818588, 1.818593, 
    1.818591, 1.818595, 1.818596, 1.818598, 1.8186, 1.818584, 1.818583, 
    1.818584, 1.818586, 1.818587, 1.818589, 1.818589, 1.818589, 1.81859, 
    1.818591, 1.818589, 1.818591, 1.818585, 1.818588, 1.818583, 1.818585, 
    1.818586, 1.818585, 1.818587, 1.818588, 1.81859, 1.818589, 1.818596, 
    1.818593, 1.818601, 1.818599, 1.818583, 1.818584, 1.818586, 1.818585, 
    1.818589, 1.81859, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818592, 1.818589, 1.81859, 1.818586, 1.818587, 1.818587, 1.818586, 
    1.818588, 1.818589, 1.818589, 1.81859, 1.818591, 1.818589, 1.818596, 
    1.818592, 1.818585, 1.818586, 1.818586, 1.818586, 1.818589, 1.818588, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.81859, 1.81859, 
    1.818588, 1.818587, 1.818586, 1.818586, 1.818587, 1.818589, 1.818591, 
    1.818591, 1.818592, 1.818588, 1.81859, 1.818589, 1.818591, 1.818588, 
    1.818591, 1.818587, 1.818587, 1.818588, 1.81859, 1.818591, 1.818591, 
    1.818591, 1.818589, 1.818589, 1.818588, 1.818588, 1.818587, 1.818586, 
    1.818587, 1.818588, 1.818589, 1.818591, 1.818593, 1.818593, 1.818595, 
    1.818594, 1.818596, 1.818594, 1.818598, 1.818591, 1.818594, 1.818588, 
    1.818589, 1.81859, 1.818592, 1.818591, 1.818593, 1.818589, 1.818587, 
    1.818587, 1.818586, 1.818587, 1.818587, 1.818588, 1.818587, 1.818589, 
    1.818588, 1.818591, 1.818593, 1.818596, 1.818598, 1.8186, 1.818601, 
    1.818601, 1.818601,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.327509e-09, 1.333351e-09, 1.332215e-09, 1.336927e-09, 1.334313e-09, 
    1.337398e-09, 1.328693e-09, 1.333583e-09, 1.330462e-09, 1.328035e-09, 
    1.346071e-09, 1.337137e-09, 1.35535e-09, 1.349652e-09, 1.363964e-09, 
    1.354463e-09, 1.36588e-09, 1.36369e-09, 1.370281e-09, 1.368393e-09, 
    1.376823e-09, 1.371152e-09, 1.381193e-09, 1.375469e-09, 1.376364e-09, 
    1.370965e-09, 1.338935e-09, 1.344959e-09, 1.338578e-09, 1.339437e-09, 
    1.339051e-09, 1.334367e-09, 1.332007e-09, 1.327063e-09, 1.32796e-09, 
    1.331591e-09, 1.339823e-09, 1.337029e-09, 1.344071e-09, 1.343912e-09, 
    1.351752e-09, 1.348217e-09, 1.361394e-09, 1.357649e-09, 1.368472e-09, 
    1.36575e-09, 1.368344e-09, 1.367557e-09, 1.368354e-09, 1.364362e-09, 
    1.366073e-09, 1.36256e-09, 1.348879e-09, 1.3529e-09, 1.340908e-09, 
    1.333698e-09, 1.328908e-09, 1.325509e-09, 1.32599e-09, 1.326906e-09, 
    1.331613e-09, 1.336038e-09, 1.33941e-09, 1.341666e-09, 1.343889e-09, 
    1.350618e-09, 1.354178e-09, 1.362152e-09, 1.360713e-09, 1.36315e-09, 
    1.365479e-09, 1.369389e-09, 1.368745e-09, 1.370468e-09, 1.363086e-09, 
    1.367992e-09, 1.359893e-09, 1.362108e-09, 1.344494e-09, 1.337783e-09, 
    1.33493e-09, 1.332433e-09, 1.326359e-09, 1.330554e-09, 1.3289e-09, 
    1.332834e-09, 1.335334e-09, 1.334098e-09, 1.341728e-09, 1.338762e-09, 
    1.354389e-09, 1.347658e-09, 1.365208e-09, 1.361008e-09, 1.366214e-09, 
    1.363557e-09, 1.368109e-09, 1.364013e-09, 1.371109e-09, 1.372654e-09, 
    1.371598e-09, 1.375655e-09, 1.363786e-09, 1.368344e-09, 1.334063e-09, 
    1.334265e-09, 1.335204e-09, 1.331075e-09, 1.330822e-09, 1.327038e-09, 
    1.330405e-09, 1.331839e-09, 1.335479e-09, 1.337632e-09, 1.339679e-09, 
    1.344179e-09, 1.349204e-09, 1.356232e-09, 1.36128e-09, 1.364664e-09, 
    1.362589e-09, 1.364421e-09, 1.362373e-09, 1.361413e-09, 1.372075e-09, 
    1.366089e-09, 1.375071e-09, 1.374574e-09, 1.370509e-09, 1.37463e-09, 
    1.334406e-09, 1.333246e-09, 1.329217e-09, 1.33237e-09, 1.326626e-09, 
    1.329841e-09, 1.33169e-09, 1.338824e-09, 1.340391e-09, 1.341844e-09, 
    1.344714e-09, 1.348398e-09, 1.35486e-09, 1.360482e-09, 1.365615e-09, 
    1.365238e-09, 1.365371e-09, 1.366517e-09, 1.363677e-09, 1.366984e-09, 
    1.367539e-09, 1.366088e-09, 1.374508e-09, 1.372102e-09, 1.374563e-09, 
    1.372997e-09, 1.333623e-09, 1.335576e-09, 1.334521e-09, 1.336505e-09, 
    1.335107e-09, 1.341322e-09, 1.343185e-09, 1.351904e-09, 1.348326e-09, 
    1.35402e-09, 1.348904e-09, 1.349811e-09, 1.354206e-09, 1.34918e-09, 
    1.360172e-09, 1.35272e-09, 1.366562e-09, 1.359121e-09, 1.367028e-09, 
    1.365592e-09, 1.36797e-09, 1.370099e-09, 1.372778e-09, 1.377721e-09, 
    1.376576e-09, 1.38071e-09, 1.338486e-09, 1.341019e-09, 1.340796e-09, 
    1.343446e-09, 1.345406e-09, 1.349654e-09, 1.356467e-09, 1.353905e-09, 
    1.358608e-09, 1.359553e-09, 1.352407e-09, 1.356794e-09, 1.342713e-09, 
    1.344989e-09, 1.343634e-09, 1.338686e-09, 1.354495e-09, 1.346382e-09, 
    1.361364e-09, 1.356969e-09, 1.369796e-09, 1.363417e-09, 1.375946e-09, 
    1.381303e-09, 1.386344e-09, 1.392235e-09, 1.342401e-09, 1.34068e-09, 
    1.343761e-09, 1.348024e-09, 1.351979e-09, 1.357237e-09, 1.357775e-09, 
    1.35876e-09, 1.361311e-09, 1.363456e-09, 1.359071e-09, 1.363994e-09, 
    1.345516e-09, 1.3552e-09, 1.34003e-09, 1.344598e-09, 1.347772e-09, 
    1.34638e-09, 1.353612e-09, 1.355317e-09, 1.362244e-09, 1.358663e-09, 
    1.379981e-09, 1.370549e-09, 1.396721e-09, 1.389407e-09, 1.340079e-09, 
    1.342395e-09, 1.350455e-09, 1.34662e-09, 1.357588e-09, 1.360287e-09, 
    1.362482e-09, 1.365287e-09, 1.36559e-09, 1.367252e-09, 1.364528e-09, 
    1.367145e-09, 1.357248e-09, 1.36167e-09, 1.349534e-09, 1.352488e-09, 
    1.351129e-09, 1.349638e-09, 1.354239e-09, 1.35914e-09, 1.359245e-09, 
    1.360816e-09, 1.365246e-09, 1.357632e-09, 1.381199e-09, 1.366645e-09, 
    1.34492e-09, 1.349381e-09, 1.350018e-09, 1.34829e-09, 1.360017e-09, 
    1.355768e-09, 1.367212e-09, 1.364119e-09, 1.369186e-09, 1.366668e-09, 
    1.366298e-09, 1.363063e-09, 1.36105e-09, 1.355963e-09, 1.351823e-09, 
    1.348541e-09, 1.349304e-09, 1.35291e-09, 1.35944e-09, 1.365618e-09, 
    1.364264e-09, 1.368801e-09, 1.356792e-09, 1.361828e-09, 1.359882e-09, 
    1.364956e-09, 1.353837e-09, 1.363306e-09, 1.351416e-09, 1.352459e-09, 
    1.355683e-09, 1.36217e-09, 1.363604e-09, 1.365137e-09, 1.364191e-09, 
    1.359606e-09, 1.358854e-09, 1.355605e-09, 1.354708e-09, 1.352232e-09, 
    1.350182e-09, 1.352055e-09, 1.354022e-09, 1.359608e-09, 1.364641e-09, 
    1.37013e-09, 1.371473e-09, 1.377885e-09, 1.372665e-09, 1.38128e-09, 
    1.373956e-09, 1.386633e-09, 1.363855e-09, 1.373741e-09, 1.35583e-09, 
    1.35776e-09, 1.36125e-09, 1.369254e-09, 1.364933e-09, 1.369986e-09, 
    1.358825e-09, 1.353034e-09, 1.351536e-09, 1.34874e-09, 1.3516e-09, 
    1.351367e-09, 1.354103e-09, 1.353224e-09, 1.359793e-09, 1.356264e-09, 
    1.366289e-09, 1.369946e-09, 1.380277e-09, 1.38661e-09, 1.393056e-09, 
    1.395902e-09, 1.396768e-09, 1.39713e-09 ;

 SOIL2_HR_S3 =
  9.482209e-11, 9.523934e-11, 9.515823e-11, 9.549478e-11, 9.530808e-11, 
    9.552846e-11, 9.490668e-11, 9.525591e-11, 9.503297e-11, 9.485964e-11, 
    9.614792e-11, 9.550979e-11, 9.68107e-11, 9.640374e-11, 9.742602e-11, 
    9.674738e-11, 9.756286e-11, 9.740643e-11, 9.787721e-11, 9.774234e-11, 
    9.834452e-11, 9.793946e-11, 9.865665e-11, 9.824778e-11, 9.831175e-11, 
    9.79261e-11, 9.56382e-11, 9.606847e-11, 9.561271e-11, 9.567407e-11, 
    9.564653e-11, 9.531195e-11, 9.514334e-11, 9.479019e-11, 9.48543e-11, 
    9.511367e-11, 9.570165e-11, 9.550205e-11, 9.600507e-11, 9.599371e-11, 
    9.655372e-11, 9.630122e-11, 9.724245e-11, 9.697494e-11, 9.774797e-11, 
    9.755356e-11, 9.773884e-11, 9.768265e-11, 9.773957e-11, 9.745445e-11, 
    9.757661e-11, 9.732572e-11, 9.634851e-11, 9.663571e-11, 9.577915e-11, 
    9.526412e-11, 9.492199e-11, 9.467923e-11, 9.471355e-11, 9.477898e-11, 
    9.511519e-11, 9.543129e-11, 9.567217e-11, 9.583331e-11, 9.599208e-11, 
    9.647268e-11, 9.672703e-11, 9.729655e-11, 9.719376e-11, 9.736788e-11, 
    9.753422e-11, 9.781349e-11, 9.776752e-11, 9.789057e-11, 9.736328e-11, 
    9.771373e-11, 9.713522e-11, 9.729344e-11, 9.603528e-11, 9.55559e-11, 
    9.535218e-11, 9.517382e-11, 9.473994e-11, 9.503957e-11, 9.492146e-11, 
    9.520246e-11, 9.538101e-11, 9.52927e-11, 9.583772e-11, 9.562583e-11, 
    9.674211e-11, 9.626129e-11, 9.751482e-11, 9.721485e-11, 9.758672e-11, 
    9.739697e-11, 9.772209e-11, 9.742948e-11, 9.793636e-11, 9.804674e-11, 
    9.797131e-11, 9.826104e-11, 9.741326e-11, 9.773884e-11, 9.529023e-11, 
    9.530463e-11, 9.537172e-11, 9.507678e-11, 9.505874e-11, 9.478843e-11, 
    9.502894e-11, 9.513137e-11, 9.539135e-11, 9.554514e-11, 9.569134e-11, 
    9.601276e-11, 9.637174e-11, 9.68737e-11, 9.72343e-11, 9.747603e-11, 
    9.73278e-11, 9.745867e-11, 9.731237e-11, 9.724381e-11, 9.800538e-11, 
    9.757775e-11, 9.821936e-11, 9.818386e-11, 9.78935e-11, 9.818786e-11, 
    9.531474e-11, 9.523186e-11, 9.49441e-11, 9.51693e-11, 9.475899e-11, 
    9.498867e-11, 9.512073e-11, 9.563027e-11, 9.574221e-11, 9.584602e-11, 
    9.605104e-11, 9.631414e-11, 9.677571e-11, 9.71773e-11, 9.75439e-11, 
    9.751704e-11, 9.752649e-11, 9.760839e-11, 9.740553e-11, 9.764169e-11, 
    9.768134e-11, 9.75777e-11, 9.81791e-11, 9.800729e-11, 9.818311e-11, 
    9.807123e-11, 9.525879e-11, 9.539826e-11, 9.53229e-11, 9.546461e-11, 
    9.536478e-11, 9.58087e-11, 9.59418e-11, 9.656457e-11, 9.630897e-11, 
    9.671574e-11, 9.635029e-11, 9.641504e-11, 9.672903e-11, 9.637003e-11, 
    9.715517e-11, 9.662289e-11, 9.761157e-11, 9.708006e-11, 9.764489e-11, 
    9.754231e-11, 9.771213e-11, 9.786423e-11, 9.805558e-11, 9.840864e-11, 
    9.832688e-11, 9.862215e-11, 9.560616e-11, 9.578705e-11, 9.577112e-11, 
    9.596042e-11, 9.610041e-11, 9.640384e-11, 9.68905e-11, 9.670749e-11, 
    9.704346e-11, 9.71109e-11, 9.660048e-11, 9.691388e-11, 9.590811e-11, 
    9.607062e-11, 9.597385e-11, 9.562044e-11, 9.674968e-11, 9.617016e-11, 
    9.724026e-11, 9.692632e-11, 9.784255e-11, 9.73869e-11, 9.828188e-11, 
    9.866449e-11, 9.902455e-11, 9.944538e-11, 9.588577e-11, 9.576286e-11, 
    9.598293e-11, 9.628742e-11, 9.65699e-11, 9.694547e-11, 9.698389e-11, 
    9.705426e-11, 9.72365e-11, 9.738974e-11, 9.707651e-11, 9.742814e-11, 
    9.610832e-11, 9.679997e-11, 9.571639e-11, 9.60427e-11, 9.626946e-11, 
    9.616998e-11, 9.668658e-11, 9.680833e-11, 9.73031e-11, 9.704734e-11, 
    9.857007e-11, 9.789637e-11, 9.976577e-11, 9.924336e-11, 9.571992e-11, 
    9.588534e-11, 9.646108e-11, 9.618715e-11, 9.697054e-11, 9.716337e-11, 
    9.732012e-11, 9.752051e-11, 9.754214e-11, 9.766087e-11, 9.746631e-11, 
    9.765318e-11, 9.694627e-11, 9.726218e-11, 9.639527e-11, 9.660627e-11, 
    9.65092e-11, 9.640273e-11, 9.673134e-11, 9.708145e-11, 9.708891e-11, 
    9.720117e-11, 9.751755e-11, 9.697371e-11, 9.865705e-11, 9.761748e-11, 
    9.606573e-11, 9.638438e-11, 9.642988e-11, 9.630644e-11, 9.714404e-11, 
    9.684055e-11, 9.765798e-11, 9.743705e-11, 9.779903e-11, 9.761916e-11, 
    9.75927e-11, 9.736167e-11, 9.721784e-11, 9.685447e-11, 9.65588e-11, 
    9.632434e-11, 9.637886e-11, 9.663641e-11, 9.710286e-11, 9.754411e-11, 
    9.744745e-11, 9.777152e-11, 9.691374e-11, 9.727343e-11, 9.713441e-11, 
    9.749689e-11, 9.670263e-11, 9.737903e-11, 9.652974e-11, 9.66042e-11, 
    9.683453e-11, 9.729784e-11, 9.740032e-11, 9.750976e-11, 9.744223e-11, 
    9.71147e-11, 9.706103e-11, 9.682893e-11, 9.676485e-11, 9.658799e-11, 
    9.644157e-11, 9.657535e-11, 9.671584e-11, 9.711483e-11, 9.747439e-11, 
    9.78664e-11, 9.796233e-11, 9.842039e-11, 9.804753e-11, 9.866283e-11, 
    9.813973e-11, 9.904524e-11, 9.741821e-11, 9.812433e-11, 9.6845e-11, 
    9.698282e-11, 9.723212e-11, 9.780387e-11, 9.749519e-11, 9.785618e-11, 
    9.705893e-11, 9.66453e-11, 9.653827e-11, 9.63386e-11, 9.654284e-11, 
    9.652622e-11, 9.672166e-11, 9.665885e-11, 9.712808e-11, 9.687603e-11, 
    9.759203e-11, 9.785332e-11, 9.85912e-11, 9.904355e-11, 9.950399e-11, 
    9.970727e-11, 9.976914e-11, 9.979501e-11 ;

 SOIL3C =
  5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782611, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782613, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782613, 
    5.782613, 5.782613 ;

 SOIL3C_TO_SOIL1C =
  2.6178e-11, 2.629317e-11, 2.627078e-11, 2.636367e-11, 2.631214e-11, 
    2.637296e-11, 2.620134e-11, 2.629774e-11, 2.62362e-11, 2.618836e-11, 
    2.654394e-11, 2.636781e-11, 2.672688e-11, 2.661455e-11, 2.689672e-11, 
    2.67094e-11, 2.693448e-11, 2.689131e-11, 2.702125e-11, 2.698402e-11, 
    2.715023e-11, 2.703843e-11, 2.723639e-11, 2.712353e-11, 2.714119e-11, 
    2.703474e-11, 2.640325e-11, 2.652202e-11, 2.639622e-11, 2.641315e-11, 
    2.640555e-11, 2.63132e-11, 2.626667e-11, 2.616919e-11, 2.618689e-11, 
    2.625848e-11, 2.642077e-11, 2.636568e-11, 2.650452e-11, 2.650138e-11, 
    2.665595e-11, 2.658626e-11, 2.684605e-11, 2.677221e-11, 2.698558e-11, 
    2.693192e-11, 2.698306e-11, 2.696755e-11, 2.698326e-11, 2.690456e-11, 
    2.693828e-11, 2.686903e-11, 2.659931e-11, 2.667858e-11, 2.644216e-11, 
    2.63e-11, 2.620557e-11, 2.613857e-11, 2.614804e-11, 2.61661e-11, 
    2.62589e-11, 2.634614e-11, 2.641263e-11, 2.645711e-11, 2.650093e-11, 
    2.663358e-11, 2.670379e-11, 2.686098e-11, 2.683261e-11, 2.688067e-11, 
    2.692658e-11, 2.700366e-11, 2.699098e-11, 2.702494e-11, 2.68794e-11, 
    2.697613e-11, 2.681645e-11, 2.686012e-11, 2.651286e-11, 2.638054e-11, 
    2.632431e-11, 2.627508e-11, 2.615532e-11, 2.623803e-11, 2.620542e-11, 
    2.628298e-11, 2.633227e-11, 2.630789e-11, 2.645833e-11, 2.639984e-11, 
    2.670795e-11, 2.657524e-11, 2.692123e-11, 2.683843e-11, 2.694107e-11, 
    2.68887e-11, 2.697844e-11, 2.689767e-11, 2.703758e-11, 2.706804e-11, 
    2.704722e-11, 2.712719e-11, 2.689319e-11, 2.698306e-11, 2.630721e-11, 
    2.631118e-11, 2.63297e-11, 2.62483e-11, 2.624331e-11, 2.616871e-11, 
    2.623509e-11, 2.626336e-11, 2.633512e-11, 2.637757e-11, 2.641792e-11, 
    2.650664e-11, 2.660572e-11, 2.674427e-11, 2.68438e-11, 2.691052e-11, 
    2.686961e-11, 2.690573e-11, 2.686535e-11, 2.684642e-11, 2.705663e-11, 
    2.69386e-11, 2.711569e-11, 2.710589e-11, 2.702574e-11, 2.710699e-11, 
    2.631398e-11, 2.62911e-11, 2.621167e-11, 2.627383e-11, 2.616058e-11, 
    2.622397e-11, 2.626043e-11, 2.640107e-11, 2.643196e-11, 2.646061e-11, 
    2.65172e-11, 2.658983e-11, 2.671722e-11, 2.682807e-11, 2.692925e-11, 
    2.692184e-11, 2.692445e-11, 2.694705e-11, 2.689106e-11, 2.695624e-11, 
    2.696719e-11, 2.693858e-11, 2.710458e-11, 2.705715e-11, 2.710568e-11, 
    2.70748e-11, 2.629853e-11, 2.633703e-11, 2.631623e-11, 2.635534e-11, 
    2.632779e-11, 2.645032e-11, 2.648705e-11, 2.665894e-11, 2.65884e-11, 
    2.670067e-11, 2.65998e-11, 2.661768e-11, 2.670434e-11, 2.660525e-11, 
    2.682196e-11, 2.667504e-11, 2.694793e-11, 2.680123e-11, 2.695712e-11, 
    2.692881e-11, 2.697569e-11, 2.701767e-11, 2.707048e-11, 2.716793e-11, 
    2.714536e-11, 2.722686e-11, 2.639441e-11, 2.644434e-11, 2.643994e-11, 
    2.649219e-11, 2.653083e-11, 2.661458e-11, 2.674891e-11, 2.669839e-11, 
    2.679112e-11, 2.680974e-11, 2.666886e-11, 2.675536e-11, 2.647775e-11, 
    2.652261e-11, 2.64959e-11, 2.639835e-11, 2.671004e-11, 2.655008e-11, 
    2.684544e-11, 2.675879e-11, 2.701168e-11, 2.688592e-11, 2.713294e-11, 
    2.723855e-11, 2.733793e-11, 2.745408e-11, 2.647159e-11, 2.643766e-11, 
    2.64984e-11, 2.658245e-11, 2.666042e-11, 2.676408e-11, 2.677468e-11, 
    2.679411e-11, 2.684441e-11, 2.68867e-11, 2.680025e-11, 2.68973e-11, 
    2.653302e-11, 2.672392e-11, 2.642484e-11, 2.65149e-11, 2.657749e-11, 
    2.655003e-11, 2.669262e-11, 2.672623e-11, 2.686279e-11, 2.67922e-11, 
    2.721249e-11, 2.702654e-11, 2.754251e-11, 2.739832e-11, 2.642581e-11, 
    2.647147e-11, 2.663038e-11, 2.655477e-11, 2.6771e-11, 2.682422e-11, 
    2.686749e-11, 2.69228e-11, 2.692877e-11, 2.696154e-11, 2.690784e-11, 
    2.695942e-11, 2.67643e-11, 2.685149e-11, 2.661222e-11, 2.667046e-11, 
    2.664366e-11, 2.661428e-11, 2.670498e-11, 2.680161e-11, 2.680367e-11, 
    2.683466e-11, 2.692198e-11, 2.677187e-11, 2.723649e-11, 2.694956e-11, 
    2.652126e-11, 2.660921e-11, 2.662177e-11, 2.65877e-11, 2.681889e-11, 
    2.673512e-11, 2.696074e-11, 2.689976e-11, 2.699967e-11, 2.695002e-11, 
    2.694272e-11, 2.687896e-11, 2.683926e-11, 2.673896e-11, 2.665736e-11, 
    2.659264e-11, 2.660769e-11, 2.667878e-11, 2.680752e-11, 2.692931e-11, 
    2.690263e-11, 2.699208e-11, 2.675532e-11, 2.68546e-11, 2.681623e-11, 
    2.691628e-11, 2.669705e-11, 2.688375e-11, 2.664933e-11, 2.666989e-11, 
    2.673346e-11, 2.686134e-11, 2.688962e-11, 2.691983e-11, 2.690119e-11, 
    2.681079e-11, 2.679598e-11, 2.673191e-11, 2.671422e-11, 2.666541e-11, 
    2.6625e-11, 2.666192e-11, 2.67007e-11, 2.681082e-11, 2.691007e-11, 
    2.701827e-11, 2.704474e-11, 2.717117e-11, 2.706826e-11, 2.723809e-11, 
    2.709371e-11, 2.734364e-11, 2.689456e-11, 2.708946e-11, 2.673635e-11, 
    2.677439e-11, 2.68432e-11, 2.700101e-11, 2.691581e-11, 2.701545e-11, 
    2.679539e-11, 2.668123e-11, 2.665169e-11, 2.659658e-11, 2.665295e-11, 
    2.664836e-11, 2.67023e-11, 2.668497e-11, 2.681448e-11, 2.674491e-11, 
    2.694254e-11, 2.701466e-11, 2.721832e-11, 2.734317e-11, 2.747026e-11, 
    2.752636e-11, 2.754344e-11, 2.755058e-11 ;

 SOIL3C_vr =
  20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00008, 20.00007, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  -7.709882e-21, -2.569961e-21, -1.003089e-36, 5.139921e-21, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, 0, 0, 1.28498e-20, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 1.027984e-20, 
    -1.28498e-20, -5.139921e-21, 5.015443e-37, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.027984e-20, 2.569961e-21, -1.541976e-20, -5.139921e-21, 
    1.28498e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    1.003089e-36, -1.28498e-20, 2.569961e-21, 2.569961e-21, 0, -5.139921e-21, 
    7.709882e-21, 1.798972e-20, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    1.003089e-36, -1.798972e-20, 2.569961e-21, 0, -7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -1.798972e-20, 2.569961e-21, -7.709882e-21, -1.28498e-20, -1.28498e-20, 
    2.569961e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    2.055969e-20, 2.569961e-21, 1.027984e-20, 7.709882e-21, -7.709882e-21, 
    7.709882e-21, -1.541976e-20, 5.139921e-21, -7.709882e-21, -7.709882e-21, 
    1.027984e-20, 2.569961e-21, -1.027984e-20, -2.569961e-21, -1.541976e-20, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    2.569961e-21, 2.055969e-20, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, 2.312965e-20, 2.569961e-21, 1.28498e-20, 7.709882e-21, 
    1.541976e-20, 2.569961e-21, 2.569961e-21, -1.027984e-20, -1.003089e-36, 
    1.003089e-36, -2.569961e-21, 1.798972e-20, 7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 5.139921e-21, 0, 1.798972e-20, 0, 
    -7.709882e-21, 5.139921e-21, 7.709882e-21, 1.541976e-20, 7.709882e-21, 0, 
    1.003089e-36, 2.055969e-20, 2.312965e-20, -2.569961e-21, -7.709882e-21, 
    1.003089e-36, 0, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -1.541976e-20, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 1.28498e-20, 2.569961e-21, -3.083953e-20, 1.027984e-20, 
    -1.28498e-20, -2.569961e-21, 5.139921e-21, 1.798972e-20, 2.055969e-20, 
    -1.28498e-20, -1.027984e-20, -2.569961e-21, -1.003089e-36, -1.28498e-20, 
    0, 2.569961e-21, -1.003089e-36, -1.28498e-20, -1.541976e-20, 1.28498e-20, 
    -1.798972e-20, 7.709882e-21, 0, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, 1.28498e-20, -7.709882e-21, 1.798972e-20, 
    -1.027984e-20, -1.027984e-20, -1.541976e-20, -5.139921e-21, 1.28498e-20, 
    2.312965e-20, -2.569961e-21, -2.055969e-20, 1.027984e-20, 2.569961e-21, 
    -1.003089e-36, 2.055969e-20, 5.139921e-21, 2.055969e-20, -1.28498e-20, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, -7.709882e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -1.541976e-20, 2.569961e-21, 7.709882e-21, 
    7.709882e-21, 7.709882e-21, 1.28498e-20, 1.28498e-20, -5.139921e-21, 
    7.709882e-21, -7.709882e-21, -2.569961e-21, -1.541976e-20, -1.541976e-20, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, 2.569961e-21, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, 2.569961e-21, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    7.709882e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, -1.003089e-36, 
    -2.569961e-21, 0, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, 1.541976e-20, -1.28498e-20, -1.027984e-20, 7.709882e-21, 
    0, -7.709882e-21, -5.139921e-21, -2.055969e-20, 1.541976e-20, 
    5.139921e-21, 1.28498e-20, 5.139921e-21, 1.541976e-20, 1.798972e-20, 
    1.541976e-20, 1.003089e-36, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.003089e-36, 0, -7.709882e-21, 
    -5.139921e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 
    -1.798972e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 1.003089e-36, 7.709882e-21, 
    2.569961e-21, -1.541976e-20, -2.569961e-21, -5.139921e-21, 2.312965e-20, 
    2.569961e-21, 2.569961e-21, 0, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -1.798972e-20, 7.709882e-21, 7.709882e-21, -1.003089e-36, 2.569961e-21, 
    7.709882e-21, -1.027984e-20, -5.139921e-21, 2.055969e-20, -1.28498e-20, 
    -5.139921e-21, 0, -2.312965e-20, -5.139921e-21, -5.139921e-21, 
    2.312965e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 1.798972e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.798972e-20, -1.027984e-20, -2.569961e-21, -1.541976e-20, -5.139921e-21, 
    0, 1.027984e-20, 1.003089e-36, 1.541976e-20, -2.569961e-21, 
    -1.027984e-20, 1.541976e-20, 1.541976e-20, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, -5.139921e-21, 1.027984e-20,
  -7.709882e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -1.003089e-36, -7.709882e-21, -1.541976e-20, 1.027984e-20, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 0, -5.139921e-21, 0, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, -1.003089e-36, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, -1.541976e-20, -2.569961e-21, -1.003089e-36, 
    2.569961e-21, -1.003089e-36, 1.027984e-20, -5.139921e-21, 0, 
    -7.709882e-21, -1.027984e-20, 7.709882e-21, 1.027984e-20, -1.027984e-20, 
    1.28498e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, 2.569961e-21, 
    5.139921e-21, 0, 0, 1.027984e-20, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, -1.003089e-36, 0, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 0, 7.709882e-21, 7.709882e-21, 2.569961e-21, 
    0, -7.709882e-21, 1.541976e-20, 5.139921e-21, 0, 0, 7.709882e-21, 
    -7.709882e-21, 7.709882e-21, 5.139921e-21, 0, 0, 1.027984e-20, 0, 
    7.709882e-21, 5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 1.003089e-36, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 
    7.709882e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 1.28498e-20, -2.569961e-21, -2.569961e-21, 
    0, -2.569961e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 7.709882e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, 1.28498e-20, 0, 2.569961e-21, 
    -1.541976e-20, -2.569961e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, 0, 
    1.28498e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 1.027984e-20, 
    -7.709882e-21, -7.709882e-21, 1.541976e-20, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -1.541976e-20, 0, -1.28498e-20, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, 1.28498e-20, 7.709882e-21, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    1.541976e-20, -1.027984e-20, 2.569961e-21, 2.569961e-21, 0, 
    -7.709882e-21, -5.139921e-21, -1.541976e-20, -1.003089e-36, 0, 0, 
    -1.027984e-20, 7.709882e-21, 1.541976e-20, -2.569961e-21, -7.709882e-21, 
    1.003089e-36, 7.709882e-21, 1.798972e-20, -1.541976e-20, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 0, 1.798972e-20, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, 0, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, -5.139921e-21, 7.709882e-21, 
    7.709882e-21, 0, 1.28498e-20, 7.709882e-21, 0, -7.709882e-21, 0, 
    1.027984e-20, 0, 1.28498e-20, 2.569961e-21, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, 
    1.003089e-36, -2.569961e-21, -1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, 1.027984e-20, -7.709882e-21, 0, 2.569961e-21, 0, 
    -1.798972e-20, 7.709882e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 1.28498e-20, 
    -1.28498e-20, 2.569961e-21, -1.541976e-20, 5.139921e-21, 7.709882e-21, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    2.312965e-20, 2.569961e-21, 7.709882e-21, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 1.003089e-36, -5.139921e-21, 
    7.709882e-21, 0, 5.139921e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -1.28498e-20, 0, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    0, 5.139921e-21, 1.003089e-36, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, 5.139921e-21, 1.027984e-20, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, -7.709882e-21, 1.798972e-20, -7.709882e-21, 
    7.709882e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 
    1.003089e-36, -7.709882e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 1.027984e-20, 1.28498e-20, 1.28498e-20, -1.798972e-20, 
    1.027984e-20,
  -1.28498e-20, -1.027984e-20, 1.003089e-36, 2.569961e-21, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 
    1.798972e-20, -5.139921e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    2.569961e-21, 0, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -7.709882e-21, 2.569961e-21, -1.003089e-36, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 1.28498e-20, 
    1.541976e-20, -2.569961e-21, 0, 7.709882e-21, 1.541976e-20, 
    -1.027984e-20, 0, 0, 1.541976e-20, -5.139921e-21, 2.312965e-20, 
    -5.139921e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 1.798972e-20, -5.139921e-21, -1.28498e-20, -2.569961e-21, 
    1.027984e-20, -1.027984e-20, -7.709882e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, 0, 
    -7.709882e-21, -7.709882e-21, -1.541976e-20, 5.139921e-21, 1.541976e-20, 
    1.027984e-20, 7.709882e-21, 1.28498e-20, 5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 0, 2.569961e-21, -2.055969e-20, 5.139921e-21, 
    -1.541976e-20, 1.541976e-20, 0, 5.139921e-21, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 7.709882e-21, 
    1.798972e-20, 5.139921e-21, -1.003089e-36, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, -7.709882e-21, -5.139921e-21, 
    1.28498e-20, 1.541976e-20, -2.569961e-21, 0, -7.709882e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 0, -2.569961e-21, 7.709882e-21, 
    1.003089e-36, 1.003089e-36, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, 2.569961e-21, 0, -2.569961e-21, 1.003089e-36, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, -1.003089e-36, 5.139921e-21, 
    1.027984e-20, 7.709882e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, 1.027984e-20, -1.541976e-20, 2.055969e-20, 
    -7.709882e-21, 5.139921e-21, -1.541976e-20, 2.312965e-20, -5.139921e-21, 
    2.569961e-21, 0, -1.027984e-20, -2.569961e-21, 1.541976e-20, 
    -1.798972e-20, -1.798972e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, -1.798972e-20, 1.541976e-20, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, -1.003089e-36, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 1.003089e-36, 2.569961e-21, 1.541976e-20, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, 0, 
    -7.709882e-21, -1.027984e-20, 1.28498e-20, 7.709882e-21, -2.569961e-21, 
    -1.027984e-20, -1.28498e-20, -1.541976e-20, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, -1.027984e-20, 1.541976e-20, 1.798972e-20, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, 1.003089e-36, -1.541976e-20, -7.709882e-21, 
    0, 1.541976e-20, 2.569961e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, 1.28498e-20, -1.003089e-36, 
    5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 1.003089e-36, 
    2.569961e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 0, 2.569961e-21, 
    1.027984e-20, 1.28498e-20, 1.541976e-20, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    0, 0, -5.139921e-21, 2.569961e-21, 1.541976e-20, -2.569961e-21, 
    2.569961e-21, -1.027984e-20, -1.003089e-36, -1.027984e-20, -2.569961e-21, 
    5.139921e-21, -1.003089e-36, 2.569961e-21, -1.541976e-20, 2.055969e-20, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 1.28498e-20, 1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    7.709882e-21, 0, -1.003089e-36, 1.798972e-20, 7.709882e-21, 
    -1.003089e-36, -5.139921e-21, -1.28498e-20, -1.28498e-20, -1.28498e-20, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, 2.569961e-21, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 2.569961e-21, -2.569961e-21, -1.003089e-36, 
    2.569961e-21, -7.709882e-21, -1.541976e-20, 0, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 0, 1.027984e-20, 7.709882e-21, 2.569961e-21, 
    0, 2.569961e-21, 7.709882e-21, -1.003089e-36, 1.541976e-20, 7.709882e-21, 
    -7.709882e-21, 0, -2.569961e-21, 0, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, -1.027984e-20, -7.709882e-21, 7.709882e-21, 5.139921e-21, 
    1.28498e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, -1.003089e-36, 0,
  1.798972e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, -1.28498e-20, 
    -1.541976e-20, -1.28498e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, 1.541976e-20, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, -1.798972e-20, 0, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    0, 5.139921e-21, -1.28498e-20, 1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, -5.139921e-21, 
    1.541976e-20, 1.003089e-36, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -1.027984e-20, -1.28498e-20, -5.139921e-21, 2.055969e-20, -2.569961e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, 1.003089e-36, 7.709882e-21, 
    -1.003089e-36, -2.569961e-21, 0, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.28498e-20, -7.709882e-21, 0, 
    7.709882e-21, -1.541976e-20, -7.709882e-21, 1.003089e-36, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 1.28498e-20, 1.798972e-20, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, -5.139921e-21, -1.28498e-20, -2.569961e-21, 
    5.139921e-21, 2.312965e-20, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.798972e-20, 1.541976e-20, 2.055969e-20, -1.003089e-36, -5.139921e-21, 
    5.139921e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, 
    1.003089e-36, -5.139921e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -1.798972e-20, -2.569961e-21, -2.569961e-21, -1.541976e-20, 5.139921e-21, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, -1.003089e-36, 5.139921e-21, 
    5.139921e-21, -7.709882e-21, 0, 1.541976e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    1.28498e-20, 5.139921e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 5.139921e-21, 1.798972e-20, -1.28498e-20, 
    1.027984e-20, 2.569961e-21, -5.139921e-21, 0, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, 7.709882e-21, 1.003089e-36, -7.709882e-21, 1.541976e-20, 
    2.569961e-21, 1.027984e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.798972e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, 2.569961e-21, -1.027984e-20, 5.139921e-21, -1.28498e-20, 
    0, 2.569961e-21, 1.003089e-36, -5.139921e-21, 0, -1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 0, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, 1.798972e-20, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 1.798972e-20, 5.139921e-21, -1.28498e-20, -7.709882e-21, 
    -1.541976e-20, 1.003089e-36, 0, 7.709882e-21, -1.28498e-20, 1.027984e-20, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, 0, 5.139921e-21, 1.027984e-20, 1.003089e-36, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, 7.709882e-21, -1.003089e-36, 
    7.709882e-21, -1.541976e-20, 1.28498e-20, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 1.541976e-20, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, 1.28498e-20, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, 0, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, 1.541976e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -2.312965e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 1.28498e-20, 
    -2.569961e-21, -1.798972e-20, 1.003089e-36, -2.569961e-21, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 1.027984e-20, -1.798972e-20, -1.003089e-36, -5.139921e-21, 
    7.709882e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 0, 5.139921e-21, 
    2.569961e-21, -7.709882e-21, 1.28498e-20, -1.541976e-20, 7.709882e-21, 
    5.139921e-21, -1.541976e-20, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    2.055969e-20, 1.027984e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, 
    -2.055969e-20, 7.709882e-21, -1.003089e-36, -1.28498e-20, -1.027984e-20, 
    -2.569961e-21, 1.003089e-36, -2.569961e-20, 1.541976e-20, -1.003089e-36, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, 0, -2.569961e-21, 
    -1.003089e-36, -1.003089e-36, 1.003089e-36, -2.569961e-21, 1.798972e-20, 
    -7.709882e-21, 5.139921e-21, 1.541976e-20, -7.709882e-21,
  -1.28498e-20, -2.569961e-21, -1.541976e-20, -1.28498e-20, 1.003089e-36, 
    1.027984e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, -2.569961e-21, -1.798972e-20, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    1.003089e-36, -5.139921e-21, 1.541976e-20, 2.312965e-20, -1.003089e-36, 
    -1.003089e-36, 2.569961e-21, -7.709882e-21, -1.798972e-20, -5.139921e-21, 
    -2.569961e-21, 1.28498e-20, 1.027984e-20, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 1.027984e-20, 1.798972e-20, 1.003089e-36, 5.139921e-21, 
    2.569961e-21, 1.28498e-20, -7.709882e-21, -1.28498e-20, -1.027984e-20, 
    -2.569961e-20, 2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    1.798972e-20, -2.569961e-21, -1.798972e-20, -7.709882e-21, -1.28498e-20, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, -2.569961e-20, 2.569961e-21, 
    1.541976e-20, 5.139921e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    1.28498e-20, 0, -5.139921e-21, 7.709882e-21, -7.709882e-21, 
    -1.027984e-20, 5.139921e-21, -1.28498e-20, 0, -3.083953e-20, 
    -1.027984e-20, 2.569961e-21, -1.798972e-20, -5.139921e-21, -5.139921e-21, 
    2.055969e-20, -1.28498e-20, -1.541976e-20, -2.569961e-21, -1.027984e-20, 
    1.027984e-20, 0, 2.569961e-21, 2.826957e-20, 7.709882e-21, -1.798972e-20, 
    1.28498e-20, -2.569961e-21, -1.28498e-20, 2.312965e-20, -2.569961e-21, 
    -2.569961e-21, 2.055969e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -1.541976e-20, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 2.312965e-20, 
    2.569961e-21, 2.569961e-21, -1.28498e-20, -1.027984e-20, 2.569961e-21, 
    1.027984e-20, -1.027984e-20, -7.709882e-21, -2.055969e-20, -5.139921e-21, 
    -1.541976e-20, -1.798972e-20, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 2.055969e-20, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 1.798972e-20, -1.003089e-36, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, -1.027984e-20, -7.709882e-21, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 1.28498e-20, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -1.798972e-20, -7.709882e-21, -1.28498e-20, 
    2.569961e-21, 1.28498e-20, -2.569961e-20, -1.798972e-20, 1.027984e-20, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, 1.003089e-36, -2.569961e-20, 
    2.569961e-21, -2.569961e-21, 2.312965e-20, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, 7.709882e-21, 0, 5.139921e-21, -7.709882e-21, -2.055969e-20, 
    -1.027984e-20, -1.027984e-20, 0, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.003089e-36, -1.027984e-20, 3.009266e-36, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -2.055969e-20, -1.027984e-20, -1.28498e-20, 
    5.139921e-21, -2.055969e-20, 2.569961e-21, -1.798972e-20, -7.709882e-21, 
    0, 1.28498e-20, -5.139921e-21, 1.28498e-20, -1.798972e-20, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -2.826957e-20, 1.28498e-20, 1.027984e-20, 
    -7.709882e-21, 5.139921e-21, 1.28498e-20, -1.027984e-20, 2.055969e-20, 
    -1.027984e-20, 1.28498e-20, 1.798972e-20, -1.003089e-36, -1.027984e-20, 
    -1.003089e-36, 2.569961e-21, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -2.826957e-20, 1.027984e-20, -1.28498e-20, -2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -1.28498e-20, -2.569961e-20, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -1.027984e-20, -2.569961e-21, 1.541976e-20, 7.709882e-21, 
    -1.027984e-20, 5.139921e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 1.003089e-36, 1.003089e-36, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 2.312965e-20, 1.027984e-20, 1.003089e-36, 
    -2.055969e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    1.003089e-36, -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.28498e-20, 
    -7.709882e-21, 3.009266e-36, 1.28498e-20, 1.027984e-20, 1.027984e-20, 
    2.569961e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -1.28498e-20, 7.709882e-21, 1.541976e-20, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, 
    7.709882e-21, 1.003089e-36, 2.569961e-21, -1.027984e-20, 1.28498e-20, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, 7.709882e-21, 1.798972e-20, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 0, -1.003089e-36, 2.569961e-21, -1.28498e-20, 
    -7.709882e-21, -7.709882e-21, 1.541976e-20, 1.541976e-20, 2.569961e-21, 
    1.003089e-36, -2.569961e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -1.003089e-36, 2.569961e-21, 5.139921e-21, -1.798972e-20, 
    1.541976e-20, 1.28498e-20, 2.569961e-21, -1.541976e-20, 2.569961e-21, 
    1.027984e-20, -2.826957e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    -1.541976e-20, -5.139921e-21, -7.709882e-21, -1.541976e-20, 0, 
    5.139921e-21, -7.709882e-21, 0, 0, -5.139921e-21, 1.027984e-20,
  6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.288484e-12, 5.311751e-12, 5.307227e-12, 5.325994e-12, 5.315583e-12, 
    5.327872e-12, 5.293201e-12, 5.312675e-12, 5.300243e-12, 5.290578e-12, 
    5.362413e-12, 5.326831e-12, 5.39937e-12, 5.376678e-12, 5.43368e-12, 
    5.395839e-12, 5.44131e-12, 5.432588e-12, 5.458838e-12, 5.451318e-12, 
    5.484896e-12, 5.462309e-12, 5.5023e-12, 5.479501e-12, 5.483068e-12, 
    5.461564e-12, 5.333991e-12, 5.357983e-12, 5.332569e-12, 5.335991e-12, 
    5.334456e-12, 5.315799e-12, 5.306397e-12, 5.286706e-12, 5.29028e-12, 
    5.304743e-12, 5.337529e-12, 5.326399e-12, 5.354448e-12, 5.353815e-12, 
    5.385041e-12, 5.370961e-12, 5.423444e-12, 5.408528e-12, 5.451632e-12, 
    5.440791e-12, 5.451123e-12, 5.44799e-12, 5.451163e-12, 5.435265e-12, 
    5.442077e-12, 5.428087e-12, 5.373598e-12, 5.389612e-12, 5.34185e-12, 
    5.313132e-12, 5.294055e-12, 5.280519e-12, 5.282432e-12, 5.286081e-12, 
    5.304828e-12, 5.322453e-12, 5.335885e-12, 5.34487e-12, 5.353724e-12, 
    5.380522e-12, 5.394704e-12, 5.426461e-12, 5.420729e-12, 5.430439e-12, 
    5.439713e-12, 5.455286e-12, 5.452722e-12, 5.459583e-12, 5.430182e-12, 
    5.449722e-12, 5.417465e-12, 5.426287e-12, 5.356133e-12, 5.329402e-12, 
    5.318042e-12, 5.308097e-12, 5.283904e-12, 5.300612e-12, 5.294025e-12, 
    5.309694e-12, 5.31965e-12, 5.314726e-12, 5.345116e-12, 5.333301e-12, 
    5.395545e-12, 5.368735e-12, 5.438631e-12, 5.421906e-12, 5.44264e-12, 
    5.43206e-12, 5.450189e-12, 5.433873e-12, 5.462136e-12, 5.468291e-12, 
    5.464085e-12, 5.48024e-12, 5.432968e-12, 5.451123e-12, 5.314588e-12, 
    5.315391e-12, 5.319132e-12, 5.302686e-12, 5.30168e-12, 5.286608e-12, 
    5.300019e-12, 5.30573e-12, 5.320227e-12, 5.328802e-12, 5.336954e-12, 
    5.354877e-12, 5.374893e-12, 5.402882e-12, 5.42299e-12, 5.436469e-12, 
    5.428203e-12, 5.4355e-12, 5.427343e-12, 5.42352e-12, 5.465985e-12, 
    5.442141e-12, 5.477917e-12, 5.475937e-12, 5.459746e-12, 5.47616e-12, 
    5.315955e-12, 5.311333e-12, 5.295288e-12, 5.307845e-12, 5.284966e-12, 
    5.297773e-12, 5.305137e-12, 5.333549e-12, 5.33979e-12, 5.345579e-12, 
    5.357011e-12, 5.371682e-12, 5.397419e-12, 5.419811e-12, 5.440253e-12, 
    5.438755e-12, 5.439282e-12, 5.443849e-12, 5.432537e-12, 5.445706e-12, 
    5.447916e-12, 5.442138e-12, 5.475672e-12, 5.466092e-12, 5.475895e-12, 
    5.469657e-12, 5.312835e-12, 5.320612e-12, 5.31641e-12, 5.324312e-12, 
    5.318745e-12, 5.343498e-12, 5.35092e-12, 5.385645e-12, 5.371393e-12, 
    5.394075e-12, 5.373697e-12, 5.377308e-12, 5.394816e-12, 5.374798e-12, 
    5.418577e-12, 5.388897e-12, 5.444026e-12, 5.414389e-12, 5.445884e-12, 
    5.440164e-12, 5.449634e-12, 5.458115e-12, 5.468784e-12, 5.488471e-12, 
    5.483912e-12, 5.500375e-12, 5.332204e-12, 5.342291e-12, 5.341403e-12, 
    5.351958e-12, 5.359764e-12, 5.376683e-12, 5.403819e-12, 5.393615e-12, 
    5.412348e-12, 5.416109e-12, 5.387648e-12, 5.405123e-12, 5.349041e-12, 
    5.358103e-12, 5.352707e-12, 5.333001e-12, 5.395967e-12, 5.363653e-12, 
    5.423322e-12, 5.405817e-12, 5.456905e-12, 5.431499e-12, 5.481402e-12, 
    5.502737e-12, 5.522814e-12, 5.546279e-12, 5.347796e-12, 5.340942e-12, 
    5.353213e-12, 5.370191e-12, 5.385943e-12, 5.406885e-12, 5.409027e-12, 
    5.41295e-12, 5.423112e-12, 5.431656e-12, 5.414192e-12, 5.433798e-12, 
    5.360205e-12, 5.398772e-12, 5.338351e-12, 5.356546e-12, 5.36919e-12, 
    5.363643e-12, 5.392449e-12, 5.399238e-12, 5.426827e-12, 5.412564e-12, 
    5.497472e-12, 5.459907e-12, 5.564143e-12, 5.535014e-12, 5.338547e-12, 
    5.347772e-12, 5.379875e-12, 5.3646e-12, 5.408283e-12, 5.419035e-12, 
    5.427775e-12, 5.438949e-12, 5.440155e-12, 5.446775e-12, 5.435927e-12, 
    5.446346e-12, 5.406929e-12, 5.424544e-12, 5.376205e-12, 5.387971e-12, 
    5.382558e-12, 5.376621e-12, 5.394944e-12, 5.414467e-12, 5.414883e-12, 
    5.421143e-12, 5.438784e-12, 5.40846e-12, 5.502322e-12, 5.444356e-12, 
    5.35783e-12, 5.375598e-12, 5.378135e-12, 5.371252e-12, 5.417957e-12, 
    5.401034e-12, 5.446614e-12, 5.434295e-12, 5.454479e-12, 5.44445e-12, 
    5.442974e-12, 5.430092e-12, 5.422072e-12, 5.401811e-12, 5.385324e-12, 
    5.37225e-12, 5.37529e-12, 5.389651e-12, 5.415661e-12, 5.440265e-12, 
    5.434875e-12, 5.452945e-12, 5.405115e-12, 5.425172e-12, 5.41742e-12, 
    5.437632e-12, 5.393344e-12, 5.43106e-12, 5.383703e-12, 5.387856e-12, 
    5.400699e-12, 5.426532e-12, 5.432247e-12, 5.43835e-12, 5.434584e-12, 
    5.416321e-12, 5.413328e-12, 5.400386e-12, 5.396813e-12, 5.386951e-12, 
    5.378787e-12, 5.386247e-12, 5.394081e-12, 5.416328e-12, 5.436377e-12, 
    5.458235e-12, 5.463584e-12, 5.489126e-12, 5.468335e-12, 5.502645e-12, 
    5.473477e-12, 5.523967e-12, 5.433244e-12, 5.472618e-12, 5.401283e-12, 
    5.408968e-12, 5.422868e-12, 5.454749e-12, 5.437537e-12, 5.457666e-12, 
    5.413211e-12, 5.390148e-12, 5.384179e-12, 5.373045e-12, 5.384434e-12, 
    5.383507e-12, 5.394405e-12, 5.390903e-12, 5.417067e-12, 5.403013e-12, 
    5.442937e-12, 5.457506e-12, 5.49865e-12, 5.523873e-12, 5.549547e-12, 
    5.560882e-12, 5.564332e-12, 5.565774e-12 ;

 SOIL3N_vr =
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818188, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.199533e-11, 3.213609e-11, 3.210873e-11, 3.222226e-11, 3.215928e-11, 
    3.223363e-11, 3.202387e-11, 3.214168e-11, 3.206647e-11, 3.2008e-11, 
    3.24426e-11, 3.222732e-11, 3.266619e-11, 3.25289e-11, 3.287377e-11, 
    3.264482e-11, 3.291993e-11, 3.286716e-11, 3.302597e-11, 3.298047e-11, 
    3.318362e-11, 3.304697e-11, 3.328891e-11, 3.315098e-11, 3.317256e-11, 
    3.304246e-11, 3.227064e-11, 3.24158e-11, 3.226205e-11, 3.228275e-11, 
    3.227345e-11, 3.216058e-11, 3.210371e-11, 3.198457e-11, 3.20062e-11, 
    3.20937e-11, 3.229205e-11, 3.222472e-11, 3.239441e-11, 3.239058e-11, 
    3.257949e-11, 3.249432e-11, 3.281184e-11, 3.272159e-11, 3.298237e-11, 
    3.291679e-11, 3.297929e-11, 3.296034e-11, 3.297954e-11, 3.288336e-11, 
    3.292457e-11, 3.283993e-11, 3.251027e-11, 3.260716e-11, 3.23182e-11, 
    3.214445e-11, 3.202904e-11, 3.194714e-11, 3.195871e-11, 3.198079e-11, 
    3.209421e-11, 3.220084e-11, 3.228211e-11, 3.233647e-11, 3.239003e-11, 
    3.255216e-11, 3.263796e-11, 3.283009e-11, 3.279541e-11, 3.285415e-11, 
    3.291026e-11, 3.300448e-11, 3.298897e-11, 3.303048e-11, 3.28526e-11, 
    3.297082e-11, 3.277566e-11, 3.282904e-11, 3.24046e-11, 3.224288e-11, 
    3.217416e-11, 3.211399e-11, 3.196762e-11, 3.20687e-11, 3.202885e-11, 
    3.212365e-11, 3.218388e-11, 3.215409e-11, 3.233795e-11, 3.226647e-11, 
    3.264305e-11, 3.248084e-11, 3.290372e-11, 3.280253e-11, 3.292797e-11, 
    3.286396e-11, 3.297364e-11, 3.287493e-11, 3.304593e-11, 3.308316e-11, 
    3.305772e-11, 3.315545e-11, 3.286946e-11, 3.297929e-11, 3.215326e-11, 
    3.215811e-11, 3.218075e-11, 3.208125e-11, 3.207516e-11, 3.198397e-11, 
    3.206511e-11, 3.209967e-11, 3.218737e-11, 3.223925e-11, 3.228857e-11, 
    3.239701e-11, 3.25181e-11, 3.268744e-11, 3.280909e-11, 3.289063e-11, 
    3.284063e-11, 3.288478e-11, 3.283543e-11, 3.281229e-11, 3.306921e-11, 
    3.292495e-11, 3.31414e-11, 3.312942e-11, 3.303147e-11, 3.313077e-11, 
    3.216153e-11, 3.213357e-11, 3.203649e-11, 3.211246e-11, 3.197404e-11, 
    3.205152e-11, 3.209608e-11, 3.226797e-11, 3.230573e-11, 3.234075e-11, 
    3.240992e-11, 3.249868e-11, 3.265438e-11, 3.278986e-11, 3.291353e-11, 
    3.290447e-11, 3.290766e-11, 3.293529e-11, 3.286685e-11, 3.294652e-11, 
    3.29599e-11, 3.292493e-11, 3.312782e-11, 3.306985e-11, 3.312917e-11, 
    3.309143e-11, 3.214265e-11, 3.21897e-11, 3.216428e-11, 3.221208e-11, 
    3.217841e-11, 3.232816e-11, 3.237306e-11, 3.258315e-11, 3.249693e-11, 
    3.263415e-11, 3.251087e-11, 3.253271e-11, 3.263863e-11, 3.251753e-11, 
    3.278239e-11, 3.260283e-11, 3.293636e-11, 3.275705e-11, 3.29476e-11, 
    3.2913e-11, 3.297028e-11, 3.302159e-11, 3.308614e-11, 3.320525e-11, 
    3.317767e-11, 3.327727e-11, 3.225984e-11, 3.232086e-11, 3.231549e-11, 
    3.237935e-11, 3.242657e-11, 3.252893e-11, 3.269311e-11, 3.263137e-11, 
    3.274471e-11, 3.276746e-11, 3.259527e-11, 3.270099e-11, 3.23617e-11, 
    3.241652e-11, 3.238388e-11, 3.226465e-11, 3.26456e-11, 3.24501e-11, 
    3.28111e-11, 3.270519e-11, 3.301428e-11, 3.286057e-11, 3.316248e-11, 
    3.329156e-11, 3.341302e-11, 3.355499e-11, 3.235416e-11, 3.23127e-11, 
    3.238694e-11, 3.248966e-11, 3.258496e-11, 3.271165e-11, 3.272461e-11, 
    3.274835e-11, 3.280983e-11, 3.286152e-11, 3.275586e-11, 3.287448e-11, 
    3.242924e-11, 3.266257e-11, 3.229703e-11, 3.24071e-11, 3.24836e-11, 
    3.245004e-11, 3.262431e-11, 3.266539e-11, 3.28323e-11, 3.274601e-11, 
    3.32597e-11, 3.303243e-11, 3.366307e-11, 3.348683e-11, 3.229821e-11, 
    3.235402e-11, 3.254825e-11, 3.245583e-11, 3.272011e-11, 3.278516e-11, 
    3.283804e-11, 3.290564e-11, 3.291294e-11, 3.295299e-11, 3.288736e-11, 
    3.29504e-11, 3.271192e-11, 3.281849e-11, 3.252604e-11, 3.259722e-11, 
    3.256448e-11, 3.252856e-11, 3.263942e-11, 3.275752e-11, 3.276004e-11, 
    3.279791e-11, 3.290464e-11, 3.272118e-11, 3.328905e-11, 3.293835e-11, 
    3.241487e-11, 3.252237e-11, 3.253772e-11, 3.249608e-11, 3.277864e-11, 
    3.267626e-11, 3.295201e-11, 3.287749e-11, 3.29996e-11, 3.293892e-11, 
    3.292999e-11, 3.285206e-11, 3.280354e-11, 3.268095e-11, 3.258121e-11, 
    3.250212e-11, 3.252051e-11, 3.260739e-11, 3.276475e-11, 3.29136e-11, 
    3.288099e-11, 3.299032e-11, 3.270095e-11, 3.282229e-11, 3.277539e-11, 
    3.289767e-11, 3.262973e-11, 3.285791e-11, 3.257141e-11, 3.259653e-11, 
    3.267422e-11, 3.283052e-11, 3.286509e-11, 3.290201e-11, 3.287923e-11, 
    3.276874e-11, 3.275064e-11, 3.267234e-11, 3.265072e-11, 3.259105e-11, 
    3.254166e-11, 3.258679e-11, 3.263419e-11, 3.276878e-11, 3.289008e-11, 
    3.302232e-11, 3.305469e-11, 3.320921e-11, 3.308343e-11, 3.3291e-11, 
    3.311454e-11, 3.342e-11, 3.287113e-11, 3.310933e-11, 3.267776e-11, 
    3.272425e-11, 3.280835e-11, 3.300123e-11, 3.28971e-11, 3.301888e-11, 
    3.274993e-11, 3.261039e-11, 3.257428e-11, 3.250692e-11, 3.257582e-11, 
    3.257022e-11, 3.263615e-11, 3.261496e-11, 3.277325e-11, 3.268823e-11, 
    3.292977e-11, 3.301791e-11, 3.326683e-11, 3.341943e-11, 3.357476e-11, 
    3.364333e-11, 3.366421e-11, 3.367293e-11 ;

 SOILC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 SOILC_HR =
  6.357484e-08, 6.385439e-08, 6.380004e-08, 6.402553e-08, 6.390044e-08, 
    6.404809e-08, 6.363151e-08, 6.386549e-08, 6.371612e-08, 6.360001e-08, 
    6.446311e-08, 6.403558e-08, 6.490716e-08, 6.463451e-08, 6.53194e-08, 
    6.486473e-08, 6.541108e-08, 6.530627e-08, 6.562168e-08, 6.553132e-08, 
    6.593476e-08, 6.566339e-08, 6.614388e-08, 6.586995e-08, 6.59128e-08, 
    6.565443e-08, 6.412161e-08, 6.440989e-08, 6.410453e-08, 6.414565e-08, 
    6.41272e-08, 6.390303e-08, 6.379007e-08, 6.355347e-08, 6.359642e-08, 
    6.377019e-08, 6.416413e-08, 6.40304e-08, 6.436741e-08, 6.43598e-08, 
    6.473498e-08, 6.456582e-08, 6.519642e-08, 6.501719e-08, 6.553509e-08, 
    6.540485e-08, 6.552898e-08, 6.549134e-08, 6.552947e-08, 6.533845e-08, 
    6.542029e-08, 6.52522e-08, 6.459751e-08, 6.478992e-08, 6.421605e-08, 
    6.387099e-08, 6.364178e-08, 6.347913e-08, 6.350213e-08, 6.354596e-08, 
    6.377121e-08, 6.398299e-08, 6.414438e-08, 6.425233e-08, 6.43587e-08, 
    6.46807e-08, 6.48511e-08, 6.523266e-08, 6.516379e-08, 6.528045e-08, 
    6.539189e-08, 6.557899e-08, 6.55482e-08, 6.563063e-08, 6.527737e-08, 
    6.551215e-08, 6.512457e-08, 6.523057e-08, 6.438765e-08, 6.406648e-08, 
    6.392999e-08, 6.38105e-08, 6.351981e-08, 6.372055e-08, 6.364142e-08, 
    6.382967e-08, 6.39493e-08, 6.389013e-08, 6.425529e-08, 6.411333e-08, 
    6.48612e-08, 6.453907e-08, 6.537889e-08, 6.517793e-08, 6.542706e-08, 
    6.529993e-08, 6.551776e-08, 6.532171e-08, 6.566131e-08, 6.573526e-08, 
    6.568472e-08, 6.587883e-08, 6.531085e-08, 6.552898e-08, 6.388848e-08, 
    6.389813e-08, 6.394308e-08, 6.374548e-08, 6.373339e-08, 6.355229e-08, 
    6.371343e-08, 6.378205e-08, 6.395624e-08, 6.405927e-08, 6.415721e-08, 
    6.437256e-08, 6.461306e-08, 6.494936e-08, 6.519095e-08, 6.53529e-08, 
    6.525359e-08, 6.534127e-08, 6.524326e-08, 6.519733e-08, 6.570755e-08, 
    6.542106e-08, 6.585091e-08, 6.582712e-08, 6.563259e-08, 6.582981e-08, 
    6.390491e-08, 6.384938e-08, 6.365659e-08, 6.380746e-08, 6.353257e-08, 
    6.368644e-08, 6.377492e-08, 6.41163e-08, 6.41913e-08, 6.426085e-08, 
    6.43982e-08, 6.457448e-08, 6.488371e-08, 6.515276e-08, 6.539837e-08, 
    6.538038e-08, 6.538671e-08, 6.544158e-08, 6.530567e-08, 6.546389e-08, 
    6.549045e-08, 6.542102e-08, 6.582394e-08, 6.570883e-08, 6.582662e-08, 
    6.575167e-08, 6.386743e-08, 6.396086e-08, 6.391037e-08, 6.400531e-08, 
    6.393843e-08, 6.423585e-08, 6.432501e-08, 6.474225e-08, 6.457101e-08, 
    6.484353e-08, 6.459869e-08, 6.464208e-08, 6.485244e-08, 6.461192e-08, 
    6.513793e-08, 6.478133e-08, 6.544371e-08, 6.508762e-08, 6.546603e-08, 
    6.539731e-08, 6.551109e-08, 6.561299e-08, 6.574118e-08, 6.597772e-08, 
    6.592295e-08, 6.612076e-08, 6.410015e-08, 6.422134e-08, 6.421067e-08, 
    6.433749e-08, 6.443128e-08, 6.463457e-08, 6.496062e-08, 6.483801e-08, 
    6.506309e-08, 6.510828e-08, 6.476632e-08, 6.497628e-08, 6.430245e-08, 
    6.441132e-08, 6.434649e-08, 6.410971e-08, 6.486627e-08, 6.447801e-08, 
    6.519495e-08, 6.498462e-08, 6.559846e-08, 6.529319e-08, 6.589279e-08, 
    6.614913e-08, 6.639036e-08, 6.667229e-08, 6.428748e-08, 6.420513e-08, 
    6.435257e-08, 6.455657e-08, 6.474583e-08, 6.499745e-08, 6.502319e-08, 
    6.507033e-08, 6.519242e-08, 6.529509e-08, 6.508524e-08, 6.532083e-08, 
    6.443658e-08, 6.489997e-08, 6.4174e-08, 6.439262e-08, 6.454454e-08, 
    6.44779e-08, 6.482399e-08, 6.490557e-08, 6.523705e-08, 6.506569e-08, 
    6.608587e-08, 6.563452e-08, 6.688694e-08, 6.653695e-08, 6.417636e-08, 
    6.428719e-08, 6.467292e-08, 6.448939e-08, 6.501424e-08, 6.514343e-08, 
    6.524845e-08, 6.538271e-08, 6.53972e-08, 6.547674e-08, 6.53464e-08, 
    6.547159e-08, 6.499798e-08, 6.520963e-08, 6.462883e-08, 6.47702e-08, 
    6.470516e-08, 6.463382e-08, 6.485399e-08, 6.508855e-08, 6.509355e-08, 
    6.516876e-08, 6.538072e-08, 6.501637e-08, 6.614414e-08, 6.544767e-08, 
    6.440805e-08, 6.462153e-08, 6.465201e-08, 6.456932e-08, 6.513049e-08, 
    6.492716e-08, 6.54748e-08, 6.532679e-08, 6.55693e-08, 6.544879e-08, 
    6.543107e-08, 6.527629e-08, 6.517993e-08, 6.493648e-08, 6.473839e-08, 
    6.458131e-08, 6.461784e-08, 6.479039e-08, 6.51029e-08, 6.539852e-08, 
    6.533376e-08, 6.555087e-08, 6.497619e-08, 6.521717e-08, 6.512403e-08, 
    6.536688e-08, 6.483475e-08, 6.528791e-08, 6.471893e-08, 6.476881e-08, 
    6.492312e-08, 6.523352e-08, 6.530218e-08, 6.53755e-08, 6.533025e-08, 
    6.511083e-08, 6.507487e-08, 6.491937e-08, 6.487644e-08, 6.475795e-08, 
    6.465985e-08, 6.474948e-08, 6.48436e-08, 6.511091e-08, 6.535181e-08, 
    6.561444e-08, 6.567871e-08, 6.598559e-08, 6.573578e-08, 6.614802e-08, 
    6.579756e-08, 6.640422e-08, 6.531416e-08, 6.578724e-08, 6.493014e-08, 
    6.502248e-08, 6.518949e-08, 6.557254e-08, 6.536574e-08, 6.560759e-08, 
    6.507346e-08, 6.479635e-08, 6.472464e-08, 6.459086e-08, 6.472769e-08, 
    6.471657e-08, 6.48475e-08, 6.480542e-08, 6.511979e-08, 6.495092e-08, 
    6.543063e-08, 6.560568e-08, 6.610003e-08, 6.640308e-08, 6.671156e-08, 
    6.684775e-08, 6.68892e-08, 6.690653e-08 ;

 SOILC_LOSS =
  6.357484e-08, 6.385439e-08, 6.380004e-08, 6.402553e-08, 6.390044e-08, 
    6.404809e-08, 6.363151e-08, 6.386549e-08, 6.371612e-08, 6.360001e-08, 
    6.446311e-08, 6.403558e-08, 6.490716e-08, 6.463451e-08, 6.53194e-08, 
    6.486473e-08, 6.541108e-08, 6.530627e-08, 6.562168e-08, 6.553132e-08, 
    6.593476e-08, 6.566339e-08, 6.614388e-08, 6.586995e-08, 6.59128e-08, 
    6.565443e-08, 6.412161e-08, 6.440989e-08, 6.410453e-08, 6.414565e-08, 
    6.41272e-08, 6.390303e-08, 6.379007e-08, 6.355347e-08, 6.359642e-08, 
    6.377019e-08, 6.416413e-08, 6.40304e-08, 6.436741e-08, 6.43598e-08, 
    6.473498e-08, 6.456582e-08, 6.519642e-08, 6.501719e-08, 6.553509e-08, 
    6.540485e-08, 6.552898e-08, 6.549134e-08, 6.552947e-08, 6.533845e-08, 
    6.542029e-08, 6.52522e-08, 6.459751e-08, 6.478992e-08, 6.421605e-08, 
    6.387099e-08, 6.364178e-08, 6.347913e-08, 6.350213e-08, 6.354596e-08, 
    6.377121e-08, 6.398299e-08, 6.414438e-08, 6.425233e-08, 6.43587e-08, 
    6.46807e-08, 6.48511e-08, 6.523266e-08, 6.516379e-08, 6.528045e-08, 
    6.539189e-08, 6.557899e-08, 6.55482e-08, 6.563063e-08, 6.527737e-08, 
    6.551215e-08, 6.512457e-08, 6.523057e-08, 6.438765e-08, 6.406648e-08, 
    6.392999e-08, 6.38105e-08, 6.351981e-08, 6.372055e-08, 6.364142e-08, 
    6.382967e-08, 6.39493e-08, 6.389013e-08, 6.425529e-08, 6.411333e-08, 
    6.48612e-08, 6.453907e-08, 6.537889e-08, 6.517793e-08, 6.542706e-08, 
    6.529993e-08, 6.551776e-08, 6.532171e-08, 6.566131e-08, 6.573526e-08, 
    6.568472e-08, 6.587883e-08, 6.531085e-08, 6.552898e-08, 6.388848e-08, 
    6.389813e-08, 6.394308e-08, 6.374548e-08, 6.373339e-08, 6.355229e-08, 
    6.371343e-08, 6.378205e-08, 6.395624e-08, 6.405927e-08, 6.415721e-08, 
    6.437256e-08, 6.461306e-08, 6.494936e-08, 6.519095e-08, 6.53529e-08, 
    6.525359e-08, 6.534127e-08, 6.524326e-08, 6.519733e-08, 6.570755e-08, 
    6.542106e-08, 6.585091e-08, 6.582712e-08, 6.563259e-08, 6.582981e-08, 
    6.390491e-08, 6.384938e-08, 6.365659e-08, 6.380746e-08, 6.353257e-08, 
    6.368644e-08, 6.377492e-08, 6.41163e-08, 6.41913e-08, 6.426085e-08, 
    6.43982e-08, 6.457448e-08, 6.488371e-08, 6.515276e-08, 6.539837e-08, 
    6.538038e-08, 6.538671e-08, 6.544158e-08, 6.530567e-08, 6.546389e-08, 
    6.549045e-08, 6.542102e-08, 6.582394e-08, 6.570883e-08, 6.582662e-08, 
    6.575167e-08, 6.386743e-08, 6.396086e-08, 6.391037e-08, 6.400531e-08, 
    6.393843e-08, 6.423585e-08, 6.432501e-08, 6.474225e-08, 6.457101e-08, 
    6.484353e-08, 6.459869e-08, 6.464208e-08, 6.485244e-08, 6.461192e-08, 
    6.513793e-08, 6.478133e-08, 6.544371e-08, 6.508762e-08, 6.546603e-08, 
    6.539731e-08, 6.551109e-08, 6.561299e-08, 6.574118e-08, 6.597772e-08, 
    6.592295e-08, 6.612076e-08, 6.410015e-08, 6.422134e-08, 6.421067e-08, 
    6.433749e-08, 6.443128e-08, 6.463457e-08, 6.496062e-08, 6.483801e-08, 
    6.506309e-08, 6.510828e-08, 6.476632e-08, 6.497628e-08, 6.430245e-08, 
    6.441132e-08, 6.434649e-08, 6.410971e-08, 6.486627e-08, 6.447801e-08, 
    6.519495e-08, 6.498462e-08, 6.559846e-08, 6.529319e-08, 6.589279e-08, 
    6.614913e-08, 6.639036e-08, 6.667229e-08, 6.428748e-08, 6.420513e-08, 
    6.435257e-08, 6.455657e-08, 6.474583e-08, 6.499745e-08, 6.502319e-08, 
    6.507033e-08, 6.519242e-08, 6.529509e-08, 6.508524e-08, 6.532083e-08, 
    6.443658e-08, 6.489997e-08, 6.4174e-08, 6.439262e-08, 6.454454e-08, 
    6.44779e-08, 6.482399e-08, 6.490557e-08, 6.523705e-08, 6.506569e-08, 
    6.608587e-08, 6.563452e-08, 6.688694e-08, 6.653695e-08, 6.417636e-08, 
    6.428719e-08, 6.467292e-08, 6.448939e-08, 6.501424e-08, 6.514343e-08, 
    6.524845e-08, 6.538271e-08, 6.53972e-08, 6.547674e-08, 6.53464e-08, 
    6.547159e-08, 6.499798e-08, 6.520963e-08, 6.462883e-08, 6.47702e-08, 
    6.470516e-08, 6.463382e-08, 6.485399e-08, 6.508855e-08, 6.509355e-08, 
    6.516876e-08, 6.538072e-08, 6.501637e-08, 6.614414e-08, 6.544767e-08, 
    6.440805e-08, 6.462153e-08, 6.465201e-08, 6.456932e-08, 6.513049e-08, 
    6.492716e-08, 6.54748e-08, 6.532679e-08, 6.55693e-08, 6.544879e-08, 
    6.543107e-08, 6.527629e-08, 6.517993e-08, 6.493648e-08, 6.473839e-08, 
    6.458131e-08, 6.461784e-08, 6.479039e-08, 6.51029e-08, 6.539852e-08, 
    6.533376e-08, 6.555087e-08, 6.497619e-08, 6.521717e-08, 6.512403e-08, 
    6.536688e-08, 6.483475e-08, 6.528791e-08, 6.471893e-08, 6.476881e-08, 
    6.492312e-08, 6.523352e-08, 6.530218e-08, 6.53755e-08, 6.533025e-08, 
    6.511083e-08, 6.507487e-08, 6.491937e-08, 6.487644e-08, 6.475795e-08, 
    6.465985e-08, 6.474948e-08, 6.48436e-08, 6.511091e-08, 6.535181e-08, 
    6.561444e-08, 6.567871e-08, 6.598559e-08, 6.573578e-08, 6.614802e-08, 
    6.579756e-08, 6.640422e-08, 6.531416e-08, 6.578724e-08, 6.493014e-08, 
    6.502248e-08, 6.518949e-08, 6.557254e-08, 6.536574e-08, 6.560759e-08, 
    6.507346e-08, 6.479635e-08, 6.472464e-08, 6.459086e-08, 6.472769e-08, 
    6.471657e-08, 6.48475e-08, 6.480542e-08, 6.511979e-08, 6.495092e-08, 
    6.543063e-08, 6.560568e-08, 6.610003e-08, 6.640308e-08, 6.671156e-08, 
    6.684775e-08, 6.68892e-08, 6.690653e-08 ;

 SOILICE =
  56.63643, 56.82955, 56.79198, 56.94802, 56.86144, 56.96366, 56.67557, 
    56.8372, 56.73399, 56.65384, 57.25174, 56.95499, 57.56158, 57.37131, 
    57.85032, 57.5319, 57.9147, 57.84118, 58.06285, 57.99929, 58.28341, 
    58.09222, 58.43122, 58.23774, 58.26795, 58.08591, 57.01468, 57.21471, 
    57.00283, 57.03131, 57.01854, 56.86321, 56.78502, 56.62174, 56.65137, 
    56.77132, 57.04413, 56.95145, 57.18539, 57.1801, 57.4414, 57.32347, 
    57.76413, 57.63863, 58.00194, 57.91039, 57.99762, 57.97117, 57.99797, 
    57.86375, 57.92123, 57.80325, 57.34553, 57.47972, 57.08019, 56.84094, 
    56.68264, 56.57048, 56.58633, 56.61653, 56.77203, 56.9186, 57.03049, 
    57.10542, 57.17934, 57.40339, 57.52241, 57.7895, 57.74128, 57.82303, 
    57.90129, 58.0328, 58.01115, 58.06913, 57.82092, 57.98576, 57.71382, 
    57.78809, 57.19923, 56.97645, 56.88178, 56.79919, 56.59851, 56.73702, 
    56.68238, 56.8125, 56.89527, 56.85433, 57.10747, 57.00894, 57.52947, 
    57.30479, 57.89216, 57.75118, 57.926, 57.83675, 57.98972, 57.85204, 
    58.09074, 58.14279, 58.10721, 58.24405, 57.84441, 57.9976, 56.85317, 
    56.85984, 56.89097, 56.75424, 56.7459, 56.62092, 56.73214, 56.77953, 
    56.90009, 56.97145, 57.03938, 57.18895, 57.35634, 57.59113, 57.76031, 
    57.87393, 57.80425, 57.86576, 57.797, 57.7648, 58.12326, 57.92175, 
    58.22435, 58.20758, 58.0705, 58.20947, 56.86454, 56.82613, 56.69287, 
    56.79713, 56.60732, 56.71348, 56.77457, 57.01095, 57.06304, 57.11131, 
    57.20679, 57.3295, 57.54524, 57.73352, 57.90586, 57.89322, 57.89767, 
    57.9362, 57.84077, 57.95187, 57.97052, 57.92175, 58.20534, 58.12421, 
    58.20723, 58.1544, 56.83862, 56.90327, 56.86832, 56.93405, 56.88772, 
    57.09389, 57.15583, 57.44641, 57.32707, 57.51716, 57.34637, 57.37659, 
    57.52328, 57.35561, 57.72309, 57.47366, 57.93769, 57.68779, 57.95338, 
    57.90511, 57.98506, 58.05671, 58.147, 58.31381, 58.27516, 58.41491, 
    56.9998, 57.08385, 57.07649, 57.16458, 57.22979, 57.37139, 57.59903, 
    57.51336, 57.67076, 57.70238, 57.4633, 57.60996, 57.1402, 57.21584, 
    57.17082, 57.0064, 57.53303, 57.26225, 57.7631, 57.61583, 58.04649, 
    57.83195, 58.25388, 58.43487, 58.6058, 58.80582, 57.12982, 57.07265, 
    57.17508, 57.31696, 57.44897, 57.62479, 57.64283, 57.67581, 57.76136, 
    57.83335, 57.6862, 57.85141, 57.23331, 57.5566, 57.05101, 57.20282, 
    57.30861, 57.26223, 57.50358, 57.56057, 57.79259, 57.67258, 58.39013, 
    58.0718, 58.9586, 58.70971, 57.05268, 57.12964, 57.39808, 57.27024, 
    57.63657, 57.72701, 57.80065, 57.89482, 57.90503, 57.96089, 57.86936, 
    57.95729, 57.62517, 57.77341, 57.3674, 57.46598, 57.42063, 57.37088, 
    57.52452, 57.6885, 57.69208, 57.74473, 57.89318, 57.63806, 58.43119, 
    57.94025, 57.21365, 57.36221, 57.38354, 57.32592, 57.71793, 57.57564, 
    57.95954, 57.8556, 58.026, 57.94127, 57.92881, 57.82016, 57.75258, 
    57.58214, 57.44378, 57.33429, 57.35973, 57.48006, 57.69856, 57.90592, 
    57.86044, 58.01303, 57.60994, 57.77866, 57.71338, 57.88373, 57.51107, 
    57.82809, 57.43023, 57.46504, 57.57281, 57.79007, 57.83833, 57.88976, 
    57.85803, 57.70413, 57.67898, 57.57021, 57.54018, 57.45747, 57.38903, 
    57.45153, 57.51723, 57.70422, 57.87312, 58.05772, 58.103, 58.31924, 
    58.14307, 58.43392, 58.18644, 58.61543, 57.8466, 58.1793, 57.57775, 
    57.64233, 57.75922, 58.02818, 57.88293, 58.05286, 57.678, 57.48419, 
    57.43421, 57.34092, 57.43634, 57.42858, 57.52, 57.49061, 57.71044, 
    57.59228, 57.92848, 58.05153, 58.40023, 58.61475, 58.83384, 58.93073, 
    58.96024, 58.97258,
  78.20255, 78.50357, 78.44503, 78.68825, 78.55334, 78.71265, 78.2636, 
    78.51546, 78.35465, 78.22973, 79.15324, 78.69914, 79.62355, 79.33496, 
    80.06183, 79.57845, 80.15962, 80.04809, 80.38474, 80.28819, 80.71954, 
    80.42934, 80.94425, 80.65029, 80.69613, 80.41974, 78.79225, 79.09707, 
    78.77377, 78.81816, 78.79828, 78.55605, 78.43407, 78.17972, 78.22588, 
    78.4128, 78.83813, 78.69367, 79.05303, 79.04501, 79.44131, 79.26243, 
    79.93111, 79.74065, 80.29222, 80.15319, 80.28565, 80.2455, 80.28617, 
    80.08235, 80.16961, 79.99052, 79.29585, 79.49943, 78.89341, 78.52119, 
    78.27459, 78.09982, 78.12451, 78.17155, 78.41389, 78.64246, 78.81694, 
    78.93174, 79.04385, 79.3834, 79.56411, 79.96955, 79.89646, 80.02047, 
    80.13937, 80.33905, 80.30619, 80.39421, 80.01734, 80.26758, 79.8548, 
    79.9675, 79.07357, 78.73266, 78.58489, 78.45626, 78.14349, 78.35933, 
    78.27417, 78.47704, 78.60608, 78.54227, 78.93485, 78.78333, 79.57483, 
    79.23403, 80.1255, 79.91148, 80.1769, 80.0414, 80.27361, 80.06461, 
    80.42706, 80.50607, 80.45205, 80.65996, 80.05302, 80.28558, 78.54045, 
    78.55084, 78.59939, 78.38617, 78.37318, 78.17841, 78.35175, 78.42561, 
    78.61362, 78.72486, 78.83077, 79.05838, 79.31219, 79.66845, 79.92532, 
    80.09785, 79.99207, 80.08544, 79.98104, 79.93218, 80.4764, 80.17039, 
    80.63003, 80.60457, 80.39628, 80.60744, 78.55816, 78.49831, 78.29055, 
    78.4531, 78.15724, 78.32265, 78.41784, 78.78638, 78.86748, 78.94064, 
    79.08547, 79.27157, 79.59885, 79.88461, 80.14633, 80.12714, 80.13389, 
    80.19236, 80.04749, 80.21617, 80.24444, 80.17044, 80.60115, 80.47792, 
    80.60403, 80.52379, 78.51778, 78.61856, 78.56408, 78.66653, 78.59428, 
    78.91412, 79.00802, 79.4488, 79.26786, 79.55621, 79.29717, 79.34297, 
    79.56529, 79.3112, 79.86868, 79.49009, 80.19463, 79.81501, 80.21845, 
    80.1452, 80.2666, 80.37537, 80.51253, 80.76586, 80.70718, 80.91953, 
    78.76908, 78.89896, 78.88788, 79.02145, 79.12032, 79.33514, 79.6805, 
    79.55053, 79.78942, 79.8374, 79.4746, 79.69706, 78.98441, 79.09904, 
    79.03088, 78.77934, 79.58026, 79.16945, 79.92954, 79.70602, 80.35983, 
    80.03399, 80.67485, 80.94968, 81.20969, 81.5136, 78.9687, 78.88206, 
    79.03739, 79.25243, 79.45281, 79.7196, 79.74702, 79.79706, 79.92696, 
    80.03623, 79.81274, 80.06366, 79.12536, 79.61607, 78.84891, 79.07928, 
    79.23981, 79.1695, 79.53573, 79.62218, 79.97427, 79.7922, 80.88165, 
    80.39816, 81.74607, 81.36751, 78.85155, 78.96848, 79.37554, 79.18167, 
    79.73752, 79.87476, 79.9866, 80.1295, 80.14505, 80.22985, 80.09091, 
    80.22441, 79.72018, 79.94521, 79.3291, 79.47861, 79.40986, 79.33438, 
    79.5675, 79.81622, 79.82178, 79.90163, 80.12657, 79.73979, 80.94378, 
    80.1981, 79.09589, 79.32105, 79.35355, 79.26618, 79.86098, 79.64502, 
    80.22781, 80.07001, 80.32876, 80.20008, 80.18115, 80.01621, 79.9136, 
    79.65487, 79.44492, 79.27888, 79.31747, 79.49996, 79.83151, 80.14635, 
    80.07727, 80.30907, 79.69711, 79.95313, 79.85402, 80.1127, 79.54704, 
    80.02781, 79.42443, 79.47723, 79.64074, 79.97036, 80.04379, 80.12182, 
    80.07371, 79.83999, 79.80185, 79.63682, 79.59119, 79.46575, 79.36192, 
    79.45673, 79.55634, 79.84018, 80.09654, 80.37688, 80.44571, 80.77389, 
    80.50633, 80.9479, 80.57188, 81.22393, 80.0561, 80.5613, 79.64826, 
    79.74628, 79.92357, 80.33188, 80.11149, 80.3694, 79.80038, 79.50615, 
    79.43046, 79.28892, 79.4337, 79.42193, 79.56063, 79.51605, 79.84962, 
    79.67031, 80.18061, 80.36742, 80.89716, 81.22313, 81.55639, 81.70374, 
    81.74864, 81.76741,
  118.5275, 119.0841, 118.9757, 119.4257, 119.176, 119.4708, 118.6402, 
    119.1062, 118.8086, 118.5776, 120.3024, 119.4458, 121.1971, 120.6473, 
    122.032, 121.1114, 122.2144, 122.0054, 122.6291, 122.4511, 123.2473, 
    122.7114, 123.6616, 123.1192, 123.2039, 122.6937, 119.6179, 120.1955, 
    119.5837, 119.6659, 119.629, 119.1811, 118.9558, 118.4851, 118.5705, 
    118.9162, 119.7029, 119.4355, 120.1104, 120.0951, 120.8497, 120.5091, 
    121.7825, 121.4196, 122.4585, 122.2023, 122.4465, 122.3724, 122.4474, 
    122.0707, 122.2326, 121.8957, 120.5728, 120.9605, 119.8069, 119.1171, 
    118.6606, 118.3375, 118.3831, 118.4702, 118.9183, 119.3408, 119.6634, 
    119.8796, 120.0929, 120.7402, 121.0839, 121.856, 121.7164, 121.953, 
    122.1768, 122.545, 122.4843, 122.6468, 121.9467, 122.4133, 121.637, 
    121.8518, 120.1509, 119.5076, 119.2348, 118.9966, 118.4182, 118.8174, 
    118.6599, 119.0348, 119.2735, 119.1554, 119.8856, 119.6013, 121.1043, 
    120.4552, 122.1512, 121.7451, 122.2459, 121.9925, 122.4244, 122.0368, 
    122.7073, 122.8531, 122.7534, 123.1368, 122.0147, 122.4465, 119.1521, 
    119.1713, 119.2611, 118.867, 118.8429, 118.4828, 118.8032, 118.9399, 
    119.2873, 119.4932, 119.6891, 120.1207, 120.6041, 121.2824, 121.7715, 
    122.1001, 121.8985, 122.0764, 121.8775, 121.7844, 122.7984, 122.2341, 
    123.0816, 123.0346, 122.6506, 123.0399, 119.1849, 119.0741, 118.6901, 
    118.9905, 118.4436, 118.7495, 118.9257, 119.6072, 119.7574, 119.8967, 
    120.1722, 120.5265, 121.1498, 121.6941, 122.1895, 122.1542, 122.1666, 
    122.2745, 122.0042, 122.3184, 122.3706, 122.2341, 123.0283, 122.801, 
    123.0336, 122.8856, 119.1101, 119.2966, 119.1958, 119.3853, 119.2518, 
    119.8465, 120.0253, 120.8643, 120.5195, 121.0687, 120.5752, 120.6625, 
    121.0866, 120.6019, 121.664, 120.9431, 122.2787, 121.562, 122.3226, 
    122.1874, 122.4113, 122.612, 122.8648, 123.3324, 123.224, 123.6158, 
    119.5749, 119.8175, 119.7962, 120.0504, 120.2386, 120.6474, 121.3052, 
    121.0576, 121.5125, 121.604, 120.9129, 121.3369, 119.9801, 120.1985, 
    120.0684, 119.5941, 121.1146, 120.3325, 121.7796, 121.3537, 122.5833, 
    121.9788, 123.1644, 123.672, 124.1513, 124.713, 119.9501, 119.7851, 
    120.0806, 120.4904, 120.8716, 121.3797, 121.4318, 121.5271, 121.7745, 
    121.9827, 121.5573, 122.0349, 120.2492, 121.1826, 119.7227, 120.1609, 
    120.4662, 120.3323, 121.0293, 121.194, 121.8649, 121.5178, 123.5465, 
    122.6544, 125.142, 124.4431, 119.7275, 119.9495, 120.7247, 120.3554, 
    121.4137, 121.6752, 121.8881, 122.1587, 122.1872, 122.3437, 122.0869, 
    122.3335, 121.3808, 121.8093, 120.6359, 120.9207, 120.7896, 120.646, 
    121.0898, 121.564, 121.5741, 121.7265, 122.1546, 121.418, 123.662, 
    122.2863, 120.192, 120.6211, 120.6826, 120.5161, 121.6489, 121.2376, 
    122.3399, 122.0471, 122.5259, 122.2887, 122.2538, 121.9445, 121.7491, 
    121.2564, 120.8566, 120.5403, 120.6138, 120.9614, 121.593, 122.1898, 
    122.0612, 122.4896, 121.3367, 121.8246, 121.6358, 122.1276, 121.051, 
    121.968, 120.8174, 120.9179, 121.2294, 121.8577, 121.9971, 122.1446, 
    122.0541, 121.6091, 121.5363, 121.2219, 121.1351, 120.896, 120.6984, 
    120.879, 121.0688, 121.6093, 122.0978, 122.6148, 122.7416, 123.3479, 
    122.8541, 123.6696, 122.9759, 124.1787, 122.0213, 122.9557, 121.2436, 
    121.4303, 121.7685, 122.5322, 122.1254, 122.6013, 121.5335, 120.9734, 
    120.8289, 120.5595, 120.8351, 120.8126, 121.0767, 120.9918, 121.6273, 
    121.2856, 122.2529, 122.5975, 123.5747, 124.1765, 124.7915, 125.0636, 
    125.1466, 125.1812,
  187.3257, 188.3278, 188.1326, 188.9433, 188.4932, 189.0245, 187.5285, 
    188.3677, 187.8316, 187.4157, 190.5242, 188.9795, 192.1386, 191.146, 
    193.6468, 191.9839, 193.9758, 193.5986, 194.7247, 194.4031, 195.8423, 
    194.8732, 196.5915, 195.6105, 195.7637, 194.8413, 189.2895, 190.3314, 
    189.2279, 189.3762, 189.3096, 188.5025, 188.0969, 187.2492, 187.4029, 
    188.0255, 189.4429, 188.9608, 190.1774, 190.1499, 191.5113, 190.8965, 
    193.1959, 192.5402, 194.4165, 193.9536, 194.3947, 194.2609, 194.3965, 
    193.7167, 194.0085, 193.4003, 191.0116, 191.7113, 189.6303, 188.3875, 
    187.5652, 186.9835, 187.0657, 187.2224, 188.0292, 188.7901, 189.3716, 
    189.7613, 190.1459, 191.3139, 191.9342, 193.3287, 193.0764, 193.5039, 
    193.9076, 194.5727, 194.4631, 194.7565, 193.4926, 194.3349, 192.9328, 
    193.321, 190.2509, 189.0907, 188.5995, 188.1701, 187.1288, 187.8475, 
    187.5639, 188.239, 188.6689, 188.4562, 189.772, 189.2596, 191.971, 
    190.7995, 193.8615, 193.1281, 194.0325, 193.5753, 194.3548, 193.6552, 
    194.8658, 195.1295, 194.9493, 195.6422, 193.6154, 194.3947, 188.4502, 
    188.4849, 188.6465, 187.9369, 187.8935, 187.245, 187.8219, 188.068, 
    188.6938, 189.0648, 189.4179, 190.1961, 191.0681, 192.2925, 193.1759, 
    193.7693, 193.4054, 193.727, 193.3675, 193.1992, 195.0307, 194.0112, 
    195.5424, 195.4574, 194.7635, 195.467, 188.5093, 188.3097, 187.6183, 
    188.1592, 187.1745, 187.7252, 188.0425, 189.2704, 189.5409, 189.7921, 
    190.2889, 190.928, 192.0531, 193.036, 193.9306, 193.8668, 193.8893, 
    194.0841, 193.5964, 194.1634, 194.2578, 194.011, 195.446, 195.0352, 
    195.4556, 195.188, 188.3746, 188.7105, 188.5289, 188.8705, 188.6298, 
    189.7018, 190.0241, 191.5378, 190.9154, 191.9066, 191.0159, 191.1735, 
    191.9391, 191.0639, 192.9818, 191.68, 194.0917, 192.7977, 194.1709, 
    193.9269, 194.3311, 194.6937, 195.1506, 195.996, 195.7999, 196.5085, 
    189.2121, 189.6494, 189.6108, 190.0692, 190.4087, 191.1462, 192.3336, 
    191.8864, 192.708, 192.8732, 191.6253, 192.3908, 189.9425, 190.3365, 
    190.1018, 189.2466, 191.9895, 190.5781, 193.1905, 192.4212, 194.642, 
    193.5506, 195.6921, 196.6104, 197.4775, 198.4949, 189.8883, 189.5908, 
    190.1237, 190.863, 191.5508, 192.4681, 192.5621, 192.7344, 193.1812, 
    193.5575, 192.789, 193.652, 190.428, 192.1123, 189.4785, 190.2688, 
    190.8194, 190.5776, 191.8353, 192.1327, 193.3448, 192.7175, 196.3835, 
    194.7704, 199.2722, 198.006, 189.487, 189.8873, 191.2856, 190.6193, 
    192.5294, 193.0019, 193.3865, 193.8751, 193.9265, 194.209, 193.7458, 
    194.1907, 192.4701, 193.2443, 191.1253, 191.6395, 191.4028, 191.1435, 
    191.9446, 192.8011, 192.8193, 193.0946, 193.8682, 192.5372, 196.5926, 
    194.1059, 190.3245, 191.0989, 191.2096, 190.9092, 192.9545, 192.2115, 
    194.2021, 193.6739, 194.5382, 194.1097, 194.0467, 193.4886, 193.1355, 
    192.2455, 191.5237, 190.9528, 191.0854, 191.713, 192.8535, 193.9312, 
    193.6995, 194.4726, 192.3905, 193.2719, 192.9309, 193.8189, 191.8746, 
    193.5314, 191.4528, 191.6344, 192.1968, 193.3319, 193.5836, 193.8495, 
    193.6866, 192.8826, 192.751, 192.1831, 192.0265, 191.5948, 191.2381, 
    191.564, 191.9068, 192.8829, 193.7654, 194.6989, 194.9278, 196.0242, 
    195.1315, 196.6065, 195.352, 197.5275, 193.6276, 195.3151, 192.2224, 
    192.5595, 193.1705, 194.5498, 193.8148, 194.6745, 192.7459, 191.7347, 
    191.4736, 190.9875, 191.4848, 191.4443, 191.921, 191.7677, 192.9153, 
    192.2982, 194.0452, 194.6677, 196.4342, 197.5234, 198.6369, 199.1301, 
    199.2803, 199.3432,
  314.8268, 316.5648, 316.2262, 317.6333, 316.8519, 317.7745, 315.1783, 
    316.634, 315.7039, 314.9827, 320.3815, 317.6962, 323.1932, 321.4637, 
    325.825, 322.9236, 326.413, 325.7408, 327.7678, 327.1858, 329.7831, 
    328.0367, 331.0963, 329.372, 329.6455, 327.9789, 318.2347, 320.0461, 
    318.1277, 318.3853, 318.2697, 316.8681, 316.1642, 314.6942, 314.9605, 
    316.0404, 318.5013, 317.6637, 319.7782, 319.7303, 322.1, 321.0295, 
    325.0376, 323.8935, 327.2101, 326.3729, 327.1707, 326.9286, 327.1739, 
    325.947, 326.4721, 325.3944, 321.2297, 322.4484, 318.8269, 316.6684, 
    315.242, 314.2337, 314.3761, 314.6477, 316.0467, 317.3673, 318.3773, 
    319.0547, 319.7234, 321.7563, 322.8369, 325.2695, 324.829, 325.5754, 
    326.2898, 327.4927, 327.2944, 327.8255, 325.5556, 327.0625, 324.5784, 
    325.256, 319.9061, 317.8894, 317.0365, 316.2913, 314.4856, 315.7315, 
    315.2398, 316.4107, 317.1569, 316.7876, 319.0732, 318.1828, 322.9011, 
    320.8606, 326.2064, 324.9194, 326.5156, 325.7001, 327.0986, 325.8397, 
    328.0233, 328.5008, 328.1744, 329.4295, 325.7701, 327.1708, 316.7773, 
    316.8375, 317.118, 315.8866, 315.8113, 314.6869, 315.6872, 316.1141, 
    317.2002, 317.8444, 318.4578, 319.8107, 321.3282, 323.4616, 325.0027, 
    326.0396, 325.4034, 325.965, 325.3372, 325.0433, 328.3218, 326.4771, 
    329.2487, 329.0947, 327.8382, 329.112, 316.8798, 316.5334, 315.334, 
    316.2723, 314.5647, 315.5195, 316.0698, 318.2015, 318.6715, 319.1082, 
    319.9721, 321.0842, 323.0441, 324.7586, 326.3314, 326.2159, 326.2565, 
    326.6088, 325.7368, 326.7522, 326.923, 326.4767, 329.0741, 328.33, 
    329.0914, 328.6067, 316.646, 317.2291, 316.9139, 317.5069, 317.0891, 
    318.9513, 319.5117, 322.1462, 321.0623, 322.7888, 321.2372, 321.5117, 
    322.8456, 321.3209, 324.664, 322.394, 326.6225, 324.3428, 326.7659, 
    326.3245, 327.0556, 327.7118, 328.5389, 330.0524, 329.709, 330.9507, 
    318.1003, 318.8602, 318.7931, 319.59, 320.1806, 321.4641, 323.5332, 
    322.7536, 324.1861, 324.4745, 322.2986, 323.633, 319.3696, 320.0549, 
    319.6466, 318.1602, 322.9333, 320.4753, 325.0282, 323.686, 327.6181, 
    325.657, 329.52, 331.1294, 332.6507, 334.4381, 319.2755, 318.7584, 
    319.6848, 320.9711, 322.1688, 323.7678, 323.9317, 324.2323, 325.012, 
    325.6691, 324.3275, 325.834, 320.2142, 323.1474, 318.5631, 319.9371, 
    320.8951, 320.4744, 322.6646, 323.1829, 325.2975, 324.2027, 330.7316, 
    327.8507, 335.8051, 333.5789, 318.5779, 319.2737, 321.7069, 320.547, 
    323.8747, 324.699, 325.3704, 326.2309, 326.3238, 326.8348, 325.9979, 
    326.8017, 323.7712, 325.122, 321.4278, 322.3232, 321.9109, 321.4594, 
    322.8551, 324.3486, 324.3804, 324.8608, 326.2186, 323.8882, 331.0983, 
    326.6484, 320.0341, 321.3818, 321.5745, 321.0515, 324.6162, 323.3203, 
    326.8223, 325.8722, 327.4303, 326.6552, 326.5413, 325.5486, 324.9322, 
    323.3796, 322.1216, 321.1273, 321.3582, 322.4514, 324.4402, 326.3323, 
    325.917, 327.3116, 323.6323, 325.1703, 324.5751, 326.1293, 322.733, 
    325.6235, 321.9981, 322.3144, 323.2946, 325.275, 325.7145, 326.1847, 
    325.8944, 324.4908, 324.2613, 323.2707, 322.9978, 322.2455, 321.6241, 
    322.1919, 322.7892, 324.4913, 326.0327, 327.7211, 328.1356, 330.102, 
    328.5043, 331.1227, 328.904, 332.7387, 325.7915, 328.8369, 323.3392, 
    323.9272, 324.9934, 327.4514, 326.122, 327.6771, 324.2523, 322.4893, 
    322.0344, 321.1877, 322.0537, 321.9832, 322.8139, 322.5467, 324.5479, 
    323.4715, 326.5385, 327.6647, 330.8204, 332.7313, 334.6876, 335.5551, 
    335.8195, 335.9301,
  523.2241, 526.4968, 525.8586, 528.5126, 527.0382, 528.7791, 523.8855, 
    526.6274, 524.8749, 523.5176, 533.7101, 528.6313, 539.0477, 535.7622, 
    544.0626, 538.535, 545.1855, 543.9018, 547.7762, 546.6628, 551.6569, 
    548.2911, 554.2677, 550.8506, 551.3835, 548.1806, 529.6483, 533.0747, 
    529.4462, 529.9329, 529.7144, 527.0687, 525.7418, 522.9748, 523.4758, 
    525.5085, 530.152, 528.5699, 532.5674, 532.4767, 536.97, 534.9384, 
    542.5602, 540.3803, 546.7092, 545.1089, 546.6339, 546.1709, 546.64, 
    544.2954, 545.2984, 543.2408, 535.3182, 537.6318, 530.7676, 526.6922, 
    524.0054, 522.1092, 522.3768, 522.8874, 525.5205, 528.0105, 529.9178, 
    531.1983, 532.4637, 536.3174, 538.3702, 543.0025, 542.1626, 543.5862, 
    544.9501, 547.2499, 546.8705, 547.8868, 543.5483, 546.427, 541.6849, 
    542.9769, 532.8096, 528.9962, 527.3863, 525.9813, 522.5826, 524.9269, 
    524.0013, 526.2064, 527.6135, 526.9169, 531.2334, 529.5502, 538.4922, 
    534.618, 544.7908, 542.3348, 545.3814, 543.8241, 546.496, 544.0906, 
    548.2656, 549.1801, 548.5549, 550.9608, 543.9576, 546.634, 526.8975, 
    527.011, 527.5402, 525.2189, 525.0772, 522.9611, 524.8434, 525.6475, 
    527.6951, 528.911, 530.0699, 532.6289, 535.5049, 539.5583, 542.4936, 
    544.4724, 543.2579, 544.3299, 543.1317, 542.5712, 548.8373, 545.3079, 
    550.614, 550.3186, 547.9111, 550.3519, 527.0907, 526.4377, 524.1785, 
    525.9455, 522.7313, 524.5276, 525.564, 529.5856, 530.4739, 531.2996, 
    532.9346, 535.0421, 538.7641, 542.0284, 545.0295, 544.8089, 544.8865, 
    545.5597, 543.8943, 545.8337, 546.1602, 545.3073, 550.2791, 548.8529, 
    550.3124, 549.3831, 526.6498, 527.7496, 527.155, 528.2739, 527.4854, 
    531.0027, 532.0629, 537.0577, 535.0006, 538.2788, 535.3324, 535.8531, 
    538.3867, 535.491, 541.848, 537.5286, 545.5859, 541.2361, 545.8599, 
    545.0165, 546.4138, 547.6691, 549.2533, 552.1918, 551.5095, 553.9781, 
    529.3943, 530.8305, 530.7036, 532.2111, 533.3294, 535.7629, 539.6946, 
    538.2119, 540.9376, 541.4869, 537.3472, 539.8845, 531.7941, 533.0914, 
    532.3184, 529.5076, 538.5534, 533.8878, 542.5424, 539.9854, 547.4899, 
    543.7419, 551.1345, 554.3337, 557.2769, 560.7277, 531.6161, 530.6379, 
    532.3907, 534.8278, 537.1006, 540.141, 540.4531, 541.0256, 542.5115, 
    543.7649, 541.2069, 544.0797, 533.3932, 538.9606, 530.2689, 532.8683, 
    534.6836, 533.8861, 538.0427, 539.0282, 543.0561, 540.9691, 553.5422, 
    547.9351, 563.3732, 559.0677, 530.2968, 531.6126, 536.2237, 534.0236, 
    540.3445, 541.9147, 543.1951, 544.8376, 545.0151, 545.9916, 544.3926, 
    545.9283, 540.1475, 542.7213, 535.6938, 537.394, 536.611, 535.7538, 
    538.4047, 541.2471, 541.3077, 542.2232, 544.8141, 540.3704, 554.2719, 
    545.6354, 533.052, 535.6067, 535.9724, 534.9802, 541.757, 539.2894, 
    545.9677, 544.1527, 547.1304, 545.6483, 545.4306, 543.5351, 542.3593, 
    539.4023, 537.011, 535.1239, 535.562, 537.6375, 541.4215, 545.0314, 
    544.2382, 546.9034, 539.8832, 542.8134, 541.6786, 544.6436, 538.1726, 
    543.6781, 536.7766, 537.3773, 539.2406, 543.0131, 543.8516, 544.7493, 
    544.1951, 541.5179, 541.0807, 539.1951, 538.6761, 537.2464, 536.0664, 
    537.1445, 538.2796, 541.5189, 544.459, 547.6871, 548.4805, 552.2903, 
    549.187, 554.3205, 549.9531, 557.4465, 543.9987, 549.8245, 539.3254, 
    540.4444, 542.476, 547.1708, 544.6296, 547.6027, 541.0636, 537.7095, 
    536.8453, 535.2385, 536.8821, 536.7482, 538.3264, 537.8186, 541.6269, 
    539.5771, 545.4252, 547.5791, 553.7189, 557.4323, 561.2101, 562.8888, 
    563.4011, 563.6154,
  947.1252, 953.998, 952.6549, 958.2488, 955.1384, 958.8117, 948.5112, 
    954.2729, 950.5876, 947.7399, 969.1228, 958.4996, 980.1627, 973.3557, 
    990.624, 979.098, 992.9788, 990.2872, 998.4282, 996.0831, 1006.636, 
    999.5141, 1012.19, 1004.926, 1006.056, 999.2809, 960.6497, 967.8149, 
    960.2222, 961.2521, 960.7896, 955.2027, 952.4093, 946.603, 947.6523, 
    951.9189, 961.7158, 958.3699, 966.7717, 966.5853, 975.8538, 971.6547, 
    987.4808, 982.934, 996.1807, 992.818, 996.0224, 995.0486, 996.0351, 
    991.1119, 993.2156, 988.9039, 972.4387, 977.2248, 963.0202, 954.4094, 
    948.7628, 944.7917, 945.3513, 946.4199, 951.944, 957.1887, 961.22, 
    963.9335, 966.5585, 974.5035, 978.756, 988.4053, 986.6502, 989.6265, 
    992.4846, 997.3192, 996.5203, 998.6613, 989.5472, 995.5871, 985.6532, 
    988.3517, 967.2695, 959.2704, 955.8721, 952.9129, 945.782, 950.6966, 
    948.754, 953.3865, 956.3511, 954.8827, 964.0079, 960.4421, 979.0092, 
    970.9939, 992.1505, 987.0099, 993.39, 990.1246, 995.7322, 990.6827, 
    999.4601, 1001.391, 1000.071, 1005.16, 990.4042, 996.0226, 954.8417, 
    955.0809, 956.1965, 951.31, 951.0124, 946.5743, 950.5213, 952.211, 
    956.5232, 959.0905, 961.5421, 966.8981, 972.8243, 981.2239, 987.3416, 
    991.4827, 988.9394, 991.1841, 988.6755, 987.5037, 1000.667, 993.2355, 
    1004.425, 1003.799, 998.7124, 1003.87, 955.2489, 953.8735, 949.1257, 
    952.8378, 946.0931, 949.8585, 952.0355, 960.517, 962.3976, 964.1482, 
    967.5267, 971.8688, 979.5736, 986.37, 992.6512, 992.1884, 992.3513, 
    993.7643, 990.2716, 994.3398, 995.0259, 993.2343, 1003.716, 1000.7, 
    1003.786, 1001.82, 954.3201, 956.6383, 955.3845, 957.7448, 956.0811, 
    963.5187, 965.735, 976.0355, 971.7831, 978.5663, 972.468, 973.5436, 
    978.7901, 972.7956, 985.9935, 977.0107, 993.8193, 984.717, 994.395, 
    992.6239, 995.5592, 998.2023, 1001.546, 1007.772, 1006.324, 1011.573, 
    960.1123, 963.1534, 962.8846, 966.0395, 968.339, 973.3571, 981.5072, 
    978.4274, 984.0947, 985.24, 976.6351, 981.9022, 965.1832, 967.8492, 
    966.2599, 960.3519, 979.1362, 969.4886, 987.4434, 982.1121, 997.8247, 
    989.9525, 1005.528, 1012.331, 1018.812, 1026.49, 964.8176, 962.7454, 
    966.4084, 971.4264, 976.1241, 982.4358, 983.0856, 984.2781, 987.379, 
    990.0006, 984.6562, 990.6598, 968.4703, 979.9818, 961.9636, 967.3904, 
    971.1291, 969.4853, 978.0765, 980.1221, 988.5173, 984.1605, 1010.644, 
    998.7629, 1032.29, 1022.79, 962.0225, 964.8105, 974.3096, 969.7685, 
    982.8596, 986.1326, 988.808, 992.2487, 992.6211, 994.6717, 991.3157, 
    994.5385, 982.4493, 987.8174, 973.2145, 976.732, 975.1108, 973.3385, 
    978.8276, 984.74, 984.8663, 986.7768, 992.1995, 982.9133, 1012.199, 
    993.9232, 967.7681, 973.0344, 973.79, 971.741, 985.8036, 980.6649, 
    994.6215, 990.8128, 997.0675, 993.9503, 993.4932, 989.5195, 987.0609, 
    980.8995, 975.9388, 972.0376, 972.9421, 977.2364, 985.1036, 992.6552, 
    990.9918, 996.5895, 981.8994, 988.0099, 985.6401, 991.8417, 978.346, 
    989.8188, 975.4534, 976.6972, 980.5634, 988.4275, 990.1821, 992.0635, 
    990.9017, 985.3047, 984.3931, 980.4689, 979.3909, 976.4261, 973.9844, 
    976.215, 978.5679, 985.3068, 991.4548, 998.2401, 999.9137, 1007.982, 
    1001.406, 1012.302, 1003.026, 1019.188, 990.4902, 1002.754, 980.7397, 
    983.0674, 987.3049, 997.1524, 991.8124, 998.0625, 984.3574, 977.3856, 
    975.5958, 972.2741, 975.6719, 975.3947, 978.665, 977.6119, 985.532, 
    981.2628, 993.4819, 998.0126, 1011.02, 1019.156, 1027.567, 1031.239, 
    1032.351, 1032.816,
  1829.886, 1849.348, 1845.52, 1861.544, 1852.608, 1863.169, 1833.786, 
    1850.133, 1839.651, 1831.614, 1893.766, 1862.268, 1928.089, 1906.809, 
    1960.685, 1924.735, 1968.115, 1959.626, 1985.501, 1977.986, 2012.206, 
    1988.998, 2030.642, 2006.59, 2010.298, 1988.246, 1868.489, 1889.765, 
    1867.249, 1870.237, 1868.894, 1852.792, 1844.821, 1828.42, 1831.368, 
    1843.427, 1871.585, 1861.894, 1886.584, 1886.016, 1914.574, 1901.55, 
    1950.842, 1936.753, 1978.298, 1967.606, 1977.792, 1974.687, 1977.833, 
    1962.22, 1968.865, 1955.288, 1903.971, 1918.857, 1875.385, 1850.523, 
    1834.495, 1823.349, 1824.913, 1827.906, 1843.498, 1858.491, 1870.144, 
    1878.052, 1885.935, 1910.37, 1923.66, 1953.728, 1948.255, 1957.552, 
    1966.552, 1981.941, 1979.383, 1986.251, 1957.303, 1976.403, 1945.158, 
    1953.561, 1888.101, 1864.495, 1854.71, 1846.254, 1826.119, 1839.96, 
    1834.47, 1847.603, 1856.084, 1851.876, 1878.27, 1867.887, 1924.456, 
    1899.514, 1965.496, 1949.375, 1969.418, 1959.115, 1976.866, 1960.869, 
    1988.824, 1995.068, 1990.795, 2007.356, 1959.994, 1977.793, 1851.759, 
    1852.443, 1855.64, 1841.699, 1840.855, 1828.339, 1839.463, 1844.257, 
    1856.578, 1863.974, 1871.08, 1886.969, 1905.163, 1931.442, 1950.408, 
    1963.389, 1955.399, 1962.448, 1954.573, 1950.913, 1992.722, 1968.928, 
    2004.949, 2002.904, 1986.415, 2003.134, 1852.924, 1848.992, 1835.518, 
    1846.04, 1826.99, 1837.588, 1843.758, 1868.104, 1873.57, 1878.68, 
    1888.885, 1902.211, 1926.232, 1947.384, 1967.079, 1965.616, 1966.131, 
    1970.605, 1959.577, 1972.433, 1974.615, 1968.925, 2002.631, 1992.829, 
    2002.861, 1996.46, 1850.268, 1856.909, 1853.312, 1860.092, 1855.309, 
    1876.84, 1883.43, 1915.141, 1901.946, 1923.064, 1904.062, 1907.391, 
    1923.767, 1905.075, 1946.214, 1918.187, 1970.779, 1942.257, 1972.608, 
    1966.992, 1976.314, 1984.775, 1995.569, 2015.952, 2011.177, 2028.578, 
    1866.931, 1875.774, 1874.989, 1884.356, 1891.367, 1906.813, 1932.338, 
    1922.628, 1940.333, 1943.877, 1917.013, 1933.58, 1881.755, 1889.87, 
    1885.026, 1867.625, 1924.855, 1894.888, 1950.725, 1934.225, 1983.562, 
    1958.575, 2008.563, 2031.113, 2053.029, 2079.234, 1880.647, 1874.583, 
    1885.478, 1900.846, 1915.417, 1935.22, 1937.22, 1940.9, 1950.524, 
    1958.726, 1942.069, 1960.797, 1891.769, 1927.519, 1872.306, 1888.469, 
    1899.93, 1894.878, 1921.526, 1927.961, 1954.078, 1940.536, 2025.48, 
    1986.578, 2099.502, 2066.699, 1872.477, 1880.625, 1909.768, 1895.747, 
    1936.524, 1946.646, 1954.988, 1965.806, 1966.984, 1973.488, 1962.862, 
    1973.064, 1935.261, 1951.892, 1906.371, 1917.316, 1912.259, 1906.755, 
    1923.885, 1942.328, 1942.719, 1948.649, 1965.651, 1936.689, 2030.672, 
    1971.109, 1889.623, 1905.814, 1908.155, 1901.817, 1945.625, 1929.674, 
    1973.328, 1961.279, 1981.135, 1971.195, 1969.745, 1957.216, 1949.533, 
    1930.416, 1914.839, 1902.732, 1905.528, 1918.894, 1943.454, 1967.091, 
    1961.842, 1979.605, 1933.572, 1952.493, 1945.117, 1964.521, 1922.372, 
    1958.155, 1913.326, 1917.207, 1929.354, 1953.797, 1959.296, 1965.221, 
    1961.558, 1944.077, 1941.255, 1929.055, 1925.657, 1916.36, 1908.758, 
    1915.701, 1923.069, 1944.084, 1963.301, 1984.896, 1990.287, 2016.644, 
    1995.115, 2031.019, 2000.38, 2054.315, 1960.264, 1999.495, 1929.911, 
    1937.164, 1950.293, 1981.406, 1964.429, 1984.326, 1941.145, 1919.361, 
    1913.769, 1903.462, 1914.007, 1913.143, 1923.374, 1920.07, 1944.782, 
    1931.565, 1969.709, 1984.166, 2026.734, 2054.207, 2082.894, 2095.755, 
    2099.718, 2101.382,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.547437, 4.565955, 4.56235, 4.577317, 4.56901, 4.578816, 4.551187, 
    4.566692, 4.556789, 4.549101, 4.606462, 4.577985, 4.636159, 4.617906, 
    4.663849, 4.633317, 4.670022, 4.662964, 4.684221, 4.678125, 4.705389, 
    4.687037, 4.719559, 4.701001, 4.703902, 4.686432, 4.583704, 4.602911, 
    4.582568, 4.585303, 4.584075, 4.569182, 4.561691, 4.546023, 4.548864, 
    4.560372, 4.586533, 4.57764, 4.600072, 4.599565, 4.624626, 4.613315, 
    4.655575, 4.643537, 4.678379, 4.669601, 4.677967, 4.675429, 4.678, 
    4.66513, 4.670641, 4.659326, 4.615432, 4.628304, 4.589988, 4.567058, 
    4.551866, 4.541109, 4.542628, 4.545527, 4.56044, 4.57449, 4.585217, 
    4.592403, 4.599492, 4.620997, 4.632403, 4.658013, 4.653382, 4.661228, 
    4.668728, 4.681341, 4.679263, 4.684826, 4.661019, 4.676833, 4.650746, 
    4.657872, 4.601428, 4.580037, 4.570973, 4.563043, 4.543797, 4.557083, 
    4.551842, 4.564314, 4.572253, 4.568325, 4.5926, 4.583152, 4.63308, 
    4.611529, 4.667853, 4.654333, 4.671097, 4.662537, 4.677211, 4.664003, 
    4.686897, 4.691893, 4.688479, 4.701601, 4.663272, 4.677968, 4.568215, 
    4.568856, 4.571839, 4.558734, 4.557933, 4.545945, 4.55661, 4.561158, 
    4.572712, 4.579558, 4.586072, 4.600416, 4.616473, 4.638988, 4.655208, 
    4.666102, 4.65942, 4.665319, 4.658725, 4.655636, 4.690021, 4.670693, 
    4.699712, 4.698102, 4.684959, 4.698284, 4.569305, 4.565621, 4.552846, 
    4.562841, 4.544641, 4.554823, 4.560686, 4.583352, 4.58834, 4.592971, 
    4.602126, 4.613894, 4.634587, 4.652642, 4.669164, 4.667952, 4.668379, 
    4.672076, 4.662923, 4.673579, 4.67537, 4.67069, 4.697887, 4.690106, 
    4.698069, 4.693001, 4.566818, 4.57302, 4.569668, 4.575973, 4.571531, 
    4.591308, 4.597248, 4.625114, 4.613662, 4.631895, 4.615511, 4.618412, 
    4.632494, 4.616395, 4.651647, 4.62773, 4.672219, 4.648268, 4.673723, 
    4.669093, 4.67676, 4.683635, 4.692292, 4.708296, 4.704587, 4.71799, 
    4.582276, 4.590341, 4.589629, 4.598078, 4.604333, 4.617909, 4.639742, 
    4.631524, 4.646618, 4.649653, 4.626723, 4.640794, 4.595743, 4.603003, 
    4.598678, 4.582913, 4.633419, 4.607452, 4.655477, 4.641352, 4.682655, 
    4.662085, 4.702546, 4.719917, 4.736298, 4.755495, 4.594745, 4.589261, 
    4.599082, 4.612699, 4.625352, 4.642213, 4.64394, 4.647104, 4.655307, 
    4.662211, 4.648107, 4.663943, 4.604691, 4.635677, 4.58719, 4.601756, 
    4.611894, 4.607443, 4.630585, 4.636051, 4.658309, 4.646792, 4.715627, 
    4.68509, 4.770141, 4.746274, 4.587346, 4.594726, 4.620475, 4.608211, 
    4.64334, 4.652015, 4.659074, 4.66811, 4.669086, 4.674446, 4.665664, 
    4.674098, 4.642249, 4.656464, 4.617525, 4.626983, 4.62263, 4.617859, 
    4.632594, 4.648329, 4.648663, 4.653717, 4.667983, 4.643482, 4.719583, 
    4.672492, 4.602782, 4.61704, 4.619076, 4.613548, 4.651145, 4.637498, 
    4.674314, 4.664345, 4.680687, 4.672562, 4.671367, 4.660946, 4.654467, 
    4.638124, 4.624855, 4.614349, 4.61679, 4.628335, 4.649292, 4.669175, 
    4.664815, 4.679443, 4.640786, 4.656971, 4.650712, 4.667044, 4.631306, 
    4.661735, 4.62355, 4.626889, 4.637228, 4.658072, 4.662688, 4.667625, 
    4.664578, 4.649825, 4.647409, 4.636976, 4.634099, 4.626162, 4.619599, 
    4.625596, 4.631899, 4.64983, 4.666029, 4.683733, 4.688072, 4.708832, 
    4.691931, 4.719847, 4.696112, 4.737245, 4.663498, 4.69541, 4.637698, 
    4.643892, 4.655111, 4.680908, 4.666967, 4.683272, 4.647315, 4.628735, 
    4.623933, 4.614988, 4.624138, 4.623393, 4.632159, 4.629341, 4.650426, 
    4.639091, 4.671338, 4.683143, 4.716585, 4.737165, 4.75817, 4.767464, 
    4.770294, 4.771478,
  5.63329, 5.656574, 5.652041, 5.670864, 5.660416, 5.67275, 5.638004, 
    5.657501, 5.645048, 5.635382, 5.707526, 5.671704, 5.744902, 5.721928, 
    5.779763, 5.741323, 5.787535, 5.778648, 5.805419, 5.79774, 5.832085, 
    5.808966, 5.849941, 5.826556, 5.830211, 5.808205, 5.678897, 5.703058, 
    5.677469, 5.680909, 5.679364, 5.660632, 5.651212, 5.631512, 5.635084, 
    5.649554, 5.682456, 5.671269, 5.699488, 5.698849, 5.730386, 5.716151, 
    5.769344, 5.754189, 5.798061, 5.787005, 5.797542, 5.794345, 5.797584, 
    5.781375, 5.788316, 5.774067, 5.718815, 5.735014, 5.686802, 5.657961, 
    5.638858, 5.625334, 5.627244, 5.630888, 5.649639, 5.667308, 5.680801, 
    5.689841, 5.698758, 5.725818, 5.740173, 5.772414, 5.766583, 5.776462, 
    5.785906, 5.801791, 5.799174, 5.806181, 5.776199, 5.796113, 5.763265, 
    5.772236, 5.701193, 5.674285, 5.662885, 5.652913, 5.628714, 5.645417, 
    5.638828, 5.654511, 5.664495, 5.659555, 5.690088, 5.678204, 5.741024, 
    5.713903, 5.784804, 5.76778, 5.788889, 5.778111, 5.796589, 5.779956, 
    5.80879, 5.815083, 5.810782, 5.827312, 5.779036, 5.797543, 5.659417, 
    5.660223, 5.663975, 5.647494, 5.646486, 5.631414, 5.644823, 5.650541, 
    5.665073, 5.673683, 5.681876, 5.699921, 5.720125, 5.748462, 5.768882, 
    5.7826, 5.774185, 5.781614, 5.77331, 5.769421, 5.812725, 5.788381, 
    5.824933, 5.822906, 5.806348, 5.823134, 5.660788, 5.656154, 5.64009, 
    5.652658, 5.629775, 5.642577, 5.649948, 5.678453, 5.684729, 5.690555, 
    5.702072, 5.716879, 5.742922, 5.765651, 5.786456, 5.784929, 5.785467, 
    5.790122, 5.778597, 5.792016, 5.794271, 5.788377, 5.822634, 5.812832, 
    5.822862, 5.816479, 5.65766, 5.66546, 5.661244, 5.669173, 5.663587, 
    5.688462, 5.695935, 5.730999, 5.716588, 5.739534, 5.718915, 5.722565, 
    5.740288, 5.720027, 5.764398, 5.734292, 5.790303, 5.760145, 5.792197, 
    5.786366, 5.796021, 5.804681, 5.815586, 5.835748, 5.831075, 5.847963, 
    5.677101, 5.687246, 5.68635, 5.696979, 5.704849, 5.721932, 5.749412, 
    5.739067, 5.758068, 5.761888, 5.733024, 5.750735, 5.694041, 5.703175, 
    5.697734, 5.677902, 5.741452, 5.708774, 5.76922, 5.751438, 5.803446, 
    5.777541, 5.828503, 5.850392, 5.871037, 5.895238, 5.692786, 5.685887, 
    5.698243, 5.715375, 5.731299, 5.752522, 5.754696, 5.75868, 5.769006, 
    5.7777, 5.759942, 5.779881, 5.705298, 5.744294, 5.683282, 5.701606, 
    5.714363, 5.708763, 5.737885, 5.744765, 5.772786, 5.758287, 5.844985, 
    5.806513, 5.913707, 5.883612, 5.683478, 5.692762, 5.725161, 5.709728, 
    5.75394, 5.764862, 5.773749, 5.785128, 5.786356, 5.793107, 5.782048, 
    5.792669, 5.752567, 5.770463, 5.721449, 5.733352, 5.727873, 5.721869, 
    5.740414, 5.760221, 5.760642, 5.767005, 5.784967, 5.754119, 5.84997, 
    5.790646, 5.702898, 5.720838, 5.723401, 5.716444, 5.763766, 5.746587, 
    5.792942, 5.780386, 5.800967, 5.790734, 5.78923, 5.776107, 5.767949, 
    5.747375, 5.730673, 5.717453, 5.720524, 5.735054, 5.761434, 5.786469, 
    5.780979, 5.799401, 5.750726, 5.771102, 5.763221, 5.783785, 5.738792, 
    5.777099, 5.729032, 5.733234, 5.746246, 5.772488, 5.778301, 5.784517, 
    5.78068, 5.762104, 5.759064, 5.745929, 5.742308, 5.732318, 5.724059, 
    5.731606, 5.73954, 5.762111, 5.782508, 5.804804, 5.810269, 5.836423, 
    5.81513, 5.850302, 5.820396, 5.872231, 5.77932, 5.819512, 5.746838, 
    5.754635, 5.76876, 5.801246, 5.783689, 5.804224, 5.758944, 5.735557, 
    5.729513, 5.718256, 5.729771, 5.728834, 5.739866, 5.736319, 5.762861, 
    5.748593, 5.789193, 5.80406, 5.846193, 5.87213, 5.898612, 5.91033, 
    5.9139, 5.915393,
  8.097958, 8.132158, 8.1255, 8.153154, 8.137803, 8.155926, 8.10488, 8.13352, 
    8.115227, 8.101029, 8.207046, 8.154389, 8.262018, 8.228224, 8.313323, 
    8.256754, 8.324766, 8.311683, 8.351101, 8.339793, 8.390382, 8.356324, 
    8.416696, 8.382236, 8.387621, 8.355203, 8.164961, 8.200477, 8.162861, 
    8.167916, 8.165647, 8.138121, 8.124281, 8.095345, 8.100592, 8.121845, 
    8.170191, 8.153751, 8.195228, 8.194289, 8.240664, 8.219728, 8.297988, 
    8.275683, 8.340264, 8.323986, 8.3395, 8.334793, 8.339561, 8.315697, 
    8.325915, 8.304939, 8.223646, 8.247472, 8.176579, 8.134196, 8.106135, 
    8.086273, 8.089079, 8.09443, 8.12197, 8.147929, 8.167759, 8.181046, 
    8.194154, 8.233946, 8.255061, 8.302505, 8.293924, 8.308463, 8.322368, 
    8.345758, 8.341904, 8.352222, 8.308077, 8.337397, 8.28904, 8.302244, 
    8.197734, 8.158183, 8.14143, 8.12678, 8.091237, 8.115769, 8.106091, 
    8.129128, 8.143796, 8.136539, 8.181409, 8.163941, 8.256314, 8.216423, 
    8.320745, 8.295685, 8.32676, 8.31089, 8.338098, 8.313608, 8.356065, 
    8.365335, 8.358999, 8.38335, 8.312253, 8.339501, 8.136335, 8.137519, 
    8.143032, 8.118819, 8.11734, 8.095202, 8.114897, 8.123296, 8.144646, 
    8.157297, 8.169338, 8.195864, 8.225573, 8.267257, 8.297307, 8.3175, 
    8.305113, 8.316049, 8.303824, 8.2981, 8.361861, 8.326012, 8.379845, 
    8.376858, 8.352468, 8.377194, 8.13835, 8.131541, 8.107945, 8.126407, 
    8.092794, 8.111596, 8.122425, 8.164309, 8.173532, 8.182095, 8.199026, 
    8.220798, 8.259107, 8.292552, 8.323176, 8.32093, 8.32172, 8.328575, 
    8.311606, 8.331363, 8.334683, 8.326005, 8.376458, 8.36202, 8.376794, 
    8.367391, 8.133754, 8.145214, 8.13902, 8.150671, 8.142462, 8.179018, 
    8.190004, 8.241567, 8.22037, 8.254122, 8.223793, 8.229161, 8.25523, 
    8.225429, 8.290708, 8.24641, 8.328841, 8.284448, 8.33163, 8.323044, 
    8.337262, 8.350014, 8.366076, 8.39578, 8.388893, 8.413781, 8.162321, 
    8.177232, 8.175916, 8.191539, 8.20311, 8.22823, 8.268655, 8.253434, 
    8.281391, 8.287013, 8.244545, 8.270601, 8.187221, 8.200648, 8.19265, 
    8.163498, 8.256943, 8.20888, 8.297805, 8.271636, 8.348194, 8.310053, 
    8.385105, 8.41736, 8.447794, 8.483485, 8.185375, 8.175234, 8.193398, 
    8.218587, 8.242007, 8.273231, 8.276429, 8.282291, 8.29749, 8.310287, 
    8.284148, 8.313497, 8.20377, 8.261124, 8.171405, 8.198341, 8.217099, 
    8.208863, 8.251695, 8.261817, 8.303052, 8.281714, 8.409392, 8.352713, 
    8.510731, 8.466338, 8.171694, 8.18534, 8.232979, 8.210284, 8.275317, 
    8.291389, 8.304471, 8.321222, 8.32303, 8.33297, 8.316688, 8.332325, 
    8.273297, 8.299633, 8.22752, 8.245027, 8.236968, 8.228138, 8.255415, 
    8.28456, 8.28518, 8.294544, 8.320984, 8.275581, 8.416738, 8.329345, 
    8.200241, 8.226622, 8.23039, 8.22016, 8.289777, 8.264498, 8.332726, 
    8.314241, 8.344544, 8.329475, 8.327261, 8.307942, 8.295934, 8.265656, 
    8.241086, 8.221642, 8.22616, 8.24753, 8.286345, 8.323195, 8.315113, 
    8.342238, 8.270588, 8.300574, 8.288976, 8.319245, 8.253031, 8.309402, 
    8.238672, 8.244854, 8.263997, 8.302614, 8.311171, 8.320323, 8.314674, 
    8.287332, 8.282857, 8.26353, 8.258203, 8.243507, 8.231359, 8.242458, 
    8.254129, 8.287341, 8.317365, 8.350196, 8.358244, 8.396774, 8.365404, 
    8.417227, 8.37316, 8.449554, 8.312672, 8.371859, 8.264868, 8.27634, 
    8.297128, 8.344954, 8.319102, 8.34934, 8.282681, 8.24827, 8.239381, 
    8.222824, 8.239759, 8.23838, 8.25461, 8.249393, 8.288445, 8.267449, 
    8.327207, 8.3491, 8.411171, 8.449406, 8.488461, 8.50575, 8.511017, 8.51322,
  12.66457, 12.72004, 12.70924, 12.7541, 12.72919, 12.7586, 12.6758, 
    12.72225, 12.69257, 12.66955, 12.84161, 12.75611, 12.93096, 12.87602, 
    13.01443, 12.9224, 13.03306, 13.01176, 13.07595, 13.05753, 13.13997, 
    13.08446, 13.18289, 13.12669, 13.13547, 13.08264, 12.77326, 12.83093, 
    12.76986, 12.77806, 12.77438, 12.72971, 12.70726, 12.66034, 12.66884, 
    12.70331, 12.78175, 12.75507, 12.82241, 12.82088, 12.89624, 12.86221, 
    12.98947, 12.95318, 13.0583, 13.03179, 13.05706, 13.04939, 13.05716, 
    13.0183, 13.03493, 13.00079, 12.86858, 12.9073, 12.79213, 12.72334, 
    12.67783, 12.64563, 12.65018, 12.65886, 12.70351, 12.74562, 12.77781, 
    12.79938, 12.82067, 12.88531, 12.91964, 12.99682, 12.98286, 13.00652, 
    13.02916, 13.06725, 13.06097, 13.07778, 13.00589, 13.05363, 12.97491, 
    12.9964, 12.82648, 12.76226, 12.73508, 12.71131, 12.65368, 12.69345, 
    12.67776, 12.71512, 12.73892, 12.72714, 12.79997, 12.77161, 12.92168, 
    12.85684, 13.02652, 12.98572, 13.03631, 13.01047, 13.05477, 13.0149, 
    13.08404, 13.09914, 13.08882, 13.12851, 13.01269, 13.05706, 12.72681, 
    12.72873, 12.73768, 12.6984, 12.696, 12.66011, 12.69204, 12.70566, 
    12.7403, 12.76083, 12.78037, 12.82344, 12.87171, 12.93948, 12.98837, 
    13.02123, 13.00107, 13.01887, 12.99897, 12.98965, 13.09348, 13.03509, 
    13.12279, 13.11793, 13.07818, 13.11847, 12.73008, 12.71904, 12.68077, 
    12.71071, 12.6562, 12.68669, 12.70425, 12.77221, 12.78718, 12.80108, 
    12.82858, 12.86395, 12.92622, 12.98063, 13.03047, 13.02682, 13.0281, 
    13.03926, 13.01164, 13.0438, 13.04921, 13.03508, 13.11727, 13.09374, 
    13.11782, 13.1025, 12.72262, 12.74122, 12.73117, 12.75007, 12.73675, 
    12.79609, 12.81393, 12.8977, 12.86325, 12.91812, 12.86882, 12.87754, 
    12.91992, 12.87147, 12.97762, 12.90558, 13.0397, 12.96744, 13.04424, 
    13.03026, 13.05341, 13.07418, 13.10035, 13.14877, 13.13754, 13.17813, 
    12.76898, 12.79319, 12.79105, 12.81642, 12.83521, 12.87603, 12.94175, 
    12.917, 12.96247, 12.97161, 12.90255, 12.94492, 12.80941, 12.83121, 
    12.81822, 12.77089, 12.9227, 12.84459, 12.98917, 12.9466, 13.07122, 
    13.00911, 13.13137, 13.18397, 13.23363, 13.29191, 12.80641, 12.78994, 
    12.81944, 12.86036, 12.89842, 12.94919, 12.9544, 12.96393, 12.98866, 
    13.00949, 12.96695, 13.01472, 12.83628, 12.9295, 12.78373, 12.82747, 
    12.85794, 12.84456, 12.91417, 12.93063, 12.99771, 12.96299, 13.17097, 
    13.07858, 13.33643, 13.26391, 12.78419, 12.80635, 12.88375, 12.84687, 
    12.95259, 12.97873, 13.00002, 13.02729, 13.03024, 13.04642, 13.01991, 
    13.04537, 12.9493, 12.99215, 12.87487, 12.90333, 12.89023, 12.87588, 
    12.92022, 12.96762, 12.96863, 12.98387, 13.0269, 12.95302, 13.18295, 
    13.04052, 12.83055, 12.87341, 12.87954, 12.86291, 12.97611, 12.93499, 
    13.04603, 13.01593, 13.06527, 13.04073, 13.03712, 13.00567, 12.98613, 
    12.93687, 12.89692, 12.86532, 12.87266, 12.9074, 12.97053, 13.03051, 
    13.01735, 13.06152, 12.94489, 12.99368, 12.97481, 13.02407, 12.91634, 
    13.00805, 12.893, 12.90305, 12.93417, 12.997, 13.01093, 13.02583, 
    13.01663, 12.97213, 12.96485, 12.93342, 12.92475, 12.90086, 12.88111, 
    12.89915, 12.91813, 12.97215, 13.02101, 13.07448, 13.08759, 13.15039, 
    13.09926, 13.18375, 13.1119, 13.2365, 13.01337, 13.10978, 12.93559, 
    12.95425, 12.98807, 13.06594, 13.02384, 13.07308, 12.96457, 12.9086, 
    12.89415, 12.86724, 12.89477, 12.89252, 12.91891, 12.91043, 12.97394, 
    12.93979, 13.03704, 13.07269, 13.17387, 13.23626, 13.30004, 13.32829, 
    13.3369, 13.3405,
  20.59555, 20.6916, 20.67289, 20.75065, 20.70747, 20.75845, 20.61498, 
    20.69543, 20.64403, 20.60417, 20.90253, 20.75413, 21.05791, 20.96234, 
    21.20336, 21.04301, 21.23585, 21.1987, 21.31072, 21.27856, 21.4226, 
    21.32558, 21.49769, 21.39938, 21.41473, 21.32239, 20.78389, 20.88399, 
    20.77798, 20.79221, 20.78582, 20.70836, 20.66946, 20.58822, 20.60294, 
    20.66262, 20.79862, 20.75233, 20.86919, 20.86654, 20.9975, 20.93834, 
    21.15984, 21.09661, 21.2799, 21.23364, 21.27773, 21.26435, 21.2779, 
    21.2101, 21.23912, 21.17956, 20.9494, 21.01675, 20.81661, 20.69733, 
    20.6185, 20.56278, 20.57064, 20.58566, 20.66297, 20.73595, 20.79177, 
    20.8292, 20.86616, 20.9785, 21.03822, 21.17266, 21.14831, 21.18956, 
    21.22904, 21.29552, 21.28456, 21.31391, 21.18847, 21.27175, 21.13446, 
    21.17191, 20.87625, 20.7648, 20.71767, 20.67648, 20.5767, 20.64555, 
    20.61838, 20.68308, 20.72432, 20.70391, 20.83022, 20.78102, 21.04177, 
    20.929, 21.22443, 21.15331, 21.24152, 21.19645, 21.27374, 21.20417, 
    21.32484, 21.35123, 21.3332, 21.40255, 21.20032, 21.27773, 20.70334, 
    20.70667, 20.72218, 20.65412, 20.64996, 20.58782, 20.6431, 20.66669, 
    20.72671, 20.76231, 20.79622, 20.87098, 20.95484, 21.07274, 21.15791, 
    21.21522, 21.18005, 21.21109, 21.1764, 21.16016, 21.34134, 21.23939, 
    21.39256, 21.38405, 21.31461, 21.38501, 20.70901, 20.68987, 20.62358, 
    20.67544, 20.58107, 20.63383, 20.66425, 20.78205, 20.80803, 20.83216, 
    20.8799, 20.94136, 21.04967, 21.14442, 21.23134, 21.22495, 21.2272, 
    21.24667, 21.19848, 21.2546, 21.26403, 21.23937, 21.38291, 21.34179, 
    21.38387, 21.35708, 20.69608, 20.72831, 20.71089, 20.74366, 20.72057, 
    20.82349, 20.85446, 21.00005, 20.94015, 21.03556, 20.94982, 20.96498, 
    21.0387, 20.95444, 21.13919, 21.01375, 21.24743, 21.12144, 21.25536, 
    21.23096, 21.27136, 21.30763, 21.35334, 21.43799, 21.41836, 21.48936, 
    20.77645, 20.81845, 20.81474, 20.85878, 20.89142, 20.96235, 21.0767, 
    21.03362, 21.11278, 21.12872, 21.00847, 21.08222, 20.84661, 20.88448, 
    20.86192, 20.77977, 21.04355, 20.90771, 21.15932, 21.08515, 21.30245, 
    21.19407, 21.40756, 21.49958, 21.58658, 21.68879, 20.84141, 20.81282, 
    20.86403, 20.93511, 21.0013, 21.08966, 21.09872, 21.11534, 21.15843, 
    21.19474, 21.1206, 21.20385, 20.89328, 21.05538, 20.80204, 20.87797, 
    20.93091, 20.90766, 21.0287, 21.05734, 21.17421, 21.1137, 21.47684, 
    21.3153, 21.76696, 21.63965, 20.80285, 20.8413, 20.97577, 20.91167, 
    21.09557, 21.14113, 21.17823, 21.22579, 21.23092, 21.25916, 21.21291, 
    21.25733, 21.08985, 21.16451, 20.96035, 21.00983, 20.98705, 20.96209, 
    21.03922, 21.12177, 21.12352, 21.15007, 21.22511, 21.09632, 21.4978, 
    21.24886, 20.88333, 20.95781, 20.96846, 20.93955, 21.13655, 21.06493, 
    21.25847, 21.20597, 21.29207, 21.24924, 21.24294, 21.18808, 21.15401, 
    21.06821, 20.99869, 20.94374, 20.9565, 21.01692, 21.12682, 21.23139, 
    21.20844, 21.28551, 21.08218, 21.16718, 21.13428, 21.22017, 21.03248, 
    21.19222, 20.99187, 21.00935, 21.06351, 21.17296, 21.19725, 21.22323, 
    21.20719, 21.12962, 21.11694, 21.06219, 21.04711, 21.00554, 20.9712, 
    21.00257, 21.03559, 21.12965, 21.21483, 21.30815, 21.33105, 21.44083, 
    21.35143, 21.4992, 21.37352, 21.59161, 21.20151, 21.36981, 21.06598, 
    21.09847, 21.1574, 21.29324, 21.21977, 21.30571, 21.11644, 21.01901, 
    20.99387, 20.94708, 20.99494, 20.99104, 21.03695, 21.02218, 21.13278, 
    21.07329, 21.24279, 21.30503, 21.48191, 21.59119, 21.70305, 21.75266, 
    21.76778, 21.77411,
  34.63898, 34.81974, 34.78448, 34.93107, 34.84964, 34.94579, 34.67551, 
    34.82695, 34.73016, 34.65519, 35.21814, 34.93763, 35.51294, 35.33147, 
    35.78992, 35.48462, 35.85194, 35.78104, 35.99503, 35.93353, 36.20937, 
    36.02347, 36.35357, 36.16483, 36.19426, 36.01736, 34.9938, 35.18304, 
    34.98264, 35.00952, 34.99745, 34.85132, 34.77803, 34.62521, 34.65288, 
    34.76515, 35.02161, 34.93423, 35.15502, 35.15001, 35.39818, 35.28597, 
    35.70694, 35.58654, 35.93609, 35.84771, 35.93194, 35.90636, 35.93227, 
    35.80278, 35.85817, 35.74453, 35.30695, 35.43474, 35.05562, 34.83053, 
    34.68213, 34.5774, 34.59218, 34.62038, 34.76581, 34.90334, 35.00868, 
    35.07941, 35.1493, 35.36214, 35.47552, 35.73137, 35.68498, 35.7636, 
    35.83894, 35.96596, 35.945, 36.00114, 35.76151, 35.92051, 35.6586, 
    35.72995, 35.1684, 34.95778, 34.86886, 34.79126, 34.60355, 34.73302, 
    34.6819, 34.80369, 34.88141, 34.84294, 35.08134, 34.98838, 35.48226, 
    35.26828, 35.83014, 35.69449, 35.86276, 35.77674, 35.92432, 35.79146, 
    36.02205, 36.07257, 36.03804, 36.17092, 35.78412, 35.93194, 34.84186, 
    34.84813, 34.87736, 34.74915, 34.74133, 34.62445, 34.72841, 34.77283, 
    34.88592, 34.95307, 35.01708, 35.15842, 35.31726, 35.54114, 35.70326, 
    35.81255, 35.74547, 35.80468, 35.7385, 35.70755, 36.05363, 35.8587, 
    36.15176, 36.13545, 36.00248, 36.13729, 34.85254, 34.81647, 34.69169, 
    34.78928, 34.61176, 34.71098, 34.76822, 34.99033, 35.03939, 35.085, 
    35.1753, 35.2917, 35.49728, 35.67757, 35.84332, 35.83113, 35.83543, 
    35.8726, 35.78062, 35.88774, 35.90577, 35.85867, 36.13327, 36.05449, 
    36.1351, 36.08378, 34.82819, 34.88893, 34.85609, 34.91788, 34.87434, 
    35.0686, 35.12716, 35.40303, 35.28941, 35.47047, 35.30774, 35.33649, 
    35.47643, 35.3165, 35.6676, 35.42903, 35.87405, 35.6338, 35.88919, 
    35.8426, 35.91978, 35.98911, 36.07661, 36.23891, 36.20123, 36.33757, 
    34.97977, 35.05909, 35.05208, 35.13534, 35.19711, 35.33151, 35.54867, 
    35.46677, 35.61732, 35.64766, 35.41902, 35.55915, 35.11231, 35.18396, 
    35.14127, 34.98602, 35.48564, 35.22794, 35.70595, 35.56473, 35.97921, 
    35.77221, 36.18051, 36.35721, 36.52464, 36.72184, 35.10248, 35.04845, 
    35.14526, 35.27986, 35.4054, 35.57332, 35.59056, 35.62218, 35.70425, 
    35.77348, 35.63219, 35.79086, 35.20063, 35.50813, 35.02807, 35.17164, 
    35.2719, 35.22786, 35.45743, 35.51186, 35.73433, 35.61906, 36.31349, 
    36.0038, 36.87302, 36.62698, 35.02961, 35.10229, 35.35696, 35.23545, 
    35.58456, 35.67129, 35.742, 35.83272, 35.84253, 35.89646, 35.80815, 
    35.89296, 35.57368, 35.71584, 35.3277, 35.4216, 35.37835, 35.33101, 
    35.47742, 35.63441, 35.63776, 35.68833, 35.83143, 35.58599, 36.35379, 
    35.87679, 35.18179, 35.32288, 35.34308, 35.28828, 35.66258, 35.52629, 
    35.89514, 35.79489, 35.95936, 35.87749, 35.86547, 35.76078, 35.69584, 
    35.53252, 35.40045, 35.29622, 35.32042, 35.43505, 35.64405, 35.84343, 
    35.79961, 35.94682, 35.55908, 35.72092, 35.65825, 35.82201, 35.4646, 
    35.76868, 35.3875, 35.42068, 35.52359, 35.73195, 35.77826, 35.82785, 
    35.79724, 35.64937, 35.62523, 35.52108, 35.49241, 35.41345, 35.34827, 
    35.40782, 35.47051, 35.64943, 35.81181, 35.9901, 36.03392, 36.24435, 
    36.07294, 36.35648, 36.11526, 36.53433, 35.78639, 36.10815, 35.52828, 
    35.59008, 35.70229, 35.96159, 35.82123, 35.98545, 35.62428, 35.43902, 
    35.3913, 35.30255, 35.39333, 35.38593, 35.4731, 35.44505, 35.65539, 
    35.54218, 35.86518, 35.98414, 36.32325, 36.53352, 36.7494, 36.84534, 
    36.87461, 36.88686,
  60.67812, 61.07083, 60.99409, 61.31372, 61.13599, 61.34589, 60.75732, 
    61.08654, 60.87596, 60.71325, 61.9436, 61.32805, 62.59598, 62.19373, 
    63.21417, 62.53307, 63.35332, 63.19427, 63.67535, 63.53676, 64.1604, 
    63.73952, 64.48857, 64.05934, 64.12612, 63.72573, 61.45091, 61.86631, 
    61.42648, 61.48533, 61.4589, 61.13967, 60.98005, 60.64828, 60.70824, 
    60.95203, 61.51183, 61.32064, 61.80466, 61.79365, 62.34135, 62.09321, 
    63.02843, 62.75974, 63.54253, 63.34382, 63.53318, 63.47564, 63.53393, 
    63.243, 63.36732, 63.11252, 62.13955, 62.42237, 61.58636, 61.09434, 
    60.77169, 60.54478, 60.57676, 60.63782, 60.95346, 61.25315, 61.48349, 
    61.63854, 61.79207, 62.26156, 62.51286, 63.08306, 62.97935, 63.15522, 
    63.32412, 63.60981, 63.5626, 63.68912, 63.15054, 63.50746, 62.92043, 
    63.0799, 61.83408, 61.3721, 61.17791, 61.00883, 60.60137, 60.88219, 
    60.77119, 61.03589, 61.20528, 61.12138, 61.6428, 61.43905, 62.52781, 
    62.05416, 63.30437, 63.0006, 63.37762, 63.18466, 63.51603, 63.21764, 
    63.73633, 63.85044, 63.77242, 64.07315, 63.20119, 63.5332, 61.11904, 
    61.13271, 61.19645, 60.91724, 60.90023, 60.64664, 60.87217, 60.96872, 
    61.21512, 61.36182, 61.5019, 61.81213, 62.16233, 62.65869, 63.02021, 
    63.26492, 63.11462, 63.24727, 63.09903, 63.02979, 63.80764, 63.36849, 
    64.02972, 63.99276, 63.69214, 63.99692, 61.14231, 61.06372, 60.79243, 
    61.00454, 60.61915, 60.8343, 60.95869, 61.44333, 61.55079, 61.65081, 
    61.84928, 62.10587, 62.56117, 62.96279, 63.33397, 63.30662, 63.31625, 
    63.39974, 63.19335, 63.43375, 63.4743, 63.36842, 63.98781, 63.80959, 
    63.99197, 63.8758, 61.08924, 61.22169, 61.15005, 61.28492, 61.18986, 
    61.61485, 61.7434, 62.35209, 62.1008, 62.50164, 62.14127, 62.20483, 
    62.51487, 62.16063, 62.94054, 62.40972, 63.40299, 62.86511, 63.43701, 
    63.33235, 63.50581, 63.66199, 63.85958, 64.22751, 64.14191, 64.4521, 
    61.4202, 61.59398, 61.57861, 61.76139, 61.89728, 62.19381, 62.67543, 
    62.49344, 62.82833, 62.89602, 62.38752, 62.69877, 61.71079, 61.86834, 
    61.77442, 61.43389, 62.53532, 61.96521, 63.02622, 62.71117, 63.63968, 
    63.17449, 64.09491, 64.49689, 64.87986, 65.33361, 61.68919, 61.57066, 
    61.7832, 62.07972, 62.35733, 62.7303, 62.7687, 62.83917, 63.02241, 
    63.17733, 62.86152, 63.21629, 61.90504, 62.58529, 61.52598, 61.84122, 
    62.06215, 61.96502, 62.4727, 62.59358, 63.08968, 62.83222, 64.39722, 
    63.69513, 65.68346, 65.11497, 61.52935, 61.68877, 62.2501, 61.98175, 
    62.75535, 62.94876, 63.10686, 63.31018, 63.33219, 63.45336, 63.25504, 
    63.44549, 62.7311, 63.04832, 62.18539, 62.39325, 62.29745, 62.19272, 
    62.51709, 62.86647, 62.87393, 62.98683, 63.30727, 62.75852, 64.48909, 
    63.40913, 61.86355, 62.17475, 62.2194, 62.09832, 62.92932, 62.62566, 
    63.4504, 63.22533, 63.59494, 63.41073, 63.38372, 63.14891, 63.00362, 
    62.63952, 62.34638, 62.11584, 62.16929, 62.42306, 62.88795, 63.3342, 
    63.23591, 63.5667, 62.69861, 63.0597, 62.91965, 63.28613, 62.48863, 
    63.16659, 62.31769, 62.39119, 62.61966, 63.08437, 63.18806, 63.29924, 
    63.23058, 62.89984, 62.84597, 62.61407, 62.55037, 62.37517, 62.23088, 
    62.3627, 62.50174, 62.89996, 63.26327, 63.66423, 63.76313, 64.23988, 
    63.8513, 64.49522, 63.94703, 64.90211, 63.20626, 63.93095, 62.63008, 
    62.76763, 63.01803, 63.59995, 63.2844, 63.65374, 62.84386, 62.43187, 
    62.3261, 62.12982, 62.33061, 62.31422, 62.50748, 62.44524, 62.91327, 
    62.66099, 63.38306, 63.65079, 64.41946, 64.90024, 65.39728, 65.61928, 
    65.68716, 65.71558,
  116.3177, 117.5456, 117.3041, 118.3151, 117.7513, 118.4176, 116.5637, 
    117.5951, 116.9338, 116.4267, 120.3481, 118.3608, 122.5137, 121.171, 
    124.6257, 122.3021, 125.1096, 124.5568, 126.2417, 125.7524, 127.9808, 
    126.4694, 129.1813, 127.615, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9486, 118.3372, 119.895, 119.8591, 121.6609, 120.8392, 
    123.9848, 123.0673, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7257, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9052, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3957, 122.2342, 124.1727, 123.8163, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4055, 125.6493, 123.6146, 
    124.1618, 119.9907, 118.5013, 117.8839, 117.3504, 116.08, 116.9533, 
    116.6069, 117.4356, 117.9706, 117.7051, 119.3704, 118.7153, 122.2844, 
    120.7108, 124.939, 123.8892, 125.1944, 124.5235, 125.6795, 124.6378, 
    126.4581, 126.8647, 126.5865, 127.6649, 124.5807, 125.7398, 117.6977, 
    117.7409, 117.9426, 117.063, 117.0098, 116.2201, 116.922, 117.2244, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9565, 
    124.8018, 124.2815, 124.7406, 124.2277, 123.9894, 126.712, 125.1625, 
    127.5082, 127.375, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.3369, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.8809, 122.3965, 123.7596, 125.0421, 124.9468, 124.9804, 
    125.2717, 124.5536, 125.3907, 125.5329, 125.1623, 127.3572, 126.7189, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9217, 
    119.2802, 119.696, 121.6967, 120.8642, 122.1966, 120.9977, 121.2077, 
    122.241, 121.0616, 123.6834, 121.8889, 125.2831, 123.4257, 125.4021, 
    125.0365, 125.6435, 126.1945, 126.8974, 128.2247, 127.9137, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1967, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8148, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3096, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4883, 127.7435, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7948, 121.7141, 122.9675, 123.0977, 123.3373, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.0139, 
    120.737, 120.4182, 122.0996, 122.5056, 124.1955, 123.3137, 128.8451, 
    126.3119, 133.7281, 131.5293, 119.0049, 119.519, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2547, 124.9592, 125.0359, 125.4594, 124.7675, 
    125.4319, 122.9702, 124.0532, 121.1434, 121.8339, 121.5149, 121.1676, 
    122.2484, 123.4304, 123.4558, 123.842, 124.9491, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1082, 121.256, 120.856, 123.645, 122.6137, 
    125.4491, 124.6644, 125.9574, 125.3102, 125.2157, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.0429, 
    124.7011, 125.8578, 122.8601, 124.0923, 123.612, 124.8756, 122.153, 
    124.461, 121.5822, 121.8271, 122.5935, 124.1772, 124.5353, 124.9212, 
    124.6826, 123.5443, 123.3605, 122.5746, 122.3602, 121.7736, 121.294, 
    121.7321, 122.1969, 123.5447, 124.7961, 126.2024, 126.5534, 128.2697, 
    126.8678, 129.2058, 127.2107, 130.7228, 124.5983, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9751, 124.8695, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5901, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6128, 133.4764, 
    133.7426, 133.8543,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02010258, -0.01977483, -0.0198381, -0.01957703, -0.01972141, 
    -0.01955111, -0.02003568, -0.01976193, -0.01993623, -0.02007286, 
    -0.01908082, -0.01956547, -0.01859121, -0.01889026, -0.01814875, 
    -0.01863739, -0.01805192, -0.01816269, -0.01783159, -0.01792577, 
    -0.01750933, -0.0177883, -0.01729765, -0.01757554, -0.01753174, 
    -0.01779758, -0.01946692, -0.01914043, -0.01948644, -0.01943947, 
    -0.01946054, -0.0197184, -0.01984971, -0.02012789, -0.02007709, 
    -0.01987294, -0.01941839, -0.01957145, -0.01918825, -0.01919682, 
    -0.01877947, -0.01896642, -0.01827957, -0.01847202, -0.01792183, 
    -0.0180585, -0.01792822, -0.01796762, -0.01792771, -0.01812861, 
    -0.01804224, -0.01822013, -0.01893124, -0.01871918, -0.01935933, 
    -0.01975552, -0.02002358, -0.02021614, -0.0201888, -0.02013678, 
    -0.01987175, -0.01962602, -0.01944094, -0.01931818, -0.01919805, 
    -0.01883919, -0.01865227, -0.01824091, -0.01831445, -0.01819008, 
    -0.01807217, -0.01787601, -0.01790814, -0.01782228, -0.01819337, 
    -0.01794581, -0.01835647, -0.01824315, -0.01916539, -0.01953004, 
    -0.01968716, -0.01982592, -0.0201678, -0.01993103, -0.020024, -0.0198036, 
    -0.01966489, -0.01973336, -0.01931483, -0.0194764, -0.01864126, 
    -0.01899615, -0.01808587, -0.01829933, -0.01803512, -0.01816943, 
    -0.01793995, -0.01814633, -0.01779045, -0.01771395, -0.01776619, 
    -0.01756647, -0.01815785, -0.01792821, -0.01973528, -0.01972409, 
    -0.01967208, -0.01990183, -0.01991599, -0.02012928, -0.01993939, 
    -0.0198591, -0.01965689, -0.0195383, -0.01942629, -0.01918245, 
    -0.01891399, -0.0185454, -0.01828541, -0.01811333, -0.01821865, 
    -0.01812563, -0.01822964, -0.01827862, -0.01774256, -0.01804143, 
    -0.01759505, -0.01761943, -0.01782024, -0.01761668, -0.01971624, 
    -0.01978069, -0.02000615, -0.01982947, -0.02015266, -0.01997104, 
    -0.01986741, -0.01947298, -0.01938748, -0.01930853, -0.01915364, 
    -0.0189568, -0.01861674, -0.01832624, -0.01806534, -0.01808432, 
    -0.01807763, -0.01801984, -0.01816334, -0.0179964, -0.01796854, 
    -0.01804148, -0.0176227, -0.01774126, -0.01761995, -0.01769704, 
    -0.01975972, -0.01965154, -0.01970991, -0.01960029, -0.01967744, 
    -0.01933684, -0.01923597, -0.01877145, -0.01896064, -0.01866054, 
    -0.01892993, -0.01888189, -0.01865078, -0.01891528, -0.0183421, 
    -0.01872857, -0.0180176, -0.01839609, -0.01799416, -0.01806645, 
    -0.01794694, -0.01784062, -0.01770785, -0.01746564, -0.01752141, 
    -0.01732094, -0.01949147, -0.01935332, -0.01936546, -0.01922194, 
    -0.01911652, -0.0188902, -0.01853321, -0.0186666, -0.01842253, 
    -0.01837394, -0.01874507, -0.01851623, -0.01926147, -0.01913888, 
    -0.01921178, -0.01948052, -0.01863573, -0.01906422, -0.01828114, 
    -0.01850722, -0.01785574, -0.01817655, -0.01755219, -0.01729235, 
    -0.01705171, -0.01677497, -0.01927839, -0.01937175, -0.01920495, 
    -0.01897667, -0.01876755, -0.01849334, -0.01846554, -0.01841473, 
    -0.01828384, -0.01817456, -0.01839867, -0.01814728, -0.01911052, 
    -0.01859905, -0.01940715, -0.01915987, -0.01899006, -0.01906437, 
    -0.01868192, -0.01859298, -0.01823623, -0.01841973, -0.01735607, 
    -0.01781822, -0.01656761, -0.0169072, -0.01940448, -0.01927872, 
    -0.01884781, -0.01905153, -0.0184752, -0.01833624, -0.01822412, 
    -0.01808184, -0.01806657, -0.01798292, -0.01812021, -0.01798833, 
    -0.01849276, -0.01826548, -0.01889656, -0.01874081, -0.0188123, 
    -0.01889103, -0.01864916, -0.01839512, -0.01838977, -0.01830912, 
    -0.01808384, -0.01847291, -0.0172973, -0.01801335, -0.01914259, 
    -0.01890459, -0.01887091, -0.01896254, -0.01835012, -0.01856951, 
    -0.01798496, -0.01814096, -0.01788612, -0.01801226, -0.0180309, 
    -0.01819452, -0.01829719, -0.01855938, -0.01877572, -0.01894922, 
    -0.01890873, -0.01871867, -0.01837971, -0.01806517, -0.01813356, 
    -0.01790535, -0.01851635, -0.01825742, -0.01835702, -0.01809856, 
    -0.01867015, -0.01818208, -0.01879715, -0.01874234, -0.01857389, 
    -0.01823998, -0.01816704, -0.01808944, -0.01813729, -0.0183712, 
    -0.01840984, -0.01857798, -0.01862467, -0.01875426, -0.01886227, 
    -0.01876355, -0.01866047, -0.01837111, -0.01811448, -0.01783911, 
    -0.01777242, -0.0174576, -0.01771337, -0.0172934, -0.01764967, 
    -0.01703792, -0.01815428, -0.01766035, -0.01856628, -0.01846632, 
    -0.01828695, -0.0178827, -0.01809976, -0.01784621, -0.01841136, 
    -0.01871213, -0.01879086, -0.01893862, -0.01878749, -0.01879974, 
    -0.01865624, -0.01870223, -0.01836159, -0.01854373, -0.01803136, 
    -0.01784821, -0.01734182, -0.01703908, -0.01673686, -0.01660528, 
    -0.01656546, -0.01654884,
  -0.05392879, -0.05288604, -0.0530871, -0.05225819, -0.05271635, 
    -0.05217599, -0.05371569, -0.05284504, -0.05339914, -0.0538341, 
    -0.05068813, -0.05222154, -0.04914599, -0.05008706, -0.04775852, 
    -0.04929113, -0.04745567, -0.04780213, -0.04676764, -0.04706157, 
    -0.04576404, -0.04663264, -0.04510658, -0.04596996, -0.04583371, 
    -0.04666157, -0.05190917, -0.05087638, -0.05197102, -0.05182223, 
    -0.05188896, -0.0527068, -0.05312401, -0.05400945, -0.05384757, 
    -0.05319784, -0.05175547, -0.05224048, -0.05102742, -0.05105449, 
    -0.04973809, -0.05032713, -0.04816814, -0.04877164, -0.04704926, 
    -0.04747625, -0.04706921, -0.04719226, -0.0470676, -0.04769551, 
    -0.0474254, -0.04798193, -0.05021623, -0.04954835, -0.05156849, 
    -0.05282469, -0.05367717, -0.05429079, -0.0542036, -0.05403776, 
    -0.05319406, -0.05241357, -0.05182686, -0.05143826, -0.05105838, 
    -0.04992617, -0.04933792, -0.04804701, -0.0482774, -0.04788786, 
    -0.04751896, -0.04690623, -0.04700652, -0.0467386, -0.04789817, 
    -0.04712413, -0.04840914, -0.04805402, -0.05095523, -0.05210918, 
    -0.05260764, -0.05304838, -0.05413665, -0.0533826, -0.05367852, 
    -0.05297742, -0.05253691, -0.05275431, -0.05142767, -0.05193919, 
    -0.04930329, -0.05042091, -0.04756183, -0.04823003, -0.04740315, 
    -0.04782321, -0.04710582, -0.04775095, -0.04663933, -0.04640089, 
    -0.04656368, -0.04594174, -0.04778698, -0.04706917, -0.0527604, 
    -0.05272487, -0.05255973, -0.05328974, -0.05333477, -0.05401387, 
    -0.0534092, -0.05315384, -0.05251152, -0.05213538, -0.05178047, 
    -0.05100908, -0.05016184, -0.04900206, -0.04818641, -0.04764771, 
    -0.0479773, -0.04768619, -0.04801172, -0.04816513, -0.04649006, 
    -0.04742287, -0.04603065, -0.04610655, -0.04673224, -0.046098, 
    -0.05269995, -0.05290463, -0.05362168, -0.05305966, -0.05408838, 
    -0.05350994, -0.05318026, -0.05192836, -0.05165759, -0.05140772, 
    -0.05091806, -0.0502968, -0.04922621, -0.04831436, -0.0474976, 
    -0.04755696, -0.04753605, -0.04735541, -0.04780415, -0.04728216, 
    -0.04719511, -0.04742302, -0.04611673, -0.04648599, -0.04610817, 
    -0.04634821, -0.05283801, -0.05249456, -0.05267985, -0.05233197, 
    -0.05257677, -0.05149732, -0.05117825, -0.04971287, -0.05030893, 
    -0.04936392, -0.0502121, -0.05006067, -0.04933325, -0.0501659, 
    -0.0483641, -0.0495779, -0.0473484, -0.04853339, -0.04727516, 
    -0.04750111, -0.04712767, -0.04679581, -0.0463819, -0.04562822, 
    -0.04580159, -0.04517883, -0.05198694, -0.05154944, -0.05158788, 
    -0.05113389, -0.05080083, -0.05008687, -0.04896375, -0.04938296, 
    -0.04861632, -0.04846391, -0.04962982, -0.04891044, -0.05125887, 
    -0.05087145, -0.0511018, -0.05195225, -0.04928592, -0.05063571, 
    -0.04817304, -0.04888215, -0.04684297, -0.04784552, -0.04589732, 
    -0.04509013, -0.04434449, -0.04348934, -0.05131239, -0.05160779, 
    -0.0510802, -0.05035948, -0.04970058, -0.04883857, -0.04875131, 
    -0.04859186, -0.04818151, -0.04783929, -0.0485415, -0.04775392, 
    -0.05078189, -0.0491706, -0.05171987, -0.05093776, -0.0504017, 
    -0.05063619, -0.04943113, -0.04915152, -0.04803238, -0.04860755, 
    -0.04528788, -0.04672594, -0.04285018, -0.04389763, -0.05171141, 
    -0.05131344, -0.0499533, -0.05059566, -0.04878163, -0.0483457, 
    -0.04799443, -0.04754922, -0.04750146, -0.04724003, -0.04766923, 
    -0.04725693, -0.04883675, -0.04812397, -0.05010691, -0.04961641, 
    -0.04984145, -0.05008948, -0.04932813, -0.04853034, -0.04851355, 
    -0.04826071, -0.0475555, -0.04877442, -0.04510553, -0.04733514, 
    -0.05088316, -0.05013224, -0.05002608, -0.0503149, -0.04838922, 
    -0.04907779, -0.0472464, -0.04773413, -0.04693778, -0.04733172, 
    -0.04738997, -0.04790176, -0.04822332, -0.04904597, -0.04972629, 
    -0.05027292, -0.05014525, -0.04954675, -0.04848201, -0.04749709, 
    -0.047711, -0.04699781, -0.04891081, -0.04809874, -0.04841087, 
    -0.04760149, -0.04939412, -0.04786285, -0.04979375, -0.04962122, 
    -0.04909156, -0.04804411, -0.04781575, -0.04757299, -0.04772265, 
    -0.04845532, -0.04857653, -0.04910439, -0.04925114, -0.04965874, 
    -0.04999884, -0.04968798, -0.0493637, -0.04845505, -0.04765129, 
    -0.04679109, -0.04658313, -0.04560323, -0.04639909, -0.04509341, 
    -0.04620073, -0.04430184, -0.04777583, -0.04623395, -0.04906764, 
    -0.04875374, -0.04819123, -0.04692712, -0.04760527, -0.04681325, 
    -0.0485813, -0.04952618, -0.04977395, -0.05023948, -0.04976336, 
    -0.0498019, -0.04935039, -0.04949502, -0.04842519, -0.04899679, 
    -0.0473914, -0.04681948, -0.04524364, -0.04430543, -0.04337175, 
    -0.04296617, -0.04284354, -0.04279238,
  -0.07870831, -0.07705726, -0.07737544, -0.07606426, -0.0767888, 
    -0.07593434, -0.07837072, -0.0769924, -0.0778694, -0.07855829, 
    -0.07358485, -0.07600633, -0.07115486, -0.07263708, -0.06897327, 
    -0.07138334, -0.06849768, -0.06904177, -0.06741803, -0.06787911, 
    -0.06584527, -0.06720632, -0.06481629, -0.06616777, -0.06595436, 
    -0.0672517, -0.07551263, -0.07388186, -0.07561037, -0.07537525, 
    -0.0754807, -0.0767737, -0.07743385, -0.07883612, -0.07857963, 
    -0.07755072, -0.07526978, -0.07603627, -0.07412019, -0.0741629, 
    -0.0720872, -0.07301552, -0.06961685, -0.0705658, -0.06785981, 
    -0.06852999, -0.06789111, -0.0680842, -0.0678886, -0.06887429, 
    -0.06845015, -0.06932423, -0.07284068, -0.07178835, -0.07497443, 
    -0.07696021, -0.0783097, -0.07928204, -0.07914381, -0.07888098, 
    -0.07754473, -0.07630993, -0.07538258, -0.07476875, -0.07416904, 
    -0.07238355, -0.071457, -0.06942651, -0.0697886, -0.06917644, 
    -0.06859704, -0.06763541, -0.06779274, -0.06737249, -0.06919263, 
    -0.06797729, -0.0699957, -0.06943751, -0.07400628, -0.07582872, 
    -0.07661686, -0.07731415, -0.0790377, -0.07784322, -0.07831183, 
    -0.07720187, -0.07650498, -0.07684885, -0.07475204, -0.07556006, 
    -0.07140247, -0.0731634, -0.06866436, -0.06971414, -0.06841522, 
    -0.06907488, -0.06794855, -0.06896137, -0.06721681, -0.066843, 
    -0.06709821, -0.06612355, -0.06901795, -0.06789105, -0.07685848, 
    -0.07680228, -0.07654107, -0.0776962, -0.07776748, -0.07884313, 
    -0.07788532, -0.07748107, -0.07646483, -0.07587013, -0.07530928, 
    -0.07409124, -0.07275495, -0.07092833, -0.06964558, -0.06879922, 
    -0.06931695, -0.06885965, -0.06937104, -0.06961212, -0.06698278, 
    -0.06844617, -0.06626283, -0.06638175, -0.0673625, -0.06636833, 
    -0.07676285, -0.07708667, -0.07822181, -0.077332, -0.07896121, 
    -0.07804485, -0.0775229, -0.07554296, -0.07511516, -0.07472054, 
    -0.07394759, -0.0729677, -0.07128113, -0.0698467, -0.06856351, 
    -0.06865671, -0.06862388, -0.06834027, -0.06904495, -0.0682253, 
    -0.06808869, -0.06844641, -0.06639769, -0.06697641, -0.06638428, 
    -0.06676042, -0.07698127, -0.076438, -0.07673106, -0.07618091, 
    -0.07656802, -0.07486203, -0.07435826, -0.07204748, -0.07298683, 
    -0.07149792, -0.07283417, -0.07259548, -0.07144965, -0.07276134, 
    -0.0699249, -0.07183488, -0.06832927, -0.07019109, -0.06821431, 
    -0.06856901, -0.06798284, -0.06746221, -0.06681323, -0.0656326, 
    -0.06590407, -0.06492931, -0.07563553, -0.07494435, -0.07500505, 
    -0.07428822, -0.07376263, -0.07263678, -0.07086805, -0.0715279, 
    -0.07032149, -0.07008183, -0.07191665, -0.07078417, -0.07448553, 
    -0.07387406, -0.07423758, -0.0755807, -0.07137513, -0.07350216, 
    -0.06962456, -0.07073966, -0.06753618, -0.06910992, -0.06605398, 
    -0.06479055, -0.06362492, -0.06228983, -0.07457002, -0.0750365, 
    -0.07420348, -0.07306654, -0.07202812, -0.07067109, -0.07053381, 
    -0.07028303, -0.06963786, -0.06910013, -0.07020383, -0.06896602, 
    -0.07373277, -0.0711936, -0.07521355, -0.0739787, -0.0731331, 
    -0.07350291, -0.07160375, -0.07116356, -0.06940351, -0.07030769, 
    -0.06509994, -0.06735264, -0.0612932, -0.06292703, -0.07520017, 
    -0.07457168, -0.07242629, -0.07343898, -0.07058151, -0.06989598, 
    -0.06934388, -0.06864456, -0.06856958, -0.06815917, -0.06883302, 
    -0.0681857, -0.07066823, -0.06954744, -0.07266837, -0.07189553, 
    -0.07225004, -0.0726409, -0.07144158, -0.07018628, -0.07015988, 
    -0.06976236, -0.06865444, -0.07057017, -0.06481466, -0.06830847, 
    -0.07389253, -0.07270829, -0.07254098, -0.07299623, -0.06996439, 
    -0.07104751, -0.06816917, -0.06893495, -0.0676849, -0.06830309, 
    -0.06839453, -0.06919828, -0.06970359, -0.07099743, -0.07206861, 
    -0.07293005, -0.07272881, -0.07178582, -0.07011028, -0.06856271, 
    -0.06889863, -0.06777907, -0.07078476, -0.0695078, -0.06999843, 
    -0.06872664, -0.07154548, -0.06913716, -0.07217488, -0.07190312, 
    -0.07106919, -0.06942195, -0.06906316, -0.06868188, -0.06891692, 
    -0.07006831, -0.07025892, -0.07108938, -0.07132037, -0.07196221, 
    -0.07249804, -0.07200826, -0.07149757, -0.0700679, -0.06880485, 
    -0.06745481, -0.0671287, -0.0655935, -0.06684019, -0.0647957, 
    -0.06652933, -0.06355829, -0.06900047, -0.06658137, -0.07103154, 
    -0.07053763, -0.06965316, -0.0676682, -0.06873257, -0.06748958, 
    -0.07026642, -0.07175343, -0.07214368, -0.07287733, -0.072127, 
    -0.07218774, -0.07147662, -0.07170435, -0.07002094, -0.07092004, 
    -0.06839678, -0.06749935, -0.06503069, -0.06356389, -0.0621064, 
    -0.06147398, -0.06128285, -0.06120312,
  -0.08618347, -0.08427344, -0.08464142, -0.08312535, -0.08396298, 
    -0.08297516, -0.08579281, -0.08419843, -0.0852128, -0.08600986, 
    -0.08026095, -0.08305837, -0.0774569, -0.07916689, -0.07494235, 
    -0.07772041, -0.07439454, -0.07502125, -0.07315145, -0.07368224, 
    -0.07134189, -0.07290778, -0.07015882, -0.07171282, -0.07146736, 
    -0.07296, -0.08248776, -0.08060391, -0.08260073, -0.08232902, 
    -0.08245087, -0.08394553, -0.08470899, -0.08633139, -0.08603456, 
    -0.08484415, -0.08220714, -0.08309298, -0.08087911, -0.08092845, 
    -0.07853236, -0.07960367, -0.07568386, -0.07677766, -0.07366001, 
    -0.07443175, -0.07369605, -0.07391837, -0.07369316, -0.07482832, 
    -0.07433979, -0.07534669, -0.07940187, -0.07818758, -0.08186588, 
    -0.08416121, -0.08572221, -0.08684752, -0.08668753, -0.08638331, 
    -0.08483724, -0.08340934, -0.08233748, -0.08162826, -0.08093555, 
    -0.07887431, -0.07780537, -0.07546453, -0.07588179, -0.07517641, 
    -0.07450897, -0.07340168, -0.07358281, -0.07309903, -0.07519505, 
    -0.07379529, -0.07612047, -0.07547721, -0.0807476, -0.08285309, 
    -0.08376419, -0.08457053, -0.0865647, -0.08518251, -0.08572468, 
    -0.08444066, -0.08363482, -0.08403243, -0.08160896, -0.08254259, 
    -0.07774247, -0.07977438, -0.07458651, -0.07579597, -0.07429956, 
    -0.07505939, -0.07376219, -0.07492863, -0.07291985, -0.07248967, 
    -0.07278335, -0.07166196, -0.07499382, -0.07369599, -0.08404357, 
    -0.08397858, -0.08367655, -0.08501244, -0.08509489, -0.0863395, 
    -0.08523121, -0.08476359, -0.08358841, -0.08290094, -0.08225279, 
    -0.0808457, -0.07930292, -0.07719567, -0.07571696, -0.07474184, 
    -0.0753383, -0.07481146, -0.07540062, -0.07567841, -0.07265051, 
    -0.07433522, -0.07182217, -0.07195897, -0.07308754, -0.07194354, 
    -0.08393298, -0.08430745, -0.08562052, -0.08459117, -0.08647616, 
    -0.08541577, -0.08481197, -0.08252282, -0.08202848, -0.08157256, 
    -0.0806798, -0.07954848, -0.07760251, -0.07594875, -0.07447036, 
    -0.07457769, -0.07453988, -0.07421325, -0.07502491, -0.07408086, 
    -0.07392354, -0.07433549, -0.0719773, -0.07264318, -0.07196187, 
    -0.07239465, -0.08418556, -0.0835574, -0.08389623, -0.08326018, 
    -0.08370771, -0.08173603, -0.08115409, -0.07848654, -0.07957056, 
    -0.07785257, -0.07939436, -0.07911889, -0.0777969, -0.07931029, 
    -0.07603887, -0.07824127, -0.07420059, -0.0763457, -0.0740682, 
    -0.07447669, -0.07380167, -0.07320231, -0.07245541, -0.07109731, 
    -0.07140951, -0.07028873, -0.08262981, -0.08183113, -0.08190126, 
    -0.08107319, -0.08046622, -0.07916654, -0.07712615, -0.07788714, 
    -0.07649601, -0.07621974, -0.0783356, -0.07702943, -0.08130109, 
    -0.08059489, -0.0810147, -0.08256644, -0.07771094, -0.08016548, 
    -0.07569274, -0.0769781, -0.07328745, -0.07509977, -0.07158194, 
    -0.07012925, -0.06878988, -0.06725694, -0.08139869, -0.0819376, 
    -0.08097532, -0.07966258, -0.0784642, -0.07689905, -0.07674078, 
    -0.07645167, -0.07570808, -0.07508849, -0.07636037, -0.07493399, 
    -0.08043175, -0.07750157, -0.08214217, -0.08071573, -0.07973941, 
    -0.08016634, -0.07797462, -0.07746693, -0.07543802, -0.0764801, 
    -0.07048488, -0.07307618, -0.06611338, -0.06798842, -0.08212671, 
    -0.0814006, -0.07892363, -0.08009252, -0.07679576, -0.07600553, 
    -0.07536931, -0.0745637, -0.07447734, -0.07400471, -0.07478078, 
    -0.07403526, -0.07689575, -0.07560387, -0.07920299, -0.07831123, 
    -0.07872024, -0.07917129, -0.07778757, -0.07634015, -0.07630972, 
    -0.07585155, -0.0745751, -0.0767827, -0.07015696, -0.07417665, 
    -0.08061621, -0.07924908, -0.07905598, -0.07958141, -0.07608438, 
    -0.07733309, -0.07401622, -0.07489821, -0.07345866, -0.07417043, 
    -0.07427573, -0.07520156, -0.07578382, -0.07727535, -0.07851092, 
    -0.07950501, -0.07927274, -0.07818467, -0.07625255, -0.07446943, 
    -0.07485636, -0.07356707, -0.07703011, -0.07555819, -0.07612362, 
    -0.07465825, -0.07790742, -0.07513117, -0.07863352, -0.07831998, 
    -0.07735809, -0.07545927, -0.07504588, -0.07460669, -0.07487743, 
    -0.07620417, -0.07642388, -0.07738137, -0.07764778, -0.07838815, 
    -0.07900643, -0.07844128, -0.07785216, -0.07620369, -0.07474834, 
    -0.07319379, -0.07281844, -0.07105237, -0.07248644, -0.07013517, 
    -0.07212877, -0.06871337, -0.07497368, -0.07218864, -0.07731467, 
    -0.07674518, -0.07572571, -0.07343943, -0.07466508, -0.07323381, 
    -0.07643252, -0.0781473, -0.07859753, -0.07944418, -0.07857829, 
    -0.07864836, -0.077828, -0.07809068, -0.07614957, -0.07718609, 
    -0.07427833, -0.07324505, -0.07040527, -0.0687198, -0.0670464, 
    -0.06632076, -0.0661015, -0.06601005,
  -0.06731972, -0.06577227, -0.0660704, -0.06484208, -0.06552074, 
    -0.06472041, -0.06700322, -0.0657115, -0.06653332, -0.06717906, 
    -0.06252129, -0.06478783, -0.06024928, -0.06163482, -0.05821183, 
    -0.0604628, -0.05776796, -0.05827576, -0.05676073, -0.05719081, 
    -0.05529455, -0.0565633, -0.05433598, -0.05559508, -0.0553962, 
    -0.0566056, -0.06432551, -0.06279916, -0.06441703, -0.06419689, 
    -0.06429562, -0.0655066, -0.06612515, -0.06743955, -0.06719907, 
    -0.06623465, -0.06409815, -0.06481586, -0.06302214, -0.06306211, 
    -0.06112069, -0.06198872, -0.05881265, -0.05969891, -0.0571728, 
    -0.0577981, -0.057202, -0.05738214, -0.05719965, -0.05811943, -0.0577236, 
    -0.05853945, -0.06182522, -0.06084133, -0.06382164, -0.06568135, 
    -0.06694602, -0.06785768, -0.06772807, -0.06748162, -0.06622905, 
    -0.06507218, -0.06420375, -0.06362912, -0.06306786, -0.06139776, 
    -0.06053163, -0.05863493, -0.05897302, -0.05840148, -0.05786068, 
    -0.05696348, -0.05711024, -0.05671826, -0.05841658, -0.05728241, 
    -0.05916642, -0.0586452, -0.06291559, -0.0646215, -0.06535968, 
    -0.06601297, -0.06762857, -0.06650878, -0.06694802, -0.06590775, 
    -0.06525487, -0.065577, -0.06361348, -0.06436993, -0.06048067, 
    -0.06212704, -0.0579235, -0.05890349, -0.057691, -0.05830666, 
    -0.05725559, -0.05820071, -0.05657308, -0.05622452, -0.05646248, 
    -0.05555387, -0.05825353, -0.05720195, -0.06558603, -0.06553337, 
    -0.06528867, -0.06637099, -0.0664378, -0.06744613, -0.06654824, 
    -0.06616938, -0.06521726, -0.06466027, -0.06413513, -0.06299506, 
    -0.06174504, -0.06003761, -0.05883947, -0.05804936, -0.05853265, 
    -0.05810577, -0.05858315, -0.05880823, -0.05635485, -0.05771989, 
    -0.05568368, -0.05579451, -0.05670895, -0.05578202, -0.06549643, 
    -0.06579982, -0.06686363, -0.06602969, -0.06755684, -0.06669775, 
    -0.06620858, -0.06435391, -0.06395338, -0.06358399, -0.06286065, 
    -0.061944, -0.06036727, -0.05902728, -0.05782939, -0.05791636, 
    -0.05788572, -0.05762107, -0.05827872, -0.0575138, -0.05738633, 
    -0.05772011, -0.05580937, -0.0563489, -0.05579687, -0.05614752, 
    -0.06570107, -0.06519213, -0.06546665, -0.06495133, -0.06531392, 
    -0.06371644, -0.06324494, -0.06108356, -0.06196189, -0.06056988, 
    -0.06181912, -0.06159592, -0.06052477, -0.06175101, -0.05910031, 
    -0.06088483, -0.0576108, -0.05934892, -0.05750354, -0.05783452, 
    -0.05728757, -0.05680194, -0.05619676, -0.05509637, -0.05534932, 
    -0.05444123, -0.06444059, -0.0637935, -0.06385031, -0.06317939, 
    -0.06268759, -0.06163453, -0.05998129, -0.06059789, -0.05947071, 
    -0.05924686, -0.06096125, -0.05990292, -0.06336404, -0.06279185, 
    -0.063132, -0.06438926, -0.06045512, -0.06244392, -0.05881985, 
    -0.05986133, -0.05687092, -0.05833938, -0.05548903, -0.05431202, 
    -0.05322686, -0.05198491, -0.06344312, -0.06387975, -0.06310008, 
    -0.06203645, -0.06106545, -0.05979728, -0.05966903, -0.05943478, 
    -0.05883227, -0.05833024, -0.05936081, -0.05820506, -0.06265967, 
    -0.06028548, -0.0640455, -0.06288976, -0.0620987, -0.06244462, 
    -0.06066877, -0.06025741, -0.05861346, -0.05945782, -0.05460016, 
    -0.05669975, -0.05105847, -0.05257753, -0.06403297, -0.06344466, 
    -0.06143771, -0.06238481, -0.05971359, -0.05907329, -0.05855778, 
    -0.05790503, -0.05783504, -0.05745209, -0.05808091, -0.05747684, 
    -0.0597946, -0.05874784, -0.06166407, -0.06094151, -0.06127292, 
    -0.06163838, -0.06051721, -0.05934442, -0.05931976, -0.05894852, 
    -0.05791427, -0.059703, -0.05433448, -0.05759142, -0.06280912, 
    -0.06170142, -0.06154495, -0.06197068, -0.05913718, -0.06014897, 
    -0.05746142, -0.05817606, -0.05700964, -0.05758637, -0.05767169, 
    -0.05842186, -0.05889364, -0.06010218, -0.06110331, -0.06190878, 
    -0.06172058, -0.06083897, -0.05927344, -0.05782864, -0.05814215, 
    -0.05709749, -0.05990347, -0.05871083, -0.05916897, -0.05798163, 
    -0.06061432, -0.05836483, -0.06120265, -0.0609486, -0.06016922, 
    -0.05863068, -0.05829572, -0.05793986, -0.05815922, -0.05923424, 
    -0.05941226, -0.06018808, -0.06040395, -0.06100384, -0.0615048, 
    -0.06104689, -0.06056955, -0.05923385, -0.05805463, -0.05679503, 
    -0.05649091, -0.05505996, -0.05622191, -0.05431682, -0.05593212, 
    -0.05316487, -0.05823722, -0.05598062, -0.06013404, -0.05967261, 
    -0.05884656, -0.05699407, -0.05798716, -0.05682747, -0.05941926, 
    -0.06080869, -0.06117349, -0.06185949, -0.06115789, -0.06121467, 
    -0.06054997, -0.06076281, -0.05919, -0.06002986, -0.0576738, -0.05683657, 
    -0.05453566, -0.05317007, -0.05181434, -0.05122647, -0.05104884, 
    -0.05097475,
  -0.06391447, -0.06222166, -0.06254755, -0.06120564, -0.06194681, 
    -0.06107282, -0.06356799, -0.06215525, -0.0630538, -0.06376047, 
    -0.05867587, -0.06114641, -0.05620678, -0.0577116, -0.0539992, 
    -0.05643849, -0.05351913, -0.05406837, -0.05243093, -0.05289538, 
    -0.05084988, -0.05221782, -0.04981819, -0.05117367, -0.05095939, 
    -0.05226349, -0.0606419, -0.05897837, -0.06074176, -0.0605016, 
    -0.06060929, -0.06193136, -0.06260741, -0.06404568, -0.06378238, 
    -0.06272715, -0.0603939, -0.06117702, -0.05922118, -0.05926472, 
    -0.05715287, -0.05809643, -0.05464952, -0.05560982, -0.05287593, 
    -0.05355172, -0.05290747, -0.0531021, -0.05290494, -0.05389924, 
    -0.05347117, -0.05435374, -0.05791861, -0.05684945, -0.06009239, 
    -0.0621223, -0.06350538, -0.0645037, -0.0643617, -0.06409176, 
    -0.06272102, -0.06145686, -0.06050907, -0.05988252, -0.05927098, 
    -0.05745393, -0.05651321, -0.0544571, -0.0548232, -0.05420442, 
    -0.05361939, -0.05264986, -0.05280836, -0.05238508, -0.05422076, 
    -0.05299434, -0.0550327, -0.05446822, -0.05910514, -0.06096487, 
    -0.06177086, -0.06248477, -0.0642527, -0.06302696, -0.06350757, 
    -0.06236975, -0.06165637, -0.06200828, -0.05986547, -0.06069036, 
    -0.05645789, -0.05824688, -0.05368733, -0.05474789, -0.05343593, 
    -0.05410181, -0.05296537, -0.05398717, -0.05222838, -0.0518523, 
    -0.05210903, -0.05112926, -0.05404432, -0.05290742, -0.06201814, 
    -0.06196061, -0.06169329, -0.06287625, -0.06294931, -0.06405289, 
    -0.06307013, -0.06265578, -0.0616153, -0.06100719, -0.06043423, 
    -0.05919169, -0.05783143, -0.05597714, -0.05467856, -0.05382345, 
    -0.05434638, -0.05388446, -0.05440104, -0.05464473, -0.05199289, 
    -0.05346716, -0.05126915, -0.05138862, -0.05237504, -0.05137514, 
    -0.06192025, -0.06225177, -0.06341521, -0.06250305, -0.06417414, 
    -0.0632337, -0.06269864, -0.06067289, -0.06023603, -0.05983333, 
    -0.05904532, -0.05804779, -0.05633481, -0.05488196, -0.05358555, 
    -0.0536796, -0.05364647, -0.05336033, -0.05407158, -0.05324438, 
    -0.05310663, -0.0534674, -0.05140464, -0.05198648, -0.05139116, 
    -0.05176925, -0.06214385, -0.06158786, -0.06188772, -0.06132491, 
    -0.06172087, -0.0599777, -0.05946387, -0.05711254, -0.05806725, 
    -0.05655472, -0.05791198, -0.05766932, -0.05650576, -0.05783793, 
    -0.05496107, -0.05689669, -0.05334923, -0.05523045, -0.0532333, 
    -0.05359109, -0.05299992, -0.05247543, -0.05182235, -0.05063646, 
    -0.05090889, -0.04993139, -0.06076746, -0.0600617, -0.06012364, 
    -0.05939246, -0.0588569, -0.05771129, -0.05591604, -0.05658513, 
    -0.05536243, -0.05511985, -0.05697969, -0.05583104, -0.05959363, 
    -0.05897041, -0.05934083, -0.06071145, -0.05643016, -0.05859167, 
    -0.05465731, -0.05578594, -0.05254991, -0.05413722, -0.0510594, 
    -0.04979242, -0.04862646, -0.04729465, -0.0596798, -0.06015574, 
    -0.05930608, -0.05814834, -0.05709287, -0.05571648, -0.05557742, 
    -0.05532349, -0.05467076, -0.05412732, -0.05524332, -0.05399187, 
    -0.05882651, -0.05624605, -0.06033648, -0.05907702, -0.05821606, 
    -0.05859243, -0.05666208, -0.05621559, -0.05443385, -0.05534846, 
    -0.05010237, -0.05236511, -0.04630303, -0.0479298, -0.06032282, 
    -0.05968148, -0.05749736, -0.05852734, -0.05562573, -0.05493181, 
    -0.05437358, -0.05366734, -0.05359167, -0.0531777, -0.05385758, 
    -0.05320444, -0.05571358, -0.05457934, -0.0577434, -0.05695825, 
    -0.05731827, -0.05771548, -0.05649755, -0.05522557, -0.05519884, 
    -0.05479667, -0.05367734, -0.05561425, -0.04981658, -0.05332828, 
    -0.05898922, -0.05778401, -0.05761391, -0.05807681, -0.05500102, 
    -0.05609793, -0.05318778, -0.0539605, -0.05269971, -0.05332283, 
    -0.05341506, -0.05422647, -0.05473723, -0.05604718, -0.05713399, 
    -0.05800948, -0.05780485, -0.05684688, -0.05514865, -0.05358474, 
    -0.05392382, -0.05279458, -0.05583163, -0.05453927, -0.05503546, 
    -0.05375019, -0.05660297, -0.05416476, -0.05724192, -0.05696594, 
    -0.05611991, -0.05445249, -0.05408997, -0.05370501, -0.05394229, 
    -0.05510618, -0.05529909, -0.05614037, -0.05637461, -0.05702594, 
    -0.05757027, -0.05707271, -0.05655436, -0.05510575, -0.05382914, 
    -0.05246797, -0.05213971, -0.05059725, -0.05184948, -0.04979759, 
    -0.05153696, -0.04855993, -0.05402667, -0.05158925, -0.05608174, 
    -0.0555813, -0.05468624, -0.05268289, -0.05375617, -0.05250299, 
    -0.05530667, -0.056814, -0.05721024, -0.05795588, -0.05719329, 
    -0.05725498, -0.0565331, -0.05676418, -0.05505824, -0.05596872, 
    -0.05341733, -0.05251282, -0.05003298, -0.04856551, -0.04711195, 
    -0.04648273, -0.04629274, -0.04621351,
  -0.04035198, -0.03907359, -0.03931955, -0.03830725, -0.03886621, 
    -0.03820712, -0.04009016, -0.03902347, -0.03970177, -0.0402356, 
    -0.03640241, -0.03826259, -0.03454811, -0.03567765, -0.03289467, 
    -0.03472191, -0.0325357, -0.03294641, -0.03172283, -0.03206963, 
    -0.03054395, -0.03156378, -0.02977613, -0.03078516, -0.03062552, 
    -0.03159786, -0.03788236, -0.03662992, -0.0379576, -0.03777665, 
    -0.03785779, -0.03885455, -0.03936473, -0.04045115, -0.04025215, 
    -0.03945512, -0.03769551, -0.03828567, -0.0368126, -0.03684536, 
    -0.03525804, -0.0359668, -0.03338129, -0.03410057, -0.03205509, 
    -0.03256006, -0.03207865, -0.03222404, -0.03207676, -0.03281991, 
    -0.03249985, -0.03315991, -0.03583318, -0.03503027, -0.03746841, 
    -0.03899861, -0.04004287, -0.0407974, -0.04069003, -0.04048597, 
    -0.0394505, -0.03849666, -0.03778228, -0.03731038, -0.03685007, 
    -0.03548411, -0.03477797, -0.03323727, -0.03351131, -0.03304819, 
    -0.03261065, -0.03188627, -0.03200463, -0.03168861, -0.03306041, 
    -0.03214354, -0.03366819, -0.03324559, -0.03672529, -0.03812575, 
    -0.03873348, -0.03927216, -0.04060763, -0.0396815, -0.04004452, 
    -0.03918534, -0.03864712, -0.03891259, -0.03729754, -0.03791887, 
    -0.03473647, -0.03607988, -0.03266144, -0.03345493, -0.0324735, 
    -0.03297142, -0.0321219, -0.03288567, -0.03157166, -0.03129108, 
    -0.0314826, -0.03075207, -0.03292842, -0.03207862, -0.03892003, 
    -0.03887662, -0.03867497, -0.0395677, -0.03962287, -0.04045659, 
    -0.0397141, -0.03940124, -0.03861614, -0.03815764, -0.03772589, 
    -0.03679041, -0.03576767, -0.03437591, -0.03340303, -0.03276323, 
    -0.03315441, -0.03280886, -0.03319531, -0.03337771, -0.03139596, 
    -0.03249685, -0.03085631, -0.03094536, -0.03168111, -0.03093531, 
    -0.03884617, -0.03909631, -0.03997475, -0.03928595, -0.04054824, 
    -0.03983764, -0.0394336, -0.03790571, -0.0375766, -0.03727334, 
    -0.03668029, -0.03593025, -0.03464414, -0.03355532, -0.03258535, 
    -0.03265566, -0.03263089, -0.032417, -0.03294881, -0.03233036, 
    -0.03222743, -0.03249703, -0.03095729, -0.03139117, -0.03094725, 
    -0.03122914, -0.03901487, -0.03859545, -0.03882163, -0.03839717, 
    -0.03869577, -0.03738204, -0.03699523, -0.03522776, -0.03594487, 
    -0.03480911, -0.0358282, -0.03564588, -0.03477238, -0.03577255, 
    -0.03361456, -0.03506573, -0.03240871, -0.03381631, -0.03232207, 
    -0.0325895, -0.03214771, -0.03175604, -0.03126875, -0.03038502, 
    -0.0305879, -0.02986032, -0.03797697, -0.0374453, -0.03749195, 
    -0.03694149, -0.03653856, -0.03567741, -0.03433011, -0.03483192, 
    -0.03391519, -0.03373347, -0.03512803, -0.03426639, -0.0370929, 
    -0.03662394, -0.03690264, -0.03793476, -0.03471566, -0.03633909, 
    -0.03338712, -0.03423258, -0.03181165, -0.03299791, -0.03070002, 
    -0.02975696, -0.02889069, -0.02790317, -0.03715776, -0.03751612, 
    -0.03687648, -0.03600582, -0.03521299, -0.03418051, -0.03407629, 
    -0.03388602, -0.03339719, -0.03299051, -0.03382596, -0.03288919, 
    -0.0365157, -0.03457757, -0.03765226, -0.03670414, -0.03605671, 
    -0.03633966, -0.03488967, -0.03455472, -0.03321987, -0.03390472, 
    -0.02998751, -0.0316737, -0.02716934, -0.02837385, -0.03764197, 
    -0.03715903, -0.03551672, -0.03629072, -0.03411249, -0.03359264, 
    -0.03317476, -0.0326465, -0.03258992, -0.03228053, -0.03278875, 
    -0.03230051, -0.03417834, -0.03332876, -0.03570153, -0.03511194, 
    -0.03538223, -0.03568055, -0.03476622, -0.03381266, -0.03379264, 
    -0.03349145, -0.03265397, -0.03410389, -0.02977493, -0.03239306, 
    -0.03663808, -0.03573204, -0.03560426, -0.03595205, -0.03364447, 
    -0.03446649, -0.03228806, -0.03286572, -0.03192349, -0.03238898, 
    -0.03245791, -0.03306468, -0.03344695, -0.03442843, -0.03524387, 
    -0.03590146, -0.0357477, -0.03502835, -0.03375505, -0.03258475, 
    -0.03283829, -0.03199434, -0.03426683, -0.03329876, -0.03367027, 
    -0.03270845, -0.03484531, -0.03301851, -0.0353249, -0.03511771, 
    -0.03448297, -0.03323382, -0.03296256, -0.03267466, -0.0328521, 
    -0.03372323, -0.03386774, -0.03449832, -0.034674, -0.03516275, 
    -0.03557148, -0.03519786, -0.03480884, -0.03372291, -0.03276749, 
    -0.03175048, -0.03150549, -0.03035583, -0.03128898, -0.02976081, 
    -0.03105594, -0.02884131, -0.03291522, -0.03109493, -0.03445435, 
    -0.03407919, -0.03340878, -0.03191093, -0.03271292, -0.03177662, 
    -0.03387342, -0.03500367, -0.03530111, -0.03586118, -0.03528839, 
    -0.0353347, -0.03479289, -0.03496628, -0.03368732, -0.03436961, 
    -0.03245961, -0.03178396, -0.02993588, -0.02884545, -0.02776788, 
    -0.02730223, -0.02716173, -0.02710316,
  -0.01970498, -0.01870054, -0.01889315, -0.01810236, -0.01853836, 
    -0.01802443, -0.01949861, -0.01866132, -0.0191931, -0.01961321, 
    -0.01662923, -0.0180676, -0.01521544, -0.01607415, -0.01397336, 
    -0.01534705, -0.01370618, -0.01401194, -0.01310463, -0.01336067, 
    -0.01224115, -0.0129875, -0.01168477, -0.01241693, -0.01230054, 
    -0.01301258, -0.01777204, -0.01680411, -0.01783047, -0.01769001, 
    -0.01775297, -0.01852925, -0.01892857, -0.01978323, -0.01962626, 
    -0.01899946, -0.01762709, -0.01808556, -0.01694474, -0.01696998, 
    -0.01575423, -0.01629523, -0.01433699, -0.01487744, -0.01334993, 
    -0.01372429, -0.01336735, -0.01347497, -0.01336595, -0.01391764, 
    -0.01367955, -0.01417136, -0.016193, -0.01558102, -0.01745117, 
    -0.01864188, -0.01946137, -0.02005681, -0.01997192, -0.01981072, 
    -0.01899583, -0.01824993, -0.01769438, -0.01732891, -0.01697361, 
    -0.01592645, -0.01538954, -0.0142292, -0.01443443, -0.0140879, 
    -0.01376189, -0.01322518, -0.01331261, -0.01307941, -0.01409703, 
    -0.01341536, -0.01455215, -0.01423542, -0.01687751, -0.01796114, 
    -0.01843468, -0.01885602, -0.0199068, -0.01917717, -0.01946267, 
    -0.01878802, -0.01836728, -0.01857461, -0.01731899, -0.01780039, 
    -0.01535808, -0.01638183, -0.01379967, -0.01439216, -0.01365998, 
    -0.0140306, -0.01339934, -0.01396665, -0.0129933, -0.01278713, 
    -0.01292779, -0.01239279, -0.01399853, -0.01336732, -0.01858043, 
    -0.0185465, -0.01838901, -0.0190878, -0.01913112, -0.01978753, 
    -0.01920278, -0.0189572, -0.01834311, -0.01798595, -0.01765065, 
    -0.01692765, -0.01614293, -0.01508524, -0.01435328, -0.01387542, 
    -0.01416725, -0.0139094, -0.01419783, -0.01433431, -0.01286412, 
    -0.01367732, -0.01246887, -0.01253393, -0.01307388, -0.01252659, 
    -0.01852271, -0.01871832, -0.01940775, -0.01886683, -0.01985989, 
    -0.01929989, -0.01898258, -0.01779017, -0.01753494, -0.01730028, 
    -0.01684286, -0.01626726, -0.01528814, -0.01446743, -0.01374308, 
    -0.01379537, -0.01377694, -0.01361804, -0.01401373, -0.01355376, 
    -0.01347748, -0.01367746, -0.01254266, -0.0128606, -0.01253532, 
    -0.0127417, -0.01865459, -0.01832696, -0.01850353, -0.01817239, 
    -0.01840525, -0.01738434, -0.01708553, -0.01573118, -0.01627845, 
    -0.01541315, -0.0161892, -0.01604989, -0.0153853, -0.01614666, 
    -0.01451188, -0.01560796, -0.01361189, -0.01466344, -0.01354762, 
    -0.01374616, -0.01341845, -0.01312911, -0.01277074, -0.01212558, 
    -0.01227314, -0.01174553, -0.01784551, -0.01743328, -0.01746939, 
    -0.01704408, -0.01673384, -0.01607397, -0.01505064, -0.01543046, 
    -0.01473782, -0.01460118, -0.01565532, -0.01500252, -0.0171609, 
    -0.01679951, -0.01701413, -0.01781273, -0.01534232, -0.01658061, 
    -0.01434136, -0.014977, -0.01317011, -0.01405037, -0.01235483, 
    -0.01167095, -0.01104943, -0.01034922, -0.01721098, -0.0174881, 
    -0.01699397, -0.0163251, -0.01571995, -0.01493772, -0.01485914, 
    -0.01471587, -0.0143489, -0.01404485, -0.0146707, -0.01396927, 
    -0.01671627, -0.01523773, -0.01759356, -0.01686122, -0.01636408, 
    -0.01658105, -0.01547426, -0.01522044, -0.01421619, -0.01472995, 
    -0.01183745, -0.01306842, -0.009834968, -0.01068182, -0.01758559, 
    -0.01721196, -0.01595132, -0.01654349, -0.01488643, -0.01449544, 
    -0.01418246, -0.01378855, -0.01374648, -0.01351682, -0.01389443, 
    -0.01353163, -0.01493608, -0.01429766, -0.0160924, -0.01564309, 
    -0.0158488, -0.01607637, -0.01538063, -0.0146607, -0.01464565, 
    -0.01441954, -0.01379411, -0.01487995, -0.0116839, -0.01360027, 
    -0.01681039, -0.0161157, -0.01601812, -0.01628395, -0.01453434, 
    -0.0151537, -0.0135224, -0.01395178, -0.01325267, -0.01359724, 
    -0.0136484, -0.01410022, -0.01438618, -0.01512493, -0.01574344, 
    -0.01624523, -0.01612766, -0.01557956, -0.01461739, -0.01374263, 
    -0.01393133, -0.01330501, -0.01500286, -0.01427521, -0.01455371, 
    -0.01383464, -0.01544061, -0.01406575, -0.01580513, -0.01564748, 
    -0.01516616, -0.01422662, -0.014024, -0.0138095, -0.01394163, 
    -0.01459348, -0.01470212, -0.01517777, -0.01531075, -0.01568172, 
    -0.0159931, -0.01570843, -0.01541295, -0.01459324, -0.01387859, 
    -0.01312501, -0.01294462, -0.01210438, -0.01278559, -0.01167372, 
    -0.01261482, -0.01101419, -0.01398868, -0.01264336, -0.01514452, 
    -0.01486133, -0.01435758, -0.0132434, -0.01383797, -0.01314428, 
    -0.01470639, -0.01556082, -0.01578701, -0.01621442, -0.01577733, 
    -0.0158126, -0.01540086, -0.01553242, -0.01456652, -0.01508047, 
    -0.01364966, -0.01314969, -0.01180012, -0.01101715, -0.01025401, 
    -0.009927695, -0.009829662, -0.009788851,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  296.8234, 298.0832, 297.838, 298.8564, 298.2913, 298.9585, 297.0786, 
    298.1332, 297.4597, 296.9368, 300.8316, 298.9019, 302.843, 301.6074, 
    304.7191, 302.6503, 305.1329, 304.6596, 306.0789, 305.6729, 307.4884, 
    306.2665, 308.4333, 307.1964, 307.3895, 306.2262, 299.2915, 300.5913, 
    299.2141, 299.4002, 299.3167, 298.3029, 297.7927, 296.7275, 296.9207, 
    297.7033, 299.4839, 298.8787, 300.4007, 300.3664, 302.0624, 301.2968, 
    304.1588, 303.3433, 305.6899, 305.1053, 305.6624, 305.4934, 305.6646, 
    304.8063, 305.1745, 304.4131, 301.44, 302.3113, 299.7183, 298.1577, 
    297.1248, 296.3932, 296.4966, 296.6935, 297.7079, 298.6643, 299.3947, 
    299.8819, 300.3615, 301.8159, 302.5886, 304.3238, 304.0103, 304.5417, 
    305.0472, 305.887, 305.7487, 306.119, 304.5278, 305.5866, 303.8318, 
    304.3145, 300.4909, 299.0419, 298.4243, 297.8851, 296.576, 297.4795, 
    297.1231, 297.9719, 298.512, 298.2448, 299.8952, 299.254, 302.6344, 
    301.1757, 304.9889, 304.0746, 305.2049, 304.6308, 305.6119, 304.7301, 
    306.2571, 306.5897, 306.3623, 307.2367, 304.6805, 305.6622, 298.2373, 
    298.2809, 298.4839, 297.5919, 297.5374, 296.7221, 297.4476, 297.7568, 
    298.5434, 299.0093, 299.4527, 300.4238, 301.5103, 303.0348, 304.134, 
    304.8724, 304.4195, 304.8193, 304.3724, 304.1631, 306.4649, 305.1779, 
    307.1108, 307.0036, 306.1278, 307.0157, 298.3115, 298.0608, 297.1915, 
    297.8716, 296.6335, 297.3259, 297.7245, 299.2672, 299.607, 299.9201, 
    300.5396, 301.3359, 302.7368, 303.9599, 305.0763, 304.9956, 305.024, 
    305.2701, 304.6569, 305.3702, 305.4893, 305.1778, 306.9893, 306.4709, 
    307.0014, 306.6638, 298.1423, 298.5643, 298.3362, 298.7652, 298.4628, 
    299.8073, 300.2091, 302.0951, 301.3202, 302.5544, 301.4455, 301.6417, 
    302.5943, 301.5054, 303.8922, 302.272, 305.2796, 303.6629, 305.3798, 
    305.0716, 305.5821, 306.0398, 306.6165, 307.6826, 307.4355, 308.3289, 
    299.1944, 299.7421, 299.6942, 300.2657, 300.6889, 301.6078, 303.0861, 
    302.5296, 303.5521, 303.7576, 302.2046, 303.1572, 300.1075, 300.5984, 
    300.3062, 299.2375, 302.6575, 300.8996, 304.1521, 303.1952, 305.9745, 
    304.5997, 307.2995, 308.4567, 309.5498, 310.83, 300.0402, 299.6693, 
    300.3338, 301.2547, 302.1116, 303.2535, 303.3706, 303.5849, 304.1408, 
    304.6087, 303.6525, 304.726, 300.712, 302.8106, 299.5287, 300.514, 
    301.2004, 300.8993, 302.4661, 302.8362, 304.3438, 303.5639, 308.1706, 
    306.1362, 311.808, 310.2148, 299.5396, 300.039, 301.7812, 300.9513, 
    303.3299, 303.9176, 304.3961, 305.0059, 305.071, 305.4278, 304.8427, 
    305.4048, 303.2559, 304.2191, 301.5819, 302.222, 301.9275, 301.6045, 
    302.6021, 303.6675, 303.6906, 304.0328, 304.9958, 303.3396, 308.4333, 
    305.2962, 300.5841, 301.5484, 301.6867, 301.3127, 303.8586, 302.9342, 
    305.4191, 304.7533, 305.8435, 305.3025, 305.2229, 304.5229, 304.0838, 
    302.9764, 302.0779, 301.367, 301.5322, 302.3135, 303.7328, 305.0768, 
    304.7848, 305.7607, 303.157, 304.2533, 303.8291, 304.9351, 302.5148, 
    304.5748, 301.9898, 302.2159, 302.9158, 304.3275, 304.641, 304.9736, 
    304.7691, 303.769, 303.6055, 302.8989, 302.7039, 302.1667, 301.7223, 
    302.1282, 302.5548, 303.7695, 304.8672, 306.0462, 306.3354, 307.7175, 
    306.5916, 308.4508, 306.8689, 309.6116, 304.695, 306.8231, 302.9478, 
    303.3674, 304.127, 305.8576, 304.9299, 306.0152, 303.5991, 302.3403, 
    302.0157, 301.4101, 302.0295, 301.9792, 302.5727, 302.3819, 303.8099, 
    303.0422, 305.2208, 306.0067, 308.2351, 309.6071, 311.0092, 311.6295, 
    311.8185, 311.8976 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.357484e-08, 6.385439e-08, 6.380004e-08, 6.402553e-08, 6.390044e-08, 
    6.404809e-08, 6.363151e-08, 6.386549e-08, 6.371612e-08, 6.360001e-08, 
    6.446311e-08, 6.403558e-08, 6.490716e-08, 6.463451e-08, 6.53194e-08, 
    6.486473e-08, 6.541108e-08, 6.530627e-08, 6.562168e-08, 6.553132e-08, 
    6.593476e-08, 6.566339e-08, 6.614388e-08, 6.586995e-08, 6.59128e-08, 
    6.565443e-08, 6.412161e-08, 6.440989e-08, 6.410453e-08, 6.414565e-08, 
    6.41272e-08, 6.390303e-08, 6.379007e-08, 6.355347e-08, 6.359642e-08, 
    6.377019e-08, 6.416413e-08, 6.40304e-08, 6.436741e-08, 6.43598e-08, 
    6.473498e-08, 6.456582e-08, 6.519642e-08, 6.501719e-08, 6.553509e-08, 
    6.540485e-08, 6.552898e-08, 6.549134e-08, 6.552947e-08, 6.533845e-08, 
    6.542029e-08, 6.52522e-08, 6.459751e-08, 6.478992e-08, 6.421605e-08, 
    6.387099e-08, 6.364178e-08, 6.347913e-08, 6.350213e-08, 6.354596e-08, 
    6.377121e-08, 6.398299e-08, 6.414438e-08, 6.425233e-08, 6.43587e-08, 
    6.46807e-08, 6.48511e-08, 6.523266e-08, 6.516379e-08, 6.528045e-08, 
    6.539189e-08, 6.557899e-08, 6.55482e-08, 6.563063e-08, 6.527737e-08, 
    6.551215e-08, 6.512457e-08, 6.523057e-08, 6.438765e-08, 6.406648e-08, 
    6.392999e-08, 6.38105e-08, 6.351981e-08, 6.372055e-08, 6.364142e-08, 
    6.382967e-08, 6.39493e-08, 6.389013e-08, 6.425529e-08, 6.411333e-08, 
    6.48612e-08, 6.453907e-08, 6.537889e-08, 6.517793e-08, 6.542706e-08, 
    6.529993e-08, 6.551776e-08, 6.532171e-08, 6.566131e-08, 6.573526e-08, 
    6.568472e-08, 6.587883e-08, 6.531085e-08, 6.552898e-08, 6.388848e-08, 
    6.389813e-08, 6.394308e-08, 6.374548e-08, 6.373339e-08, 6.355229e-08, 
    6.371343e-08, 6.378205e-08, 6.395624e-08, 6.405927e-08, 6.415721e-08, 
    6.437256e-08, 6.461306e-08, 6.494936e-08, 6.519095e-08, 6.53529e-08, 
    6.525359e-08, 6.534127e-08, 6.524326e-08, 6.519733e-08, 6.570755e-08, 
    6.542106e-08, 6.585091e-08, 6.582712e-08, 6.563259e-08, 6.582981e-08, 
    6.390491e-08, 6.384938e-08, 6.365659e-08, 6.380746e-08, 6.353257e-08, 
    6.368644e-08, 6.377492e-08, 6.41163e-08, 6.41913e-08, 6.426085e-08, 
    6.43982e-08, 6.457448e-08, 6.488371e-08, 6.515276e-08, 6.539837e-08, 
    6.538038e-08, 6.538671e-08, 6.544158e-08, 6.530567e-08, 6.546389e-08, 
    6.549045e-08, 6.542102e-08, 6.582394e-08, 6.570883e-08, 6.582662e-08, 
    6.575167e-08, 6.386743e-08, 6.396086e-08, 6.391037e-08, 6.400531e-08, 
    6.393843e-08, 6.423585e-08, 6.432501e-08, 6.474225e-08, 6.457101e-08, 
    6.484353e-08, 6.459869e-08, 6.464208e-08, 6.485244e-08, 6.461192e-08, 
    6.513793e-08, 6.478133e-08, 6.544371e-08, 6.508762e-08, 6.546603e-08, 
    6.539731e-08, 6.551109e-08, 6.561299e-08, 6.574118e-08, 6.597772e-08, 
    6.592295e-08, 6.612076e-08, 6.410015e-08, 6.422134e-08, 6.421067e-08, 
    6.433749e-08, 6.443128e-08, 6.463457e-08, 6.496062e-08, 6.483801e-08, 
    6.506309e-08, 6.510828e-08, 6.476632e-08, 6.497628e-08, 6.430245e-08, 
    6.441132e-08, 6.434649e-08, 6.410971e-08, 6.486627e-08, 6.447801e-08, 
    6.519495e-08, 6.498462e-08, 6.559846e-08, 6.529319e-08, 6.589279e-08, 
    6.614913e-08, 6.639036e-08, 6.667229e-08, 6.428748e-08, 6.420513e-08, 
    6.435257e-08, 6.455657e-08, 6.474583e-08, 6.499745e-08, 6.502319e-08, 
    6.507033e-08, 6.519242e-08, 6.529509e-08, 6.508524e-08, 6.532083e-08, 
    6.443658e-08, 6.489997e-08, 6.4174e-08, 6.439262e-08, 6.454454e-08, 
    6.44779e-08, 6.482399e-08, 6.490557e-08, 6.523705e-08, 6.506569e-08, 
    6.608587e-08, 6.563452e-08, 6.688694e-08, 6.653695e-08, 6.417636e-08, 
    6.428719e-08, 6.467292e-08, 6.448939e-08, 6.501424e-08, 6.514343e-08, 
    6.524845e-08, 6.538271e-08, 6.53972e-08, 6.547674e-08, 6.53464e-08, 
    6.547159e-08, 6.499798e-08, 6.520963e-08, 6.462883e-08, 6.47702e-08, 
    6.470516e-08, 6.463382e-08, 6.485399e-08, 6.508855e-08, 6.509355e-08, 
    6.516876e-08, 6.538072e-08, 6.501637e-08, 6.614414e-08, 6.544767e-08, 
    6.440805e-08, 6.462153e-08, 6.465201e-08, 6.456932e-08, 6.513049e-08, 
    6.492716e-08, 6.54748e-08, 6.532679e-08, 6.55693e-08, 6.544879e-08, 
    6.543107e-08, 6.527629e-08, 6.517993e-08, 6.493648e-08, 6.473839e-08, 
    6.458131e-08, 6.461784e-08, 6.479039e-08, 6.51029e-08, 6.539852e-08, 
    6.533376e-08, 6.555087e-08, 6.497619e-08, 6.521717e-08, 6.512403e-08, 
    6.536688e-08, 6.483475e-08, 6.528791e-08, 6.471893e-08, 6.476881e-08, 
    6.492312e-08, 6.523352e-08, 6.530218e-08, 6.53755e-08, 6.533025e-08, 
    6.511083e-08, 6.507487e-08, 6.491937e-08, 6.487644e-08, 6.475795e-08, 
    6.465985e-08, 6.474948e-08, 6.48436e-08, 6.511091e-08, 6.535181e-08, 
    6.561444e-08, 6.567871e-08, 6.598559e-08, 6.573578e-08, 6.614802e-08, 
    6.579756e-08, 6.640422e-08, 6.531416e-08, 6.578724e-08, 6.493014e-08, 
    6.502248e-08, 6.518949e-08, 6.557254e-08, 6.536574e-08, 6.560759e-08, 
    6.507346e-08, 6.479635e-08, 6.472464e-08, 6.459086e-08, 6.472769e-08, 
    6.471657e-08, 6.48475e-08, 6.480542e-08, 6.511979e-08, 6.495092e-08, 
    6.543063e-08, 6.560568e-08, 6.610003e-08, 6.640308e-08, 6.671156e-08, 
    6.684775e-08, 6.68892e-08, 6.690653e-08 ;

 SOM_C_LEACHED =
  4.887949e-20, -5.476003e-20, -2.83453e-20, 4.010503e-21, -3.068273e-21, 
    -2.686305e-20, 1.660543e-20, 5.183759e-20, 8.246297e-21, -6.252845e-21, 
    -5.037543e-20, -3.63907e-20, -3.403394e-20, -4.144622e-20, 1.522268e-20, 
    1.989003e-20, -2.196207e-20, -7.771551e-20, 3.61981e-22, 8.374906e-20, 
    8.510362e-20, 3.600625e-22, 9.415408e-21, -1.235119e-19, -3.870513e-20, 
    -1.174637e-20, 3.741559e-20, -7.533419e-21, -5.874145e-20, 5.186635e-20, 
    1.419277e-20, 3.094447e-20, -9.036269e-21, 1.76617e-20, 3.147943e-20, 
    4.016613e-20, 2.89712e-21, 6.438378e-20, 4.990581e-21, 2.928121e-20, 
    -3.754243e-20, -4.955224e-20, 7.29246e-20, -1.81893e-20, 4.070844e-20, 
    -6.052358e-20, 1.386919e-20, -7.046415e-20, -3.892646e-21, -1.667877e-20, 
    2.252856e-21, 9.655536e-21, -6.802784e-20, 4.585479e-21, -4.128332e-20, 
    2.906953e-20, -1.95061e-20, -2.344152e-20, -6.992234e-21, -5.946788e-20, 
    1.62008e-20, -7.889739e-20, 1.824867e-20, 2.556382e-20, -3.47742e-21, 
    -4.870982e-20, -4.910719e-20, 5.895402e-20, -9.357565e-20, -2.467978e-20, 
    3.380025e-20, 4.417665e-20, 3.799082e-20, -1.328042e-20, -1.817947e-20, 
    -2.458276e-20, 3.835964e-20, -6.263518e-21, 2.91531e-20, -1.969907e-20, 
    2.21151e-20, 2.312829e-21, -3.55326e-20, -6.366651e-20, 4.980995e-20, 
    3.303848e-20, -7.149312e-20, 2.128834e-20, 1.824491e-20, -4.251213e-20, 
    -3.846727e-20, 6.68254e-20, 5.097931e-20, -2.493963e-20, -3.875258e-21, 
    -2.920529e-20, -1.920486e-21, 2.862985e-20, -4.281699e-20, -1.235165e-20, 
    8.091319e-20, -3.480049e-20, -1.444186e-20, -2.12188e-20, 8.147318e-21, 
    1.690571e-20, -4.229542e-21, 2.998889e-20, -3.886879e-20, 8.420063e-20, 
    -5.445758e-20, 8.563336e-21, -3.654602e-20, 2.850773e-20, -1.287444e-20, 
    5.600885e-20, 3.823339e-20, -2.560838e-20, -9.159649e-20, 7.301193e-21, 
    -1.197522e-20, -3.960556e-21, 2.152507e-20, 3.815034e-20, 3.493224e-20, 
    -6.26781e-20, 2.0945e-20, 1.37984e-20, 2.46643e-20, 3.15408e-20, 
    3.462566e-20, -4.778415e-21, 3.233882e-20, -1.733824e-20, 4.612486e-20, 
    -1.062799e-20, -3.059459e-20, 5.839649e-21, -2.725919e-20, 8.415558e-20, 
    5.375985e-20, -6.259959e-20, -3.390862e-20, -8.118199e-21, 2.378198e-20, 
    -1.872176e-20, 4.97189e-20, -4.835428e-20, -5.789356e-20, 3.330422e-21, 
    8.745703e-21, -6.167397e-22, 2.291095e-22, 1.427401e-20, -4.551848e-20, 
    -6.260594e-21, -2.916638e-21, 2.539956e-20, 3.516103e-20, -7.372494e-21, 
    3.097053e-20, 4.243502e-20, 4.95359e-21, 1.50018e-20, 3.833981e-21, 
    2.071968e-21, 5.425549e-21, -2.887593e-20, 3.659444e-20, -1.501169e-20, 
    -1.395215e-20, 7.75523e-20, -1.012113e-20, -6.041346e-20, -1.216795e-20, 
    5.264768e-20, 3.673522e-20, 4.899914e-20, -1.220133e-20, -4.365536e-20, 
    2.140084e-20, -3.466208e-20, 2.723099e-20, -1.631687e-20, -1.385572e-20, 
    -1.737551e-20, -8.962816e-21, -1.66315e-20, 2.100649e-20, 3.570785e-20, 
    1.028667e-20, -2.772572e-20, 8.309171e-21, 3.091598e-20, -2.724806e-20, 
    3.929374e-20, -3.535225e-20, 5.427066e-20, 4.195767e-21, -8.163412e-21, 
    3.125688e-20, -8.923902e-20, -5.942076e-20, -9.723117e-21, -2.946989e-20, 
    -3.193372e-20, -2.028688e-20, -3.159316e-20, 3.500381e-20, -1.999898e-20, 
    -1.677525e-20, 5.957222e-20, -2.277433e-20, 3.316598e-20, 5.739845e-21, 
    -5.567857e-20, -5.975283e-20, 2.488331e-20, -6.279382e-21, -2.29639e-20, 
    -5.922664e-20, 8.829133e-20, 5.480649e-20, 7.964235e-20, -5.867716e-21, 
    3.656962e-20, 1.517981e-20, 4.929643e-20, -6.230083e-21, 1.238183e-20, 
    1.140453e-20, 2.068306e-20, 2.58046e-21, 2.86536e-20, -1.091748e-19, 
    -4.708939e-21, -1.33068e-20, -2.941628e-20, 1.728351e-20, -4.738223e-21, 
    1.424161e-20, -2.232234e-20, -1.592083e-20, 1.793136e-20, -2.402293e-20, 
    1.259581e-20, 1.323337e-20, 2.699384e-20, 3.00741e-20, -4.683159e-20, 
    6.897048e-20, 2.157327e-20, 3.219616e-20, -1.772899e-20, -3.945079e-20, 
    1.05684e-19, -2.223598e-20, -4.911028e-21, 1.149049e-19, 5.18453e-20, 
    -2.608253e-20, -4.672852e-20, -1.076185e-20, -5.977739e-21, 5.53099e-20, 
    -2.612201e-21, -2.693962e-20, 1.877151e-21, -2.933541e-20, -7.236351e-21, 
    -1.542372e-20, -3.238278e-20, -4.200418e-20, 4.941256e-20, -5.043964e-20, 
    1.667019e-20, 3.604947e-20, -5.182012e-20, 1.693447e-20, -1.330087e-20, 
    5.182486e-20, 8.83483e-20, 2.525955e-21, 1.873117e-20, -3.569233e-20, 
    -1.429228e-21, 3.112471e-21, 1.991299e-20, 1.203659e-20, 6.387845e-21, 
    4.167287e-20, -8.989901e-21, 2.562716e-20, -5.547451e-20, 5.300113e-20, 
    6.608241e-20, 3.766674e-20, 5.493633e-20, -5.941181e-20, -5.863934e-20, 
    5.315291e-21, 4.237484e-21, -5.984115e-20, -3.215916e-21, 7.920039e-21, 
    3.485043e-20, 1.815891e-20, 4.602636e-20, 6.194392e-20, -3.769548e-20, 
    3.880114e-20, 7.71703e-21, 4.255706e-20, -2.144052e-20, 1.095242e-20, 
    -3.664954e-20, -4.403486e-20, -1.426652e-20, 2.36827e-20, -2.113285e-20, 
    5.880754e-20, -6.027657e-20, 1.812145e-21, -2.596402e-20, -2.142309e-20, 
    4.094303e-20, -2.151247e-21, 1.705521e-20, 1.392472e-20, 7.751489e-21, 
    -3.113971e-20, -2.666007e-20, -2.937998e-20, -4.000667e-20, 2.335482e-20, 
    -1.513648e-21, -1.399694e-20, 2.81515e-20 ;

 SR =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371698e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441075e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379093e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377207e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523353e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.56315e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529406e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.532169e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547246e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.46224e-08, 6.465288e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532766e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472856e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999936, 0.9999937, 0.9999937, 
    0.9999937, 0.9999936, 0.9999934, 0.9999935, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999936, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 0.9999936, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999937, 0.9999936, 0.9999937, 
    0.9999936, 0.9999936, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999937, 0.9999936, 
    0.9999937, 0.9999937, 0.9999936, 0.9999937, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999937, 0.9999937, 0.9999937, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999935, 0.9999935, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999937, 0.9999937, 
    0.9999937, 0.9999937, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999935, 0.9999935, 0.9999935, 0.9999934, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999937, 0.9999937, 0.9999937, 0.9999937, 0.9999935, 0.9999934, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 0.9999936, 
    0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999936, 0.9999938, 0.9999937, 
    0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999935, 0.9999936, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999937, 0.9999936, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 
    0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999937, 0.9999937, 0.9999937, 0.9999937, 0.9999937, 
    0.9999936, 0.9999937, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999937, 0.9999938, 0.9999938, 
    0.9999938, 0.9999938 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.1477094, -0.1477245, -0.1477216, -0.1477333, -0.147727, -0.1477344, 
    -0.1477125, -0.147725, -0.1477171, -0.1477109, -0.1477537, -0.1477338, 
    -0.1477685, -0.1477599, -0.1477925, -0.1477671, -0.1477954, -0.1477923, 
    -0.1478021, -0.1477993, -0.1478115, -0.1478034, -0.1478181, -0.1478097, 
    -0.1478109, -0.1478031, -0.1477383, -0.1477517, -0.1477374, -0.1477394, 
    -0.1477386, -0.1477271, -0.1477208, -0.1477084, -0.1477107, -0.1477199, 
    -0.1477403, -0.1477337, -0.1477508, -0.1477504, -0.1477632, -0.1477577, 
    -0.1477889, -0.147772, -0.1477994, -0.1477954, -0.1477992, -0.1477981, 
    -0.1477992, -0.1477933, -0.1477958, -0.1477906, -0.1477587, -0.147765, 
    -0.147743, -0.147725, -0.1477131, -0.1477043, -0.1477056, -0.1477079, 
    -0.1477199, -0.1477313, -0.1477395, -0.1477449, -0.1477503, -0.1477611, 
    -0.1477668, -0.1477899, -0.1477879, -0.1477914, -0.147795, -0.1478007, 
    -0.1477998, -0.1478023, -0.1477914, -0.1477986, -0.1477753, -0.14779, 
    -0.1477509, -0.1477355, -0.1477282, -0.1477221, -0.1477065, -0.1477172, 
    -0.147713, -0.1477233, -0.1477296, -0.1477266, -0.1477451, -0.1477379, 
    -0.1477671, -0.1477567, -0.1477946, -0.1477883, -0.1477961, -0.1477921, 
    -0.1477988, -0.1477928, -0.1478033, -0.1478055, -0.147804, -0.1478101, 
    -0.1477925, -0.1477991, -0.1477264, -0.1477269, -0.1477294, -0.1477186, 
    -0.147718, -0.1477083, -0.147717, -0.1477206, -0.14773, -0.1477352, 
    -0.1477401, -0.1477509, -0.1477591, -0.1477698, -0.1477887, -0.1477938, 
    -0.1477907, -0.1477934, -0.1477904, -0.147789, -0.1478046, -0.1477958, 
    -0.1478092, -0.1478085, -0.1478024, -0.1478085, -0.1477273, -0.1477244, 
    -0.1477139, -0.1477221, -0.1477072, -0.1477154, -0.1477201, -0.1477379, 
    -0.1477419, -0.1477453, -0.1477519, -0.147758, -0.1477679, -0.1477875, 
    -0.1477952, -0.1477946, -0.1477948, -0.1477965, -0.1477923, -0.1477972, 
    -0.147798, -0.1477959, -0.1478084, -0.1478048, -0.1478084, -0.1478061, 
    -0.1477253, -0.1477302, -0.1477276, -0.1477324, -0.147729, -0.1477439, 
    -0.1477483, -0.1477633, -0.1477578, -0.1477666, -0.1477588, -0.1477602, 
    -0.1477667, -0.1477592, -0.1477869, -0.1477645, -0.1477966, -0.1477738, 
    -0.1477973, -0.1477952, -0.1477987, -0.1478018, -0.1478058, -0.147813, 
    -0.1478114, -0.1478175, -0.1477373, -0.1477432, -0.1477429, -0.1477492, 
    -0.147753, -0.14776, -0.1477702, -0.1477666, -0.1477734, -0.1477747, 
    -0.1477643, -0.1477707, -0.1477473, -0.1477521, -0.1477496, -0.1477376, 
    -0.1477673, -0.1477546, -0.1477888, -0.147771, -0.1478013, -0.1477918, 
    -0.1478104, -0.1478181, -0.1478259, -0.1478343, -0.1477467, -0.1477426, 
    -0.14775, -0.1477572, -0.1477636, -0.1477713, -0.1477722, -0.1477735, 
    -0.1477888, -0.147792, -0.1477739, -0.1477928, -0.1477528, -0.1477684, 
    -0.1477409, -0.1477514, -0.1477569, -0.1477547, -0.1477662, -0.1477686, 
    -0.1477901, -0.1477735, -0.1478161, -0.1478023, -0.1478412, -0.1478302, 
    -0.1477411, -0.1477467, -0.1477611, -0.1477552, -0.1477719, -0.1477872, 
    -0.1477906, -0.1477946, -0.1477951, -0.1477976, -0.1477936, -0.1477975, 
    -0.1477714, -0.1477893, -0.1477598, -0.1477644, -0.1477623, -0.14776, 
    -0.1477671, -0.147774, -0.1477743, -0.147788, -0.147794, -0.147772, 
    -0.1478176, -0.1477962, -0.1477522, -0.1477593, -0.1477605, -0.1477579, 
    -0.1477754, -0.1477692, -0.1477975, -0.147793, -0.1478005, -0.1477967, 
    -0.1477962, -0.1477914, -0.1477884, -0.1477695, -0.1477633, -0.1477583, 
    -0.1477595, -0.147765, -0.1477744, -0.1477951, -0.1477931, -0.1477999, 
    -0.1477707, -0.1477895, -0.1477751, -0.1477942, -0.1477665, -0.1477912, 
    -0.1477628, -0.1477644, -0.1477691, -0.1477899, -0.1477922, -0.1477944, 
    -0.1477931, -0.1477747, -0.1477737, -0.147769, -0.1477677, -0.1477641, 
    -0.1477608, -0.1477637, -0.1477667, -0.1477748, -0.1477937, -0.1478018, 
    -0.1478039, -0.147813, -0.1478053, -0.1478177, -0.1478068, -0.1478258, 
    -0.1477922, -0.1478069, -0.1477694, -0.1477722, -0.1477885, -0.1478004, 
    -0.1477942, -0.1478015, -0.1477737, -0.1477651, -0.147763, -0.1477585, 
    -0.147763, -0.1477627, -0.1477669, -0.1477656, -0.1477751, -0.14777, 
    -0.1477961, -0.1478015, -0.1478168, -0.1478261, -0.1478358, -0.14784, 
    -0.1478413, -0.1478418 ;

 TAUY =
  -0.1477094, -0.1477245, -0.1477216, -0.1477333, -0.147727, -0.1477344, 
    -0.1477125, -0.147725, -0.1477171, -0.1477109, -0.1477537, -0.1477338, 
    -0.1477685, -0.1477599, -0.1477925, -0.1477671, -0.1477954, -0.1477923, 
    -0.1478021, -0.1477993, -0.1478115, -0.1478034, -0.1478181, -0.1478097, 
    -0.1478109, -0.1478031, -0.1477383, -0.1477517, -0.1477374, -0.1477394, 
    -0.1477386, -0.1477271, -0.1477208, -0.1477084, -0.1477107, -0.1477199, 
    -0.1477403, -0.1477337, -0.1477508, -0.1477504, -0.1477632, -0.1477577, 
    -0.1477889, -0.147772, -0.1477994, -0.1477954, -0.1477992, -0.1477981, 
    -0.1477992, -0.1477933, -0.1477958, -0.1477906, -0.1477587, -0.147765, 
    -0.147743, -0.147725, -0.1477131, -0.1477043, -0.1477056, -0.1477079, 
    -0.1477199, -0.1477313, -0.1477395, -0.1477449, -0.1477503, -0.1477611, 
    -0.1477668, -0.1477899, -0.1477879, -0.1477914, -0.147795, -0.1478007, 
    -0.1477998, -0.1478023, -0.1477914, -0.1477986, -0.1477753, -0.14779, 
    -0.1477509, -0.1477355, -0.1477282, -0.1477221, -0.1477065, -0.1477172, 
    -0.147713, -0.1477233, -0.1477296, -0.1477266, -0.1477451, -0.1477379, 
    -0.1477671, -0.1477567, -0.1477946, -0.1477883, -0.1477961, -0.1477921, 
    -0.1477988, -0.1477928, -0.1478033, -0.1478055, -0.147804, -0.1478101, 
    -0.1477925, -0.1477991, -0.1477264, -0.1477269, -0.1477294, -0.1477186, 
    -0.147718, -0.1477083, -0.147717, -0.1477206, -0.14773, -0.1477352, 
    -0.1477401, -0.1477509, -0.1477591, -0.1477698, -0.1477887, -0.1477938, 
    -0.1477907, -0.1477934, -0.1477904, -0.147789, -0.1478046, -0.1477958, 
    -0.1478092, -0.1478085, -0.1478024, -0.1478085, -0.1477273, -0.1477244, 
    -0.1477139, -0.1477221, -0.1477072, -0.1477154, -0.1477201, -0.1477379, 
    -0.1477419, -0.1477453, -0.1477519, -0.147758, -0.1477679, -0.1477875, 
    -0.1477952, -0.1477946, -0.1477948, -0.1477965, -0.1477923, -0.1477972, 
    -0.147798, -0.1477959, -0.1478084, -0.1478048, -0.1478084, -0.1478061, 
    -0.1477253, -0.1477302, -0.1477276, -0.1477324, -0.147729, -0.1477439, 
    -0.1477483, -0.1477633, -0.1477578, -0.1477666, -0.1477588, -0.1477602, 
    -0.1477667, -0.1477592, -0.1477869, -0.1477645, -0.1477966, -0.1477738, 
    -0.1477973, -0.1477952, -0.1477987, -0.1478018, -0.1478058, -0.147813, 
    -0.1478114, -0.1478175, -0.1477373, -0.1477432, -0.1477429, -0.1477492, 
    -0.147753, -0.14776, -0.1477702, -0.1477666, -0.1477734, -0.1477747, 
    -0.1477643, -0.1477707, -0.1477473, -0.1477521, -0.1477496, -0.1477376, 
    -0.1477673, -0.1477546, -0.1477888, -0.147771, -0.1478013, -0.1477918, 
    -0.1478104, -0.1478181, -0.1478259, -0.1478343, -0.1477467, -0.1477426, 
    -0.14775, -0.1477572, -0.1477636, -0.1477713, -0.1477722, -0.1477735, 
    -0.1477888, -0.147792, -0.1477739, -0.1477928, -0.1477528, -0.1477684, 
    -0.1477409, -0.1477514, -0.1477569, -0.1477547, -0.1477662, -0.1477686, 
    -0.1477901, -0.1477735, -0.1478161, -0.1478023, -0.1478412, -0.1478302, 
    -0.1477411, -0.1477467, -0.1477611, -0.1477552, -0.1477719, -0.1477872, 
    -0.1477906, -0.1477946, -0.1477951, -0.1477976, -0.1477936, -0.1477975, 
    -0.1477714, -0.1477893, -0.1477598, -0.1477644, -0.1477623, -0.14776, 
    -0.1477671, -0.147774, -0.1477743, -0.147788, -0.147794, -0.147772, 
    -0.1478176, -0.1477962, -0.1477522, -0.1477593, -0.1477605, -0.1477579, 
    -0.1477754, -0.1477692, -0.1477975, -0.147793, -0.1478005, -0.1477967, 
    -0.1477962, -0.1477914, -0.1477884, -0.1477695, -0.1477633, -0.1477583, 
    -0.1477595, -0.147765, -0.1477744, -0.1477951, -0.1477931, -0.1477999, 
    -0.1477707, -0.1477895, -0.1477751, -0.1477942, -0.1477665, -0.1477912, 
    -0.1477628, -0.1477644, -0.1477691, -0.1477899, -0.1477922, -0.1477944, 
    -0.1477931, -0.1477747, -0.1477737, -0.147769, -0.1477677, -0.1477641, 
    -0.1477608, -0.1477637, -0.1477667, -0.1477748, -0.1477937, -0.1478018, 
    -0.1478039, -0.147813, -0.1478053, -0.1478177, -0.1478068, -0.1478258, 
    -0.1477922, -0.1478069, -0.1477694, -0.1477722, -0.1477885, -0.1478004, 
    -0.1477942, -0.1478015, -0.1477737, -0.1477651, -0.147763, -0.1477585, 
    -0.147763, -0.1477627, -0.1477669, -0.1477656, -0.1477751, -0.14777, 
    -0.1477961, -0.1478015, -0.1478168, -0.1478261, -0.1478358, -0.14784, 
    -0.1478413, -0.1478418 ;

 TBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.6911, 261.7076, 261.7044, 261.7177, 261.7103, 261.719, 261.6944, 
    261.7082, 261.6994, 261.6926, 261.7435, 261.7183, 261.7699, 261.7537, 
    261.7942, 261.7673, 261.7996, 261.7934, 261.8121, 261.8068, 261.8306, 
    261.8146, 261.843, 261.8268, 261.8293, 261.8141, 261.7234, 261.7403, 
    261.7224, 261.7248, 261.7237, 261.7104, 261.7037, 261.6898, 261.6924, 
    261.7026, 261.7259, 261.718, 261.7379, 261.7375, 261.7597, 261.7497, 
    261.7869, 261.7765, 261.807, 261.7993, 261.8066, 261.8044, 261.8067, 
    261.7953, 261.8002, 261.7903, 261.7516, 261.7629, 261.729, 261.7085, 
    261.695, 261.6854, 261.6868, 261.6894, 261.7027, 261.7152, 261.7248, 
    261.7311, 261.7374, 261.7564, 261.7665, 261.7891, 261.785, 261.7919, 
    261.7985, 261.8096, 261.8078, 261.8127, 261.7917, 261.8056, 261.7828, 
    261.789, 261.739, 261.7201, 261.712, 261.705, 261.6878, 261.6997, 
    261.695, 261.7061, 261.7132, 261.7097, 261.7313, 261.7229, 261.7672, 
    261.7481, 261.7977, 261.7858, 261.8006, 261.7931, 261.806, 261.7944, 
    261.8145, 261.8188, 261.8159, 261.8274, 261.7937, 261.8066, 261.7096, 
    261.7102, 261.7129, 261.7011, 261.7004, 261.6898, 261.6993, 261.7033, 
    261.7136, 261.7197, 261.7255, 261.7382, 261.7524, 261.7724, 261.7866, 
    261.7962, 261.7903, 261.7955, 261.7897, 261.787, 261.8172, 261.8002, 
    261.8257, 261.8243, 261.8128, 261.8245, 261.7106, 261.7073, 261.6959, 
    261.7048, 261.6886, 261.6977, 261.7029, 261.7231, 261.7275, 261.7316, 
    261.7397, 261.7502, 261.7685, 261.7843, 261.7989, 261.7979, 261.7982, 
    261.8015, 261.7934, 261.8028, 261.8044, 261.8002, 261.8241, 261.8173, 
    261.8243, 261.8198, 261.7084, 261.7139, 261.7109, 261.7165, 261.7126, 
    261.7301, 261.7354, 261.7601, 261.75, 261.7661, 261.7516, 261.7542, 
    261.7666, 261.7524, 261.7834, 261.7624, 261.8016, 261.7805, 261.8029, 
    261.7989, 261.8056, 261.8116, 261.8192, 261.8332, 261.83, 261.8417, 
    261.7221, 261.7293, 261.7287, 261.7361, 261.7417, 261.7538, 261.7731, 
    261.7658, 261.7792, 261.7818, 261.7616, 261.774, 261.7341, 261.7405, 
    261.7367, 261.7227, 261.7675, 261.7444, 261.7868, 261.7745, 261.8108, 
    261.7926, 261.8282, 261.8433, 261.8576, 261.8742, 261.7332, 261.7283, 
    261.7371, 261.7491, 261.7603, 261.7753, 261.7768, 261.7796, 261.7867, 
    261.7928, 261.7804, 261.7943, 261.7419, 261.7695, 261.7265, 261.7393, 
    261.7484, 261.7445, 261.765, 261.7698, 261.7893, 261.7793, 261.8395, 
    261.8128, 261.887, 261.8663, 261.7267, 261.7332, 261.756, 261.7451, 
    261.7763, 261.7838, 261.79, 261.7979, 261.7988, 261.8035, 261.7958, 
    261.8033, 261.7753, 261.7877, 261.7534, 261.7618, 261.758, 261.7537, 
    261.7668, 261.7806, 261.781, 261.7853, 261.7977, 261.7764, 261.8429, 
    261.8017, 261.7404, 261.7529, 261.7548, 261.7499, 261.7831, 261.7711, 
    261.8034, 261.7947, 261.809, 261.8019, 261.8008, 261.7917, 261.7859, 
    261.7716, 261.7599, 261.7506, 261.7528, 261.763, 261.7815, 261.7989, 
    261.795, 261.808, 261.774, 261.7881, 261.7827, 261.797, 261.7656, 
    261.7922, 261.7588, 261.7617, 261.7708, 261.7891, 261.7932, 261.7975, 
    261.7949, 261.782, 261.7798, 261.7707, 261.7681, 261.7611, 261.7553, 
    261.7606, 261.7661, 261.782, 261.7961, 261.8117, 261.8155, 261.8336, 
    261.8188, 261.8431, 261.8224, 261.8583, 261.7938, 261.8218, 261.7713, 
    261.7768, 261.7865, 261.8092, 261.797, 261.8112, 261.7798, 261.7633, 
    261.7591, 261.7512, 261.7593, 261.7586, 261.7664, 261.7639, 261.7825, 
    261.7725, 261.8008, 261.8112, 261.8404, 261.8583, 261.8766, 261.8847, 
    261.8871, 261.8882 ;

 TG_R =
  261.6911, 261.7076, 261.7044, 261.7177, 261.7103, 261.719, 261.6944, 
    261.7082, 261.6994, 261.6926, 261.7435, 261.7183, 261.7699, 261.7537, 
    261.7942, 261.7673, 261.7996, 261.7934, 261.8121, 261.8068, 261.8306, 
    261.8146, 261.843, 261.8268, 261.8293, 261.8141, 261.7234, 261.7403, 
    261.7224, 261.7248, 261.7237, 261.7104, 261.7037, 261.6898, 261.6924, 
    261.7026, 261.7259, 261.718, 261.7379, 261.7375, 261.7597, 261.7497, 
    261.7869, 261.7765, 261.807, 261.7993, 261.8066, 261.8044, 261.8067, 
    261.7953, 261.8002, 261.7903, 261.7516, 261.7629, 261.729, 261.7085, 
    261.695, 261.6854, 261.6868, 261.6894, 261.7027, 261.7152, 261.7248, 
    261.7311, 261.7374, 261.7564, 261.7665, 261.7891, 261.785, 261.7919, 
    261.7985, 261.8096, 261.8078, 261.8127, 261.7917, 261.8056, 261.7828, 
    261.789, 261.739, 261.7201, 261.712, 261.705, 261.6878, 261.6997, 
    261.695, 261.7061, 261.7132, 261.7097, 261.7313, 261.7229, 261.7672, 
    261.7481, 261.7977, 261.7858, 261.8006, 261.7931, 261.806, 261.7944, 
    261.8145, 261.8188, 261.8159, 261.8274, 261.7937, 261.8066, 261.7096, 
    261.7102, 261.7129, 261.7011, 261.7004, 261.6898, 261.6993, 261.7033, 
    261.7136, 261.7197, 261.7255, 261.7382, 261.7524, 261.7724, 261.7866, 
    261.7962, 261.7903, 261.7955, 261.7897, 261.787, 261.8172, 261.8002, 
    261.8257, 261.8243, 261.8128, 261.8245, 261.7106, 261.7073, 261.6959, 
    261.7048, 261.6886, 261.6977, 261.7029, 261.7231, 261.7275, 261.7316, 
    261.7397, 261.7502, 261.7685, 261.7843, 261.7989, 261.7979, 261.7982, 
    261.8015, 261.7934, 261.8028, 261.8044, 261.8002, 261.8241, 261.8173, 
    261.8243, 261.8198, 261.7084, 261.7139, 261.7109, 261.7165, 261.7126, 
    261.7301, 261.7354, 261.7601, 261.75, 261.7661, 261.7516, 261.7542, 
    261.7666, 261.7524, 261.7834, 261.7624, 261.8016, 261.7805, 261.8029, 
    261.7989, 261.8056, 261.8116, 261.8192, 261.8332, 261.83, 261.8417, 
    261.7221, 261.7293, 261.7287, 261.7361, 261.7417, 261.7538, 261.7731, 
    261.7658, 261.7792, 261.7818, 261.7616, 261.774, 261.7341, 261.7405, 
    261.7367, 261.7227, 261.7675, 261.7444, 261.7868, 261.7745, 261.8108, 
    261.7926, 261.8282, 261.8433, 261.8576, 261.8742, 261.7332, 261.7283, 
    261.7371, 261.7491, 261.7603, 261.7753, 261.7768, 261.7796, 261.7867, 
    261.7928, 261.7804, 261.7943, 261.7419, 261.7695, 261.7265, 261.7393, 
    261.7484, 261.7445, 261.765, 261.7698, 261.7893, 261.7793, 261.8395, 
    261.8128, 261.887, 261.8663, 261.7267, 261.7332, 261.756, 261.7451, 
    261.7763, 261.7838, 261.79, 261.7979, 261.7988, 261.8035, 261.7958, 
    261.8033, 261.7753, 261.7877, 261.7534, 261.7618, 261.758, 261.7537, 
    261.7668, 261.7806, 261.781, 261.7853, 261.7977, 261.7764, 261.8429, 
    261.8017, 261.7404, 261.7529, 261.7548, 261.7499, 261.7831, 261.7711, 
    261.8034, 261.7947, 261.809, 261.8019, 261.8008, 261.7917, 261.7859, 
    261.7716, 261.7599, 261.7506, 261.7528, 261.763, 261.7815, 261.7989, 
    261.795, 261.808, 261.774, 261.7881, 261.7827, 261.797, 261.7656, 
    261.7922, 261.7588, 261.7617, 261.7708, 261.7891, 261.7932, 261.7975, 
    261.7949, 261.782, 261.7798, 261.7707, 261.7681, 261.7611, 261.7553, 
    261.7606, 261.7661, 261.782, 261.7961, 261.8117, 261.8155, 261.8336, 
    261.8188, 261.8431, 261.8224, 261.8583, 261.7938, 261.8218, 261.7713, 
    261.7768, 261.7865, 261.8092, 261.797, 261.8112, 261.7798, 261.7633, 
    261.7591, 261.7512, 261.7593, 261.7586, 261.7664, 261.7639, 261.7825, 
    261.7725, 261.8008, 261.8112, 261.8404, 261.8583, 261.8766, 261.8847, 
    261.8871, 261.8882 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.0153, 254.0171, 254.0168, 254.0182, 254.0174, 254.0184, 254.0157, 
    254.0172, 254.0162, 254.0155, 254.021, 254.0183, 254.024, 254.0223, 
    254.0267, 254.0237, 254.0273, 254.0267, 254.0288, 254.0282, 254.0308, 
    254.029, 254.0322, 254.0304, 254.0306, 254.029, 254.0189, 254.0207, 
    254.0188, 254.019, 254.0189, 254.0175, 254.0167, 254.0152, 254.0155, 
    254.0166, 254.0192, 254.0183, 254.0205, 254.0205, 254.0229, 254.0218, 
    254.026, 254.0248, 254.0282, 254.0273, 254.0282, 254.0279, 254.0282, 
    254.0269, 254.0274, 254.0263, 254.022, 254.0233, 254.0195, 254.0172, 
    254.0157, 254.0147, 254.0148, 254.0151, 254.0166, 254.018, 254.0191, 
    254.0198, 254.0205, 254.0225, 254.0237, 254.0262, 254.0257, 254.0265, 
    254.0273, 254.0285, 254.0283, 254.0288, 254.0265, 254.028, 254.0255, 
    254.0262, 254.0205, 254.0185, 254.0176, 254.0168, 254.0149, 254.0163, 
    254.0157, 254.017, 254.0178, 254.0174, 254.0198, 254.0189, 254.0237, 
    254.0216, 254.0272, 254.0258, 254.0275, 254.0266, 254.0281, 254.0268, 
    254.029, 254.0295, 254.0292, 254.0305, 254.0267, 254.0281, 254.0174, 
    254.0174, 254.0177, 254.0164, 254.0163, 254.0152, 254.0162, 254.0167, 
    254.0178, 254.0185, 254.0191, 254.0206, 254.0221, 254.0243, 254.0259, 
    254.027, 254.0264, 254.0269, 254.0263, 254.026, 254.0293, 254.0274, 
    254.0303, 254.0301, 254.0288, 254.0301, 254.0175, 254.0171, 254.0158, 
    254.0168, 254.015, 254.016, 254.0166, 254.0188, 254.0194, 254.0198, 
    254.0207, 254.0219, 254.0239, 254.0257, 254.0273, 254.0272, 254.0272, 
    254.0276, 254.0267, 254.0277, 254.0279, 254.0274, 254.0301, 254.0293, 
    254.0301, 254.0296, 254.0172, 254.0179, 254.0175, 254.0181, 254.0177, 
    254.0196, 254.0202, 254.0229, 254.0219, 254.0236, 254.022, 254.0223, 
    254.0236, 254.0221, 254.0255, 254.0232, 254.0276, 254.0252, 254.0277, 
    254.0273, 254.028, 254.0287, 254.0295, 254.0311, 254.0307, 254.032, 
    254.0188, 254.0195, 254.0195, 254.0203, 254.0209, 254.0223, 254.0244, 
    254.0236, 254.0251, 254.0254, 254.0231, 254.0245, 254.0201, 254.0208, 
    254.0204, 254.0188, 254.0238, 254.0212, 254.0259, 254.0246, 254.0286, 
    254.0266, 254.0305, 254.0322, 254.0338, 254.0356, 254.02, 254.0195, 
    254.0204, 254.0217, 254.023, 254.0247, 254.0248, 254.0251, 254.0259, 
    254.0266, 254.0252, 254.0268, 254.0209, 254.024, 254.0192, 254.0206, 
    254.0217, 254.0212, 254.0235, 254.0241, 254.0262, 254.0251, 254.0318, 
    254.0288, 254.0371, 254.0347, 254.0193, 254.02, 254.0225, 254.0213, 
    254.0248, 254.0256, 254.0263, 254.0272, 254.0273, 254.0278, 254.0269, 
    254.0278, 254.0247, 254.026, 254.0222, 254.0232, 254.0228, 254.0223, 
    254.0237, 254.0252, 254.0253, 254.0258, 254.027, 254.0248, 254.0321, 
    254.0275, 254.0208, 254.0222, 254.0224, 254.0219, 254.0255, 254.0242, 
    254.0278, 254.0268, 254.0284, 254.0276, 254.0275, 254.0265, 254.0258, 
    254.0242, 254.0229, 254.0219, 254.0222, 254.0233, 254.0253, 254.0273, 
    254.0268, 254.0283, 254.0245, 254.0261, 254.0255, 254.0271, 254.0236, 
    254.0265, 254.0228, 254.0232, 254.0242, 254.0262, 254.0267, 254.0271, 
    254.0268, 254.0254, 254.0252, 254.0242, 254.0238, 254.0231, 254.0224, 
    254.023, 254.0236, 254.0254, 254.027, 254.0287, 254.0291, 254.0311, 
    254.0294, 254.0321, 254.0298, 254.0338, 254.0267, 254.0298, 254.0242, 
    254.0248, 254.0259, 254.0284, 254.0271, 254.0286, 254.0252, 254.0233, 
    254.0229, 254.022, 254.0229, 254.0228, 254.0237, 254.0234, 254.0255, 
    254.0244, 254.0275, 254.0286, 254.0319, 254.0339, 254.0359, 254.0368, 
    254.0371, 254.0372 ;

 THBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23998, 18.23999, 18.23999, 18.24, 18.23999, 18.23999, 
    18.23997, 18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 
    18.23991, 18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 
    18.23994, 18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 
    18.23991, 18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 
    18.23988, 18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 
    18.23996, 18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 
    18.23993, 18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 
    18.23992, 18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 
    18.23985, 18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 
    18.23993, 18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 
    18.23993, 18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 
    18.23992, 18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 
    18.23996, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 
    18.23994, 18.23994, 18.23995, 18.23994, 18.23992, 18.23992, 18.23992, 
    18.23991, 18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 
    18.23995, 18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23991, 18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 
    18.23994, 18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 
    18.23992, 18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 
    18.23992, 18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 
    18.23993, 18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 
    18.2399, 18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 
    18.23991, 18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 
    18.2399, 18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 
    18.23994, 18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 
    18.23986, 18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTCOLCH4 =
  1.357287e-05, 1.336598e-05, 1.34061e-05, 1.323997e-05, 1.333202e-05, 
    1.32234e-05, 1.353082e-05, 1.335779e-05, 1.346815e-05, 1.355419e-05, 
    1.292026e-05, 1.323258e-05, 1.268327e-05, 1.289255e-05, 1.237232e-05, 
    1.271565e-05, 1.230412e-05, 1.238211e-05, 1.214884e-05, 1.221522e-05, 
    1.192171e-05, 1.211832e-05, 1.17726e-05, 1.196835e-05, 1.193749e-05, 
    1.212486e-05, 1.316945e-05, 1.295894e-05, 1.318197e-05, 1.315184e-05, 
    1.316535e-05, 1.333012e-05, 1.341348e-05, 1.358873e-05, 1.355685e-05, 
    1.342816e-05, 1.31383e-05, 1.323639e-05, 1.298984e-05, 1.299539e-05, 
    1.28151e-05, 1.29457e-05, 1.246436e-05, 1.25996e-05, 1.221244e-05, 
    1.230874e-05, 1.221695e-05, 1.224471e-05, 1.221659e-05, 1.235812e-05, 
    1.229729e-05, 1.242253e-05, 1.292116e-05, 1.277292e-05, 1.310031e-05, 
    1.335375e-05, 1.352321e-05, 1.364397e-05, 1.362687e-05, 1.359431e-05, 
    1.342741e-05, 1.327124e-05, 1.315276e-05, 1.307378e-05, 1.299618e-05, 
    1.285691e-05, 1.272607e-05, 1.243717e-05, 1.248888e-05, 1.24014e-05, 
    1.231836e-05, 1.218015e-05, 1.22028e-05, 1.214228e-05, 1.24037e-05, 
    1.222935e-05, 1.251842e-05, 1.243873e-05, 1.297512e-05, 1.320989e-05, 
    1.331026e-05, 1.339838e-05, 1.361374e-05, 1.346488e-05, 1.352348e-05, 
    1.338422e-05, 1.329603e-05, 1.333962e-05, 1.307163e-05, 1.317552e-05, 
    1.271835e-05, 1.296645e-05, 1.232802e-05, 1.247825e-05, 1.229227e-05, 
    1.238684e-05, 1.222522e-05, 1.237059e-05, 1.211984e-05, 1.206592e-05, 
    1.210274e-05, 1.196195e-05, 1.237869e-05, 1.221695e-05, 1.334084e-05, 
    1.333373e-05, 1.330061e-05, 1.344644e-05, 1.345538e-05, 1.35896e-05, 
    1.347014e-05, 1.34194e-05, 1.329093e-05, 1.321518e-05, 1.314336e-05, 
    1.298609e-05, 1.290912e-05, 1.265112e-05, 1.246846e-05, 1.234735e-05, 
    1.242149e-05, 1.235601e-05, 1.242922e-05, 1.246368e-05, 1.208609e-05, 
    1.229672e-05, 1.198209e-05, 1.199928e-05, 1.214085e-05, 1.199734e-05, 
    1.332873e-05, 1.336968e-05, 1.351224e-05, 1.340062e-05, 1.360425e-05, 
    1.349012e-05, 1.342467e-05, 1.317334e-05, 1.311841e-05, 1.306756e-05, 
    1.296743e-05, 1.293899e-05, 1.270115e-05, 1.249718e-05, 1.231355e-05, 
    1.232692e-05, 1.232221e-05, 1.228151e-05, 1.238256e-05, 1.226499e-05, 
    1.224537e-05, 1.229675e-05, 1.200158e-05, 1.208516e-05, 1.199965e-05, 
    1.205398e-05, 1.335636e-05, 1.328752e-05, 1.33247e-05, 1.325483e-05, 
    1.330404e-05, 1.308583e-05, 1.302074e-05, 1.280951e-05, 1.294167e-05, 
    1.273185e-05, 1.292024e-05, 1.28867e-05, 1.272505e-05, 1.291e-05, 
    1.250835e-05, 1.277951e-05, 1.227993e-05, 1.254631e-05, 1.226341e-05, 
    1.231434e-05, 1.223014e-05, 1.215521e-05, 1.206161e-05, 1.18909e-05, 
    1.19302e-05, 1.178898e-05, 1.318518e-05, 1.309644e-05, 1.310424e-05, 
    1.301164e-05, 1.294337e-05, 1.28925e-05, 1.264256e-05, 1.273608e-05, 
    1.256484e-05, 1.25307e-05, 1.279102e-05, 1.263065e-05, 1.30372e-05, 
    1.295789e-05, 1.300508e-05, 1.317817e-05, 1.271447e-05, 1.290943e-05, 
    1.246546e-05, 1.262432e-05, 1.216586e-05, 1.239188e-05, 1.195189e-05, 
    1.176888e-05, 1.159964e-05, 1.140567e-05, 1.304812e-05, 1.310829e-05, 
    1.300065e-05, 1.295287e-05, 1.280676e-05, 1.261458e-05, 1.259505e-05, 
    1.255937e-05, 1.246735e-05, 1.239046e-05, 1.25481e-05, 1.237126e-05, 
    1.293953e-05, 1.268875e-05, 1.313107e-05, 1.29715e-05, 1.29622e-05, 
    1.290951e-05, 1.27468e-05, 1.268447e-05, 1.243388e-05, 1.256287e-05, 
    1.181375e-05, 1.213944e-05, 1.126087e-05, 1.149826e-05, 1.312934e-05, 
    1.304833e-05, 1.286289e-05, 1.290116e-05, 1.260184e-05, 1.25042e-05, 
    1.242534e-05, 1.232519e-05, 1.231442e-05, 1.225549e-05, 1.23522e-05, 
    1.22593e-05, 1.261417e-05, 1.245444e-05, 1.289693e-05, 1.278805e-05, 
    1.283805e-05, 1.289307e-05, 1.272386e-05, 1.254561e-05, 1.254182e-05, 
    1.248514e-05, 1.232667e-05, 1.260022e-05, 1.177241e-05, 1.2277e-05, 
    1.296027e-05, 1.290258e-05, 1.287902e-05, 1.294298e-05, 1.251396e-05, 
    1.266802e-05, 1.225693e-05, 1.236681e-05, 1.218727e-05, 1.227617e-05, 
    1.22893e-05, 1.240451e-05, 1.247674e-05, 1.266092e-05, 1.281248e-05, 
    1.293369e-05, 1.290543e-05, 1.277256e-05, 1.253477e-05, 1.231344e-05, 
    1.236161e-05, 1.220083e-05, 1.263072e-05, 1.244878e-05, 1.251883e-05, 
    1.233695e-05, 1.273857e-05, 1.239583e-05, 1.282745e-05, 1.278911e-05, 
    1.26711e-05, 1.243653e-05, 1.238517e-05, 1.233054e-05, 1.236422e-05, 
    1.252879e-05, 1.255594e-05, 1.267396e-05, 1.27067e-05, 1.279745e-05, 
    1.287297e-05, 1.280396e-05, 1.27318e-05, 1.252872e-05, 1.234817e-05, 
    1.215414e-05, 1.210713e-05, 1.188527e-05, 1.206553e-05, 1.176967e-05, 
    1.202069e-05, 1.159001e-05, 1.237623e-05, 1.202817e-05, 1.266575e-05, 
    1.25956e-05, 1.246956e-05, 1.218489e-05, 1.23378e-05, 1.215917e-05, 
    1.2557e-05, 1.276799e-05, 1.282306e-05, 1.29263e-05, 1.28207e-05, 
    1.282927e-05, 1.272882e-05, 1.276103e-05, 1.252202e-05, 1.264993e-05, 
    1.228963e-05, 1.216057e-05, 1.180369e-05, 1.159079e-05, 1.137899e-05, 
    1.128712e-05, 1.125936e-05, 1.124778e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23998, 18.23999, 18.23999, 18.24, 18.23999, 18.23999, 
    18.23997, 18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 
    18.23991, 18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 
    18.23994, 18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 
    18.23991, 18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 
    18.23988, 18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 
    18.23996, 18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 
    18.23993, 18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 
    18.23992, 18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 
    18.23985, 18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 
    18.23993, 18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 
    18.23993, 18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 
    18.23992, 18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 
    18.23996, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 
    18.23994, 18.23994, 18.23995, 18.23994, 18.23992, 18.23992, 18.23992, 
    18.23991, 18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 
    18.23995, 18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23991, 18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 
    18.23994, 18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 
    18.23992, 18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 
    18.23992, 18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 
    18.23993, 18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 
    18.2399, 18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 
    18.23991, 18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 
    18.2399, 18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 
    18.23994, 18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 
    18.23986, 18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976202e-05, 5.976187e-05, 5.97619e-05, 5.976178e-05, 5.976185e-05, 
    5.976177e-05, 5.976199e-05, 5.976186e-05, 5.976194e-05, 5.9762e-05, 
    5.976155e-05, 5.976178e-05, 5.976132e-05, 5.976146e-05, 5.976111e-05, 
    5.976134e-05, 5.976106e-05, 5.976111e-05, 5.976095e-05, 5.9761e-05, 
    5.976079e-05, 5.976093e-05, 5.976068e-05, 5.976082e-05, 5.97608e-05, 
    5.976094e-05, 5.976173e-05, 5.976158e-05, 5.976174e-05, 5.976172e-05, 
    5.976173e-05, 5.976185e-05, 5.97619e-05, 5.976203e-05, 5.976201e-05, 
    5.976191e-05, 5.976171e-05, 5.976178e-05, 5.97616e-05, 5.976161e-05, 
    5.976141e-05, 5.97615e-05, 5.976117e-05, 5.976126e-05, 5.9761e-05, 
    5.976106e-05, 5.9761e-05, 5.976102e-05, 5.9761e-05, 5.97611e-05, 
    5.976106e-05, 5.976114e-05, 5.976148e-05, 5.976138e-05, 5.976168e-05, 
    5.976186e-05, 5.976198e-05, 5.976206e-05, 5.976205e-05, 5.976203e-05, 
    5.976191e-05, 5.97618e-05, 5.976172e-05, 5.976166e-05, 5.976161e-05, 
    5.976144e-05, 5.976135e-05, 5.976115e-05, 5.976119e-05, 5.976113e-05, 
    5.976107e-05, 5.976097e-05, 5.976099e-05, 5.976095e-05, 5.976113e-05, 
    5.976101e-05, 5.976121e-05, 5.976115e-05, 5.976159e-05, 5.976176e-05, 
    5.976183e-05, 5.976189e-05, 5.976205e-05, 5.976194e-05, 5.976198e-05, 
    5.976188e-05, 5.976182e-05, 5.976185e-05, 5.976166e-05, 5.976174e-05, 
    5.976135e-05, 5.976151e-05, 5.976108e-05, 5.976118e-05, 5.976105e-05, 
    5.976112e-05, 5.976101e-05, 5.976111e-05, 5.976093e-05, 5.976089e-05, 
    5.976092e-05, 5.976082e-05, 5.976111e-05, 5.9761e-05, 5.976185e-05, 
    5.976185e-05, 5.976182e-05, 5.976193e-05, 5.976193e-05, 5.976203e-05, 
    5.976194e-05, 5.976191e-05, 5.976182e-05, 5.976176e-05, 5.976171e-05, 
    5.97616e-05, 5.976147e-05, 5.97613e-05, 5.976118e-05, 5.976109e-05, 
    5.976114e-05, 5.97611e-05, 5.976115e-05, 5.976117e-05, 5.976091e-05, 
    5.976106e-05, 5.976083e-05, 5.976085e-05, 5.976095e-05, 5.976085e-05, 
    5.976184e-05, 5.976187e-05, 5.976197e-05, 5.976189e-05, 5.976204e-05, 
    5.976196e-05, 5.976191e-05, 5.976173e-05, 5.976169e-05, 5.976166e-05, 
    5.976159e-05, 5.97615e-05, 5.976133e-05, 5.976119e-05, 5.976107e-05, 
    5.976108e-05, 5.976107e-05, 5.976105e-05, 5.976111e-05, 5.976103e-05, 
    5.976102e-05, 5.976106e-05, 5.976085e-05, 5.976091e-05, 5.976085e-05, 
    5.976089e-05, 5.976186e-05, 5.976181e-05, 5.976184e-05, 5.976179e-05, 
    5.976183e-05, 5.976167e-05, 5.976162e-05, 5.976141e-05, 5.97615e-05, 
    5.976135e-05, 5.976148e-05, 5.976146e-05, 5.976135e-05, 5.976147e-05, 
    5.97612e-05, 5.976139e-05, 5.976105e-05, 5.976123e-05, 5.976103e-05, 
    5.976107e-05, 5.976101e-05, 5.976096e-05, 5.976089e-05, 5.976077e-05, 
    5.97608e-05, 5.976069e-05, 5.976174e-05, 5.976168e-05, 5.976169e-05, 
    5.976162e-05, 5.976157e-05, 5.976146e-05, 5.976129e-05, 5.976136e-05, 
    5.976124e-05, 5.976122e-05, 5.976139e-05, 5.976129e-05, 5.976163e-05, 
    5.976158e-05, 5.976161e-05, 5.976174e-05, 5.976134e-05, 5.976154e-05, 
    5.976117e-05, 5.976128e-05, 5.976097e-05, 5.976112e-05, 5.976081e-05, 
    5.976068e-05, 5.976055e-05, 5.976041e-05, 5.976165e-05, 5.976169e-05, 
    5.976161e-05, 5.97615e-05, 5.976141e-05, 5.976127e-05, 5.976126e-05, 
    5.976124e-05, 5.976117e-05, 5.976112e-05, 5.976123e-05, 5.976111e-05, 
    5.976157e-05, 5.976133e-05, 5.97617e-05, 5.976159e-05, 5.976151e-05, 
    5.976154e-05, 5.976137e-05, 5.976132e-05, 5.976115e-05, 5.976124e-05, 
    5.976071e-05, 5.976095e-05, 5.97603e-05, 5.976048e-05, 5.97617e-05, 
    5.976165e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 5.97612e-05, 
    5.976114e-05, 5.976107e-05, 5.976107e-05, 5.976103e-05, 5.97611e-05, 
    5.976103e-05, 5.976127e-05, 5.976117e-05, 5.976147e-05, 5.976139e-05, 
    5.976143e-05, 5.976146e-05, 5.976135e-05, 5.976123e-05, 5.976123e-05, 
    5.976119e-05, 5.976108e-05, 5.976127e-05, 5.976068e-05, 5.976104e-05, 
    5.976158e-05, 5.976147e-05, 5.976146e-05, 5.97615e-05, 5.976121e-05, 
    5.976131e-05, 5.976103e-05, 5.97611e-05, 5.976098e-05, 5.976104e-05, 
    5.976105e-05, 5.976113e-05, 5.976118e-05, 5.976131e-05, 5.976141e-05, 
    5.976149e-05, 5.976147e-05, 5.976138e-05, 5.976122e-05, 5.976107e-05, 
    5.97611e-05, 5.976099e-05, 5.976129e-05, 5.976116e-05, 5.976121e-05, 
    5.976109e-05, 5.976136e-05, 5.976113e-05, 5.976142e-05, 5.976139e-05, 
    5.976131e-05, 5.976115e-05, 5.976112e-05, 5.976108e-05, 5.97611e-05, 
    5.976122e-05, 5.976123e-05, 5.976131e-05, 5.976134e-05, 5.97614e-05, 
    5.976145e-05, 5.976141e-05, 5.976135e-05, 5.976122e-05, 5.976109e-05, 
    5.976095e-05, 5.976092e-05, 5.976076e-05, 5.976089e-05, 5.976068e-05, 
    5.976086e-05, 5.976055e-05, 5.976111e-05, 5.976087e-05, 5.976131e-05, 
    5.976126e-05, 5.976118e-05, 5.976098e-05, 5.976109e-05, 5.976096e-05, 
    5.976123e-05, 5.976138e-05, 5.976142e-05, 5.976149e-05, 5.976142e-05, 
    5.976142e-05, 5.976135e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976105e-05, 5.976096e-05, 5.97607e-05, 5.976055e-05, 5.976039e-05, 
    5.976032e-05, 5.97603e-05, 5.976029e-05 ;

 TOTLITC_1m =
  5.976202e-05, 5.976187e-05, 5.97619e-05, 5.976178e-05, 5.976185e-05, 
    5.976177e-05, 5.976199e-05, 5.976186e-05, 5.976194e-05, 5.9762e-05, 
    5.976155e-05, 5.976178e-05, 5.976132e-05, 5.976146e-05, 5.976111e-05, 
    5.976134e-05, 5.976106e-05, 5.976111e-05, 5.976095e-05, 5.9761e-05, 
    5.976079e-05, 5.976093e-05, 5.976068e-05, 5.976082e-05, 5.97608e-05, 
    5.976094e-05, 5.976173e-05, 5.976158e-05, 5.976174e-05, 5.976172e-05, 
    5.976173e-05, 5.976185e-05, 5.97619e-05, 5.976203e-05, 5.976201e-05, 
    5.976191e-05, 5.976171e-05, 5.976178e-05, 5.97616e-05, 5.976161e-05, 
    5.976141e-05, 5.97615e-05, 5.976117e-05, 5.976126e-05, 5.9761e-05, 
    5.976106e-05, 5.9761e-05, 5.976102e-05, 5.9761e-05, 5.97611e-05, 
    5.976106e-05, 5.976114e-05, 5.976148e-05, 5.976138e-05, 5.976168e-05, 
    5.976186e-05, 5.976198e-05, 5.976206e-05, 5.976205e-05, 5.976203e-05, 
    5.976191e-05, 5.97618e-05, 5.976172e-05, 5.976166e-05, 5.976161e-05, 
    5.976144e-05, 5.976135e-05, 5.976115e-05, 5.976119e-05, 5.976113e-05, 
    5.976107e-05, 5.976097e-05, 5.976099e-05, 5.976095e-05, 5.976113e-05, 
    5.976101e-05, 5.976121e-05, 5.976115e-05, 5.976159e-05, 5.976176e-05, 
    5.976183e-05, 5.976189e-05, 5.976205e-05, 5.976194e-05, 5.976198e-05, 
    5.976188e-05, 5.976182e-05, 5.976185e-05, 5.976166e-05, 5.976174e-05, 
    5.976135e-05, 5.976151e-05, 5.976108e-05, 5.976118e-05, 5.976105e-05, 
    5.976112e-05, 5.976101e-05, 5.976111e-05, 5.976093e-05, 5.976089e-05, 
    5.976092e-05, 5.976082e-05, 5.976111e-05, 5.9761e-05, 5.976185e-05, 
    5.976185e-05, 5.976182e-05, 5.976193e-05, 5.976193e-05, 5.976203e-05, 
    5.976194e-05, 5.976191e-05, 5.976182e-05, 5.976176e-05, 5.976171e-05, 
    5.97616e-05, 5.976147e-05, 5.97613e-05, 5.976118e-05, 5.976109e-05, 
    5.976114e-05, 5.97611e-05, 5.976115e-05, 5.976117e-05, 5.976091e-05, 
    5.976106e-05, 5.976083e-05, 5.976085e-05, 5.976095e-05, 5.976085e-05, 
    5.976184e-05, 5.976187e-05, 5.976197e-05, 5.976189e-05, 5.976204e-05, 
    5.976196e-05, 5.976191e-05, 5.976173e-05, 5.976169e-05, 5.976166e-05, 
    5.976159e-05, 5.97615e-05, 5.976133e-05, 5.976119e-05, 5.976107e-05, 
    5.976108e-05, 5.976107e-05, 5.976105e-05, 5.976111e-05, 5.976103e-05, 
    5.976102e-05, 5.976106e-05, 5.976085e-05, 5.976091e-05, 5.976085e-05, 
    5.976089e-05, 5.976186e-05, 5.976181e-05, 5.976184e-05, 5.976179e-05, 
    5.976183e-05, 5.976167e-05, 5.976162e-05, 5.976141e-05, 5.97615e-05, 
    5.976135e-05, 5.976148e-05, 5.976146e-05, 5.976135e-05, 5.976147e-05, 
    5.97612e-05, 5.976139e-05, 5.976105e-05, 5.976123e-05, 5.976103e-05, 
    5.976107e-05, 5.976101e-05, 5.976096e-05, 5.976089e-05, 5.976077e-05, 
    5.97608e-05, 5.976069e-05, 5.976174e-05, 5.976168e-05, 5.976169e-05, 
    5.976162e-05, 5.976157e-05, 5.976146e-05, 5.976129e-05, 5.976136e-05, 
    5.976124e-05, 5.976122e-05, 5.976139e-05, 5.976129e-05, 5.976163e-05, 
    5.976158e-05, 5.976161e-05, 5.976174e-05, 5.976134e-05, 5.976154e-05, 
    5.976117e-05, 5.976128e-05, 5.976097e-05, 5.976112e-05, 5.976081e-05, 
    5.976068e-05, 5.976055e-05, 5.976041e-05, 5.976165e-05, 5.976169e-05, 
    5.976161e-05, 5.97615e-05, 5.976141e-05, 5.976127e-05, 5.976126e-05, 
    5.976124e-05, 5.976117e-05, 5.976112e-05, 5.976123e-05, 5.976111e-05, 
    5.976157e-05, 5.976133e-05, 5.97617e-05, 5.976159e-05, 5.976151e-05, 
    5.976154e-05, 5.976137e-05, 5.976132e-05, 5.976115e-05, 5.976124e-05, 
    5.976071e-05, 5.976095e-05, 5.97603e-05, 5.976048e-05, 5.97617e-05, 
    5.976165e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 5.97612e-05, 
    5.976114e-05, 5.976107e-05, 5.976107e-05, 5.976103e-05, 5.97611e-05, 
    5.976103e-05, 5.976127e-05, 5.976117e-05, 5.976147e-05, 5.976139e-05, 
    5.976143e-05, 5.976146e-05, 5.976135e-05, 5.976123e-05, 5.976123e-05, 
    5.976119e-05, 5.976108e-05, 5.976127e-05, 5.976068e-05, 5.976104e-05, 
    5.976158e-05, 5.976147e-05, 5.976146e-05, 5.97615e-05, 5.976121e-05, 
    5.976131e-05, 5.976103e-05, 5.97611e-05, 5.976098e-05, 5.976104e-05, 
    5.976105e-05, 5.976113e-05, 5.976118e-05, 5.976131e-05, 5.976141e-05, 
    5.976149e-05, 5.976147e-05, 5.976138e-05, 5.976122e-05, 5.976107e-05, 
    5.97611e-05, 5.976099e-05, 5.976129e-05, 5.976116e-05, 5.976121e-05, 
    5.976109e-05, 5.976136e-05, 5.976113e-05, 5.976142e-05, 5.976139e-05, 
    5.976131e-05, 5.976115e-05, 5.976112e-05, 5.976108e-05, 5.97611e-05, 
    5.976122e-05, 5.976123e-05, 5.976131e-05, 5.976134e-05, 5.97614e-05, 
    5.976145e-05, 5.976141e-05, 5.976135e-05, 5.976122e-05, 5.976109e-05, 
    5.976095e-05, 5.976092e-05, 5.976076e-05, 5.976089e-05, 5.976068e-05, 
    5.976086e-05, 5.976055e-05, 5.976111e-05, 5.976087e-05, 5.976131e-05, 
    5.976126e-05, 5.976118e-05, 5.976098e-05, 5.976109e-05, 5.976096e-05, 
    5.976123e-05, 5.976138e-05, 5.976142e-05, 5.976149e-05, 5.976142e-05, 
    5.976142e-05, 5.976135e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976105e-05, 5.976096e-05, 5.97607e-05, 5.976055e-05, 5.976039e-05, 
    5.976032e-05, 5.97603e-05, 5.976029e-05 ;

 TOTLITN =
  1.375929e-06, 1.375925e-06, 1.375925e-06, 1.375922e-06, 1.375924e-06, 
    1.375922e-06, 1.375928e-06, 1.375924e-06, 1.375927e-06, 1.375928e-06, 
    1.375916e-06, 1.375922e-06, 1.375909e-06, 1.375913e-06, 1.375903e-06, 
    1.37591e-06, 1.375902e-06, 1.375903e-06, 1.375899e-06, 1.3759e-06, 
    1.375894e-06, 1.375898e-06, 1.375891e-06, 1.375895e-06, 1.375894e-06, 
    1.375898e-06, 1.375921e-06, 1.375916e-06, 1.375921e-06, 1.37592e-06, 
    1.375921e-06, 1.375924e-06, 1.375925e-06, 1.375929e-06, 1.375928e-06, 
    1.375926e-06, 1.37592e-06, 1.375922e-06, 1.375917e-06, 1.375917e-06, 
    1.375912e-06, 1.375914e-06, 1.375905e-06, 1.375907e-06, 1.3759e-06, 
    1.375902e-06, 1.3759e-06, 1.375901e-06, 1.3759e-06, 1.375903e-06, 
    1.375902e-06, 1.375904e-06, 1.375914e-06, 1.375911e-06, 1.375919e-06, 
    1.375924e-06, 1.375928e-06, 1.37593e-06, 1.37593e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.37592e-06, 1.375919e-06, 1.375917e-06, 
    1.375912e-06, 1.37591e-06, 1.375904e-06, 1.375905e-06, 1.375904e-06, 
    1.375902e-06, 1.375899e-06, 1.3759e-06, 1.375899e-06, 1.375904e-06, 
    1.3759e-06, 1.375906e-06, 1.375904e-06, 1.375917e-06, 1.375921e-06, 
    1.375923e-06, 1.375925e-06, 1.375929e-06, 1.375926e-06, 1.375928e-06, 
    1.375925e-06, 1.375923e-06, 1.375924e-06, 1.375919e-06, 1.375921e-06, 
    1.37591e-06, 1.375915e-06, 1.375902e-06, 1.375905e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375903e-06, 1.375898e-06, 1.375897e-06, 
    1.375898e-06, 1.375895e-06, 1.375903e-06, 1.3759e-06, 1.375924e-06, 
    1.375924e-06, 1.375923e-06, 1.375926e-06, 1.375926e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375923e-06, 1.375921e-06, 1.37592e-06, 
    1.375917e-06, 1.375913e-06, 1.375908e-06, 1.375905e-06, 1.375903e-06, 
    1.375904e-06, 1.375903e-06, 1.375904e-06, 1.375905e-06, 1.375897e-06, 
    1.375902e-06, 1.375895e-06, 1.375896e-06, 1.375898e-06, 1.375896e-06, 
    1.375924e-06, 1.375925e-06, 1.375927e-06, 1.375925e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375921e-06, 1.37592e-06, 1.375918e-06, 
    1.375917e-06, 1.375914e-06, 1.375909e-06, 1.375906e-06, 1.375902e-06, 
    1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 1.375901e-06, 
    1.375901e-06, 1.375902e-06, 1.375896e-06, 1.375897e-06, 1.375896e-06, 
    1.375897e-06, 1.375924e-06, 1.375923e-06, 1.375924e-06, 1.375922e-06, 
    1.375923e-06, 1.375919e-06, 1.375918e-06, 1.375912e-06, 1.375914e-06, 
    1.37591e-06, 1.375914e-06, 1.375913e-06, 1.37591e-06, 1.375913e-06, 
    1.375906e-06, 1.375911e-06, 1.375901e-06, 1.375906e-06, 1.375901e-06, 
    1.375902e-06, 1.3759e-06, 1.375899e-06, 1.375897e-06, 1.375893e-06, 
    1.375894e-06, 1.375891e-06, 1.375921e-06, 1.375919e-06, 1.375919e-06, 
    1.375917e-06, 1.375916e-06, 1.375913e-06, 1.375908e-06, 1.37591e-06, 
    1.375907e-06, 1.375906e-06, 1.375911e-06, 1.375908e-06, 1.375918e-06, 
    1.375916e-06, 1.375917e-06, 1.375921e-06, 1.37591e-06, 1.375915e-06, 
    1.375905e-06, 1.375908e-06, 1.375899e-06, 1.375903e-06, 1.375895e-06, 
    1.375891e-06, 1.375887e-06, 1.375883e-06, 1.375918e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375911e-06, 1.375908e-06, 1.375907e-06, 
    1.375907e-06, 1.375905e-06, 1.375903e-06, 1.375906e-06, 1.375903e-06, 
    1.375916e-06, 1.375909e-06, 1.37592e-06, 1.375917e-06, 1.375914e-06, 
    1.375915e-06, 1.37591e-06, 1.375909e-06, 1.375904e-06, 1.375907e-06, 
    1.375892e-06, 1.375898e-06, 1.37588e-06, 1.375885e-06, 1.37592e-06, 
    1.375918e-06, 1.375912e-06, 1.375915e-06, 1.375908e-06, 1.375906e-06, 
    1.375904e-06, 1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 
    1.375901e-06, 1.375908e-06, 1.375905e-06, 1.375913e-06, 1.375911e-06, 
    1.375912e-06, 1.375913e-06, 1.37591e-06, 1.375906e-06, 1.375906e-06, 
    1.375905e-06, 1.375902e-06, 1.375907e-06, 1.375891e-06, 1.375901e-06, 
    1.375916e-06, 1.375913e-06, 1.375913e-06, 1.375914e-06, 1.375906e-06, 
    1.375909e-06, 1.375901e-06, 1.375903e-06, 1.375899e-06, 1.375901e-06, 
    1.375901e-06, 1.375904e-06, 1.375905e-06, 1.375909e-06, 1.375912e-06, 
    1.375914e-06, 1.375913e-06, 1.375911e-06, 1.375906e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375908e-06, 1.375905e-06, 1.375906e-06, 
    1.375902e-06, 1.37591e-06, 1.375903e-06, 1.375912e-06, 1.375911e-06, 
    1.375909e-06, 1.375904e-06, 1.375903e-06, 1.375902e-06, 1.375903e-06, 
    1.375906e-06, 1.375907e-06, 1.375909e-06, 1.37591e-06, 1.375911e-06, 
    1.375913e-06, 1.375911e-06, 1.37591e-06, 1.375906e-06, 1.375903e-06, 
    1.375899e-06, 1.375898e-06, 1.375893e-06, 1.375897e-06, 1.375891e-06, 
    1.375896e-06, 1.375887e-06, 1.375903e-06, 1.375896e-06, 1.375909e-06, 
    1.375907e-06, 1.375905e-06, 1.375899e-06, 1.375902e-06, 1.375899e-06, 
    1.375907e-06, 1.375911e-06, 1.375912e-06, 1.375914e-06, 1.375912e-06, 
    1.375912e-06, 1.37591e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375901e-06, 1.375899e-06, 1.375892e-06, 1.375887e-06, 1.375883e-06, 
    1.375881e-06, 1.37588e-06, 1.37588e-06 ;

 TOTLITN_1m =
  1.375929e-06, 1.375925e-06, 1.375925e-06, 1.375922e-06, 1.375924e-06, 
    1.375922e-06, 1.375928e-06, 1.375924e-06, 1.375927e-06, 1.375928e-06, 
    1.375916e-06, 1.375922e-06, 1.375909e-06, 1.375913e-06, 1.375903e-06, 
    1.37591e-06, 1.375902e-06, 1.375903e-06, 1.375899e-06, 1.3759e-06, 
    1.375894e-06, 1.375898e-06, 1.375891e-06, 1.375895e-06, 1.375894e-06, 
    1.375898e-06, 1.375921e-06, 1.375916e-06, 1.375921e-06, 1.37592e-06, 
    1.375921e-06, 1.375924e-06, 1.375925e-06, 1.375929e-06, 1.375928e-06, 
    1.375926e-06, 1.37592e-06, 1.375922e-06, 1.375917e-06, 1.375917e-06, 
    1.375912e-06, 1.375914e-06, 1.375905e-06, 1.375907e-06, 1.3759e-06, 
    1.375902e-06, 1.3759e-06, 1.375901e-06, 1.3759e-06, 1.375903e-06, 
    1.375902e-06, 1.375904e-06, 1.375914e-06, 1.375911e-06, 1.375919e-06, 
    1.375924e-06, 1.375928e-06, 1.37593e-06, 1.37593e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.37592e-06, 1.375919e-06, 1.375917e-06, 
    1.375912e-06, 1.37591e-06, 1.375904e-06, 1.375905e-06, 1.375904e-06, 
    1.375902e-06, 1.375899e-06, 1.3759e-06, 1.375899e-06, 1.375904e-06, 
    1.3759e-06, 1.375906e-06, 1.375904e-06, 1.375917e-06, 1.375921e-06, 
    1.375923e-06, 1.375925e-06, 1.375929e-06, 1.375926e-06, 1.375928e-06, 
    1.375925e-06, 1.375923e-06, 1.375924e-06, 1.375919e-06, 1.375921e-06, 
    1.37591e-06, 1.375915e-06, 1.375902e-06, 1.375905e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375903e-06, 1.375898e-06, 1.375897e-06, 
    1.375898e-06, 1.375895e-06, 1.375903e-06, 1.3759e-06, 1.375924e-06, 
    1.375924e-06, 1.375923e-06, 1.375926e-06, 1.375926e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375923e-06, 1.375921e-06, 1.37592e-06, 
    1.375917e-06, 1.375913e-06, 1.375908e-06, 1.375905e-06, 1.375903e-06, 
    1.375904e-06, 1.375903e-06, 1.375904e-06, 1.375905e-06, 1.375897e-06, 
    1.375902e-06, 1.375895e-06, 1.375896e-06, 1.375898e-06, 1.375896e-06, 
    1.375924e-06, 1.375925e-06, 1.375927e-06, 1.375925e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375921e-06, 1.37592e-06, 1.375918e-06, 
    1.375917e-06, 1.375914e-06, 1.375909e-06, 1.375906e-06, 1.375902e-06, 
    1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 1.375901e-06, 
    1.375901e-06, 1.375902e-06, 1.375896e-06, 1.375897e-06, 1.375896e-06, 
    1.375897e-06, 1.375924e-06, 1.375923e-06, 1.375924e-06, 1.375922e-06, 
    1.375923e-06, 1.375919e-06, 1.375918e-06, 1.375912e-06, 1.375914e-06, 
    1.37591e-06, 1.375914e-06, 1.375913e-06, 1.37591e-06, 1.375913e-06, 
    1.375906e-06, 1.375911e-06, 1.375901e-06, 1.375906e-06, 1.375901e-06, 
    1.375902e-06, 1.3759e-06, 1.375899e-06, 1.375897e-06, 1.375893e-06, 
    1.375894e-06, 1.375891e-06, 1.375921e-06, 1.375919e-06, 1.375919e-06, 
    1.375917e-06, 1.375916e-06, 1.375913e-06, 1.375908e-06, 1.37591e-06, 
    1.375907e-06, 1.375906e-06, 1.375911e-06, 1.375908e-06, 1.375918e-06, 
    1.375916e-06, 1.375917e-06, 1.375921e-06, 1.37591e-06, 1.375915e-06, 
    1.375905e-06, 1.375908e-06, 1.375899e-06, 1.375903e-06, 1.375895e-06, 
    1.375891e-06, 1.375887e-06, 1.375883e-06, 1.375918e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375911e-06, 1.375908e-06, 1.375907e-06, 
    1.375907e-06, 1.375905e-06, 1.375903e-06, 1.375906e-06, 1.375903e-06, 
    1.375916e-06, 1.375909e-06, 1.37592e-06, 1.375917e-06, 1.375914e-06, 
    1.375915e-06, 1.37591e-06, 1.375909e-06, 1.375904e-06, 1.375907e-06, 
    1.375892e-06, 1.375898e-06, 1.37588e-06, 1.375885e-06, 1.37592e-06, 
    1.375918e-06, 1.375912e-06, 1.375915e-06, 1.375908e-06, 1.375906e-06, 
    1.375904e-06, 1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 
    1.375901e-06, 1.375908e-06, 1.375905e-06, 1.375913e-06, 1.375911e-06, 
    1.375912e-06, 1.375913e-06, 1.37591e-06, 1.375906e-06, 1.375906e-06, 
    1.375905e-06, 1.375902e-06, 1.375907e-06, 1.375891e-06, 1.375901e-06, 
    1.375916e-06, 1.375913e-06, 1.375913e-06, 1.375914e-06, 1.375906e-06, 
    1.375909e-06, 1.375901e-06, 1.375903e-06, 1.375899e-06, 1.375901e-06, 
    1.375901e-06, 1.375904e-06, 1.375905e-06, 1.375909e-06, 1.375912e-06, 
    1.375914e-06, 1.375913e-06, 1.375911e-06, 1.375906e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375908e-06, 1.375905e-06, 1.375906e-06, 
    1.375902e-06, 1.37591e-06, 1.375903e-06, 1.375912e-06, 1.375911e-06, 
    1.375909e-06, 1.375904e-06, 1.375903e-06, 1.375902e-06, 1.375903e-06, 
    1.375906e-06, 1.375907e-06, 1.375909e-06, 1.37591e-06, 1.375911e-06, 
    1.375913e-06, 1.375911e-06, 1.37591e-06, 1.375906e-06, 1.375903e-06, 
    1.375899e-06, 1.375898e-06, 1.375893e-06, 1.375897e-06, 1.375891e-06, 
    1.375896e-06, 1.375887e-06, 1.375903e-06, 1.375896e-06, 1.375909e-06, 
    1.375907e-06, 1.375905e-06, 1.375899e-06, 1.375902e-06, 1.375899e-06, 
    1.375907e-06, 1.375911e-06, 1.375912e-06, 1.375914e-06, 1.375912e-06, 
    1.375912e-06, 1.37591e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375901e-06, 1.375899e-06, 1.375892e-06, 1.375887e-06, 1.375883e-06, 
    1.375881e-06, 1.37588e-06, 1.37588e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMC_1m =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMN =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773752, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773751, 1.773751, 1.77375, 1.773748, 1.773747, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTSOMN_1m =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773752, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773751, 1.773751, 1.77375, 1.773748, 1.773747, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  243.0876, 243.0908, 243.0902, 243.0928, 243.0914, 243.093, 243.0883, 
    243.0909, 243.0892, 243.0879, 243.0977, 243.0929, 243.1028, 243.0998, 
    243.1075, 243.1023, 243.1086, 243.1074, 243.111, 243.11, 243.1144, 
    243.1115, 243.1168, 243.1138, 243.1142, 243.1114, 243.0939, 243.0971, 
    243.0937, 243.0942, 243.094, 243.0914, 243.09, 243.0874, 243.0879, 
    243.0898, 243.0944, 243.0929, 243.0968, 243.0967, 243.1009, 243.099, 
    243.1062, 243.1042, 243.11, 243.1085, 243.1099, 243.1095, 243.11, 
    243.1078, 243.1087, 243.1068, 243.0994, 243.1015, 243.095, 243.0909, 
    243.0884, 243.0865, 243.0868, 243.0873, 243.0899, 243.0923, 243.0942, 
    243.0954, 243.0966, 243.1002, 243.1022, 243.1066, 243.1058, 243.1071, 
    243.1084, 243.1105, 243.1102, 243.1111, 243.1071, 243.1097, 243.1054, 
    243.1066, 243.0968, 243.0933, 243.0916, 243.0903, 243.087, 243.0893, 
    243.0884, 243.0906, 243.0919, 243.0913, 243.0955, 243.0938, 243.1023, 
    243.0987, 243.1082, 243.106, 243.1088, 243.1074, 243.1098, 243.1076, 
    243.1114, 243.1122, 243.1117, 243.1139, 243.1075, 243.1099, 243.0912, 
    243.0914, 243.0919, 243.0896, 243.0894, 243.0874, 243.0892, 243.09, 
    243.092, 243.0932, 243.0943, 243.0968, 243.0995, 243.1033, 243.1061, 
    243.108, 243.1068, 243.1078, 243.1067, 243.1062, 243.1119, 243.1087, 
    243.1136, 243.1133, 243.1111, 243.1133, 243.0914, 243.0908, 243.0885, 
    243.0903, 243.0871, 243.0889, 243.0899, 243.0938, 243.0947, 243.0955, 
    243.0971, 243.0991, 243.1026, 243.1057, 243.1085, 243.1083, 243.1084, 
    243.109, 243.1074, 243.1092, 243.1095, 243.1087, 243.1133, 243.112, 
    243.1133, 243.1125, 243.091, 243.0921, 243.0915, 243.0926, 243.0918, 
    243.0952, 243.0962, 243.101, 243.0991, 243.1021, 243.0994, 243.0999, 
    243.1022, 243.0995, 243.1055, 243.1014, 243.109, 243.1049, 243.1092, 
    243.1085, 243.1098, 243.1109, 243.1123, 243.115, 243.1144, 243.1166, 
    243.0937, 243.095, 243.095, 243.0964, 243.0975, 243.0998, 243.1035, 
    243.1021, 243.1047, 243.1052, 243.1013, 243.1037, 243.096, 243.0972, 
    243.0965, 243.0938, 243.1024, 243.098, 243.1062, 243.1038, 243.1107, 
    243.1072, 243.114, 243.1168, 243.1196, 243.1227, 243.0958, 243.0949, 
    243.0966, 243.0989, 243.1011, 243.1039, 243.1042, 243.1048, 243.1062, 
    243.1073, 243.1049, 243.1076, 243.0974, 243.1028, 243.0945, 243.097, 
    243.0987, 243.098, 243.102, 243.1029, 243.1066, 243.1047, 243.1161, 
    243.1111, 243.1251, 243.1212, 243.0946, 243.0958, 243.1002, 243.0981, 
    243.1041, 243.1056, 243.1068, 243.1083, 243.1085, 243.1093, 243.1079, 
    243.1093, 243.1039, 243.1063, 243.0997, 243.1013, 243.1006, 243.0998, 
    243.1023, 243.1049, 243.105, 243.1059, 243.1081, 243.1042, 243.1166, 
    243.1089, 243.0972, 243.0996, 243.1, 243.0991, 243.1054, 243.1031, 
    243.1093, 243.1077, 243.1104, 243.109, 243.1088, 243.1071, 243.106, 
    243.1032, 243.101, 243.0992, 243.0996, 243.1015, 243.1051, 243.1085, 
    243.1077, 243.1102, 243.1037, 243.1064, 243.1053, 243.1081, 243.1021, 
    243.1071, 243.1008, 243.1013, 243.1031, 243.1065, 243.1074, 243.1082, 
    243.1077, 243.1052, 243.1048, 243.103, 243.1025, 243.1012, 243.1001, 
    243.1011, 243.1022, 243.1052, 243.1079, 243.1109, 243.1116, 243.1149, 
    243.1122, 243.1167, 243.1127, 243.1196, 243.1074, 243.1127, 243.1032, 
    243.1042, 243.1061, 243.1104, 243.1081, 243.1108, 243.1048, 243.1016, 
    243.1008, 243.0993, 243.1009, 243.1007, 243.1022, 243.1018, 243.1053, 
    243.1034, 243.1088, 243.1108, 243.1163, 243.1197, 243.1232, 243.1247, 
    243.1251, 243.1253 ;

 TREFMNAV_R =
  243.0876, 243.0908, 243.0902, 243.0928, 243.0914, 243.093, 243.0883, 
    243.0909, 243.0892, 243.0879, 243.0977, 243.0929, 243.1028, 243.0998, 
    243.1075, 243.1023, 243.1086, 243.1074, 243.111, 243.11, 243.1144, 
    243.1115, 243.1168, 243.1138, 243.1142, 243.1114, 243.0939, 243.0971, 
    243.0937, 243.0942, 243.094, 243.0914, 243.09, 243.0874, 243.0879, 
    243.0898, 243.0944, 243.0929, 243.0968, 243.0967, 243.1009, 243.099, 
    243.1062, 243.1042, 243.11, 243.1085, 243.1099, 243.1095, 243.11, 
    243.1078, 243.1087, 243.1068, 243.0994, 243.1015, 243.095, 243.0909, 
    243.0884, 243.0865, 243.0868, 243.0873, 243.0899, 243.0923, 243.0942, 
    243.0954, 243.0966, 243.1002, 243.1022, 243.1066, 243.1058, 243.1071, 
    243.1084, 243.1105, 243.1102, 243.1111, 243.1071, 243.1097, 243.1054, 
    243.1066, 243.0968, 243.0933, 243.0916, 243.0903, 243.087, 243.0893, 
    243.0884, 243.0906, 243.0919, 243.0913, 243.0955, 243.0938, 243.1023, 
    243.0987, 243.1082, 243.106, 243.1088, 243.1074, 243.1098, 243.1076, 
    243.1114, 243.1122, 243.1117, 243.1139, 243.1075, 243.1099, 243.0912, 
    243.0914, 243.0919, 243.0896, 243.0894, 243.0874, 243.0892, 243.09, 
    243.092, 243.0932, 243.0943, 243.0968, 243.0995, 243.1033, 243.1061, 
    243.108, 243.1068, 243.1078, 243.1067, 243.1062, 243.1119, 243.1087, 
    243.1136, 243.1133, 243.1111, 243.1133, 243.0914, 243.0908, 243.0885, 
    243.0903, 243.0871, 243.0889, 243.0899, 243.0938, 243.0947, 243.0955, 
    243.0971, 243.0991, 243.1026, 243.1057, 243.1085, 243.1083, 243.1084, 
    243.109, 243.1074, 243.1092, 243.1095, 243.1087, 243.1133, 243.112, 
    243.1133, 243.1125, 243.091, 243.0921, 243.0915, 243.0926, 243.0918, 
    243.0952, 243.0962, 243.101, 243.0991, 243.1021, 243.0994, 243.0999, 
    243.1022, 243.0995, 243.1055, 243.1014, 243.109, 243.1049, 243.1092, 
    243.1085, 243.1098, 243.1109, 243.1123, 243.115, 243.1144, 243.1166, 
    243.0937, 243.095, 243.095, 243.0964, 243.0975, 243.0998, 243.1035, 
    243.1021, 243.1047, 243.1052, 243.1013, 243.1037, 243.096, 243.0972, 
    243.0965, 243.0938, 243.1024, 243.098, 243.1062, 243.1038, 243.1107, 
    243.1072, 243.114, 243.1168, 243.1196, 243.1227, 243.0958, 243.0949, 
    243.0966, 243.0989, 243.1011, 243.1039, 243.1042, 243.1048, 243.1062, 
    243.1073, 243.1049, 243.1076, 243.0974, 243.1028, 243.0945, 243.097, 
    243.0987, 243.098, 243.102, 243.1029, 243.1066, 243.1047, 243.1161, 
    243.1111, 243.1251, 243.1212, 243.0946, 243.0958, 243.1002, 243.0981, 
    243.1041, 243.1056, 243.1068, 243.1083, 243.1085, 243.1093, 243.1079, 
    243.1093, 243.1039, 243.1063, 243.0997, 243.1013, 243.1006, 243.0998, 
    243.1023, 243.1049, 243.105, 243.1059, 243.1081, 243.1042, 243.1166, 
    243.1089, 243.0972, 243.0996, 243.1, 243.0991, 243.1054, 243.1031, 
    243.1093, 243.1077, 243.1104, 243.109, 243.1088, 243.1071, 243.106, 
    243.1032, 243.101, 243.0992, 243.0996, 243.1015, 243.1051, 243.1085, 
    243.1077, 243.1102, 243.1037, 243.1064, 243.1053, 243.1081, 243.1021, 
    243.1071, 243.1008, 243.1013, 243.1031, 243.1065, 243.1074, 243.1082, 
    243.1077, 243.1052, 243.1048, 243.103, 243.1025, 243.1012, 243.1001, 
    243.1011, 243.1022, 243.1052, 243.1079, 243.1109, 243.1116, 243.1149, 
    243.1122, 243.1167, 243.1127, 243.1196, 243.1074, 243.1127, 243.1032, 
    243.1042, 243.1061, 243.1104, 243.1081, 243.1108, 243.1048, 243.1016, 
    243.1008, 243.0993, 243.1009, 243.1007, 243.1022, 243.1018, 243.1053, 
    243.1034, 243.1088, 243.1108, 243.1163, 243.1197, 243.1232, 243.1247, 
    243.1251, 243.1253 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  270.7643, 270.7622, 270.7626, 270.7609, 270.7618, 270.7607, 270.7638, 
    270.7621, 270.7632, 270.7641, 270.7577, 270.7608, 270.7543, 270.7563, 
    270.7512, 270.7546, 270.7505, 270.7512, 270.7488, 270.7495, 270.7466, 
    270.7485, 270.745, 270.747, 270.7467, 270.7486, 270.7601, 270.7581, 
    270.7603, 270.76, 270.7601, 270.7618, 270.7627, 270.7644, 270.7641, 
    270.7628, 270.7598, 270.7608, 270.7583, 270.7583, 270.7555, 270.7568, 
    270.752, 270.7534, 270.7495, 270.7505, 270.7495, 270.7498, 270.7495, 
    270.751, 270.7504, 270.7516, 270.7566, 270.7551, 270.7594, 270.7621, 
    270.7638, 270.765, 270.7648, 270.7645, 270.7628, 270.7612, 270.7599, 
    270.7592, 270.7583, 270.756, 270.7547, 270.7518, 270.7523, 270.7514, 
    270.7506, 270.7492, 270.7494, 270.7488, 270.7514, 270.7497, 270.7526, 
    270.7518, 270.7583, 270.7606, 270.7617, 270.7625, 270.7647, 270.7632, 
    270.7638, 270.7623, 270.7614, 270.7619, 270.7591, 270.7602, 270.7546, 
    270.757, 270.7507, 270.7522, 270.7503, 270.7513, 270.7496, 270.7511, 
    270.7485, 270.748, 270.7484, 270.7469, 270.7512, 270.7495, 270.7619, 
    270.7618, 270.7615, 270.763, 270.7631, 270.7644, 270.7632, 270.7627, 
    270.7614, 270.7606, 270.7599, 270.7582, 270.7565, 270.7539, 270.7521, 
    270.7509, 270.7516, 270.7509, 270.7517, 270.752, 270.7482, 270.7504, 
    270.7471, 270.7473, 270.7488, 270.7473, 270.7618, 270.7622, 270.7636, 
    270.7625, 270.7646, 270.7634, 270.7628, 270.7602, 270.7596, 270.7591, 
    270.7581, 270.7567, 270.7544, 270.7524, 270.7505, 270.7506, 270.7506, 
    270.7502, 270.7512, 270.75, 270.7498, 270.7504, 270.7473, 270.7482, 
    270.7473, 270.7479, 270.7621, 270.7614, 270.7617, 270.761, 270.7615, 
    270.7593, 270.7586, 270.7555, 270.7568, 270.7547, 270.7565, 270.7562, 
    270.7547, 270.7564, 270.7525, 270.7552, 270.7502, 270.7529, 270.75, 
    270.7505, 270.7497, 270.7489, 270.748, 270.7462, 270.7466, 270.7451, 
    270.7603, 270.7594, 270.7595, 270.7585, 270.7578, 270.7563, 270.7538, 
    270.7547, 270.7531, 270.7527, 270.7553, 270.7537, 270.7588, 270.758, 
    270.7585, 270.7602, 270.7546, 270.7575, 270.7521, 270.7536, 270.749, 
    270.7513, 270.7468, 270.7449, 270.7431, 270.741, 270.7589, 270.7595, 
    270.7584, 270.7569, 270.7554, 270.7535, 270.7533, 270.753, 270.7521, 
    270.7513, 270.7529, 270.7511, 270.7579, 270.7543, 270.7597, 270.7581, 
    270.757, 270.7574, 270.7548, 270.7542, 270.7518, 270.753, 270.7454, 
    270.7488, 270.7394, 270.742, 270.7597, 270.7589, 270.756, 270.7574, 
    270.7534, 270.7524, 270.7516, 270.7506, 270.7505, 270.7499, 270.7509, 
    270.75, 270.7535, 270.752, 270.7563, 270.7552, 270.7557, 270.7563, 
    270.7546, 270.7529, 270.7528, 270.7523, 270.7508, 270.7534, 270.7451, 
    270.7503, 270.758, 270.7564, 270.7561, 270.7567, 270.7525, 270.7541, 
    270.7499, 270.7511, 270.7492, 270.7502, 270.7503, 270.7514, 270.7522, 
    270.754, 270.7555, 270.7567, 270.7564, 270.7551, 270.7528, 270.7505, 
    270.751, 270.7494, 270.7537, 270.7519, 270.7526, 270.7508, 270.7548, 
    270.7515, 270.7556, 270.7552, 270.7541, 270.7518, 270.7513, 270.7507, 
    270.751, 270.7527, 270.753, 270.7541, 270.7545, 270.7553, 270.7561, 
    270.7554, 270.7547, 270.7527, 270.7509, 270.7489, 270.7484, 270.7462, 
    270.748, 270.7451, 270.7477, 270.7431, 270.7512, 270.7477, 270.754, 
    270.7534, 270.7521, 270.7493, 270.7508, 270.749, 270.753, 270.7551, 
    270.7556, 270.7566, 270.7556, 270.7556, 270.7547, 270.755, 270.7526, 
    270.7539, 270.7503, 270.749, 270.7453, 270.743, 270.7407, 270.7397, 
    270.7393, 270.7392 ;

 TREFMXAV_R =
  270.7643, 270.7622, 270.7626, 270.7609, 270.7618, 270.7607, 270.7638, 
    270.7621, 270.7632, 270.7641, 270.7577, 270.7608, 270.7543, 270.7563, 
    270.7512, 270.7546, 270.7505, 270.7512, 270.7488, 270.7495, 270.7466, 
    270.7485, 270.745, 270.747, 270.7467, 270.7486, 270.7601, 270.7581, 
    270.7603, 270.76, 270.7601, 270.7618, 270.7627, 270.7644, 270.7641, 
    270.7628, 270.7598, 270.7608, 270.7583, 270.7583, 270.7555, 270.7568, 
    270.752, 270.7534, 270.7495, 270.7505, 270.7495, 270.7498, 270.7495, 
    270.751, 270.7504, 270.7516, 270.7566, 270.7551, 270.7594, 270.7621, 
    270.7638, 270.765, 270.7648, 270.7645, 270.7628, 270.7612, 270.7599, 
    270.7592, 270.7583, 270.756, 270.7547, 270.7518, 270.7523, 270.7514, 
    270.7506, 270.7492, 270.7494, 270.7488, 270.7514, 270.7497, 270.7526, 
    270.7518, 270.7583, 270.7606, 270.7617, 270.7625, 270.7647, 270.7632, 
    270.7638, 270.7623, 270.7614, 270.7619, 270.7591, 270.7602, 270.7546, 
    270.757, 270.7507, 270.7522, 270.7503, 270.7513, 270.7496, 270.7511, 
    270.7485, 270.748, 270.7484, 270.7469, 270.7512, 270.7495, 270.7619, 
    270.7618, 270.7615, 270.763, 270.7631, 270.7644, 270.7632, 270.7627, 
    270.7614, 270.7606, 270.7599, 270.7582, 270.7565, 270.7539, 270.7521, 
    270.7509, 270.7516, 270.7509, 270.7517, 270.752, 270.7482, 270.7504, 
    270.7471, 270.7473, 270.7488, 270.7473, 270.7618, 270.7622, 270.7636, 
    270.7625, 270.7646, 270.7634, 270.7628, 270.7602, 270.7596, 270.7591, 
    270.7581, 270.7567, 270.7544, 270.7524, 270.7505, 270.7506, 270.7506, 
    270.7502, 270.7512, 270.75, 270.7498, 270.7504, 270.7473, 270.7482, 
    270.7473, 270.7479, 270.7621, 270.7614, 270.7617, 270.761, 270.7615, 
    270.7593, 270.7586, 270.7555, 270.7568, 270.7547, 270.7565, 270.7562, 
    270.7547, 270.7564, 270.7525, 270.7552, 270.7502, 270.7529, 270.75, 
    270.7505, 270.7497, 270.7489, 270.748, 270.7462, 270.7466, 270.7451, 
    270.7603, 270.7594, 270.7595, 270.7585, 270.7578, 270.7563, 270.7538, 
    270.7547, 270.7531, 270.7527, 270.7553, 270.7537, 270.7588, 270.758, 
    270.7585, 270.7602, 270.7546, 270.7575, 270.7521, 270.7536, 270.749, 
    270.7513, 270.7468, 270.7449, 270.7431, 270.741, 270.7589, 270.7595, 
    270.7584, 270.7569, 270.7554, 270.7535, 270.7533, 270.753, 270.7521, 
    270.7513, 270.7529, 270.7511, 270.7579, 270.7543, 270.7597, 270.7581, 
    270.757, 270.7574, 270.7548, 270.7542, 270.7518, 270.753, 270.7454, 
    270.7488, 270.7394, 270.742, 270.7597, 270.7589, 270.756, 270.7574, 
    270.7534, 270.7524, 270.7516, 270.7506, 270.7505, 270.7499, 270.7509, 
    270.75, 270.7535, 270.752, 270.7563, 270.7552, 270.7557, 270.7563, 
    270.7546, 270.7529, 270.7528, 270.7523, 270.7508, 270.7534, 270.7451, 
    270.7503, 270.758, 270.7564, 270.7561, 270.7567, 270.7525, 270.7541, 
    270.7499, 270.7511, 270.7492, 270.7502, 270.7503, 270.7514, 270.7522, 
    270.754, 270.7555, 270.7567, 270.7564, 270.7551, 270.7528, 270.7505, 
    270.751, 270.7494, 270.7537, 270.7519, 270.7526, 270.7508, 270.7548, 
    270.7515, 270.7556, 270.7552, 270.7541, 270.7518, 270.7513, 270.7507, 
    270.751, 270.7527, 270.753, 270.7541, 270.7545, 270.7553, 270.7561, 
    270.7554, 270.7547, 270.7527, 270.7509, 270.7489, 270.7484, 270.7462, 
    270.748, 270.7451, 270.7477, 270.7431, 270.7512, 270.7477, 270.754, 
    270.7534, 270.7521, 270.7493, 270.7508, 270.749, 270.753, 270.7551, 
    270.7556, 270.7566, 270.7556, 270.7556, 270.7547, 270.755, 270.7526, 
    270.7539, 270.7503, 270.749, 270.7453, 270.743, 270.7407, 270.7397, 
    270.7393, 270.7392 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  255.2032, 255.203, 255.2031, 255.203, 255.203, 255.2029, 255.2032, 255.203, 
    255.2031, 255.2032, 255.2027, 255.2029, 255.2025, 255.2026, 255.2022, 
    255.2025, 255.2022, 255.2022, 255.2021, 255.2021, 255.2019, 255.202, 
    255.2018, 255.2019, 255.2019, 255.202, 255.2029, 255.2028, 255.2029, 
    255.2029, 255.2029, 255.203, 255.2031, 255.2032, 255.2032, 255.2031, 
    255.2029, 255.2029, 255.2028, 255.2028, 255.2026, 255.2027, 255.2023, 
    255.2024, 255.2021, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2022, 255.2023, 255.2026, 255.2025, 255.2029, 255.203, 255.2032, 
    255.2032, 255.2032, 255.2032, 255.2031, 255.203, 255.2029, 255.2028, 
    255.2028, 255.2026, 255.2025, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2021, 255.2021, 255.2021, 255.2023, 255.2021, 255.2023, 255.2023, 
    255.2028, 255.2029, 255.203, 255.2031, 255.2032, 255.2031, 255.2032, 
    255.2031, 255.203, 255.203, 255.2028, 255.2029, 255.2025, 255.2027, 
    255.2022, 255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.203, 255.2031, 255.2031, 255.2032, 255.2031, 255.2031, 255.203, 
    255.2029, 255.2029, 255.2028, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2023, 255.2023, 255.202, 255.2022, 255.2019, 
    255.2019, 255.2021, 255.2019, 255.203, 255.203, 255.2032, 255.2031, 
    255.2032, 255.2031, 255.2031, 255.2029, 255.2029, 255.2028, 255.2027, 
    255.2027, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2022, 
    255.2022, 255.2021, 255.2021, 255.2022, 255.2019, 255.202, 255.2019, 
    255.202, 255.203, 255.203, 255.203, 255.203, 255.203, 255.2028, 255.2028, 
    255.2026, 255.2027, 255.2025, 255.2026, 255.2026, 255.2025, 255.2026, 
    255.2023, 255.2025, 255.2022, 255.2024, 255.2021, 255.2022, 255.2021, 
    255.2021, 255.202, 255.2019, 255.2019, 255.2018, 255.2029, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2025, 255.2024, 
    255.2023, 255.2025, 255.2024, 255.2028, 255.2027, 255.2028, 255.2029, 
    255.2025, 255.2027, 255.2023, 255.2024, 255.2021, 255.2022, 255.2019, 
    255.2018, 255.2016, 255.2015, 255.2028, 255.2029, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2024, 255.2024, 255.2023, 255.2022, 255.2024, 
    255.2022, 255.2027, 255.2025, 255.2029, 255.2028, 255.2027, 255.2027, 
    255.2025, 255.2025, 255.2023, 255.2024, 255.2018, 255.2021, 255.2013, 
    255.2015, 255.2029, 255.2028, 255.2026, 255.2027, 255.2024, 255.2023, 
    255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.2021, 255.2024, 
    255.2023, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 255.2024, 
    255.2024, 255.2023, 255.2022, 255.2024, 255.2018, 255.2022, 255.2027, 
    255.2026, 255.2026, 255.2027, 255.2023, 255.2025, 255.2021, 255.2022, 
    255.2021, 255.2021, 255.2022, 255.2023, 255.2023, 255.2025, 255.2026, 
    255.2027, 255.2026, 255.2025, 255.2023, 255.2022, 255.2022, 255.2021, 
    255.2024, 255.2023, 255.2023, 255.2022, 255.2025, 255.2023, 255.2026, 
    255.2025, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2023, 
    255.2024, 255.2025, 255.2025, 255.2025, 255.2026, 255.2025, 255.2025, 
    255.2023, 255.2022, 255.2021, 255.202, 255.2019, 255.202, 255.2018, 
    255.202, 255.2016, 255.2022, 255.202, 255.2025, 255.2024, 255.2023, 
    255.2021, 255.2022, 255.2021, 255.2024, 255.2025, 255.2026, 255.2026, 
    255.2026, 255.2026, 255.2025, 255.2025, 255.2023, 255.2024, 255.2022, 
    255.2021, 255.2018, 255.2016, 255.2014, 255.2014, 255.2013, 255.2013 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  255.2032, 255.203, 255.2031, 255.203, 255.203, 255.2029, 255.2032, 255.203, 
    255.2031, 255.2032, 255.2027, 255.2029, 255.2025, 255.2026, 255.2022, 
    255.2025, 255.2022, 255.2022, 255.2021, 255.2021, 255.2019, 255.202, 
    255.2018, 255.2019, 255.2019, 255.202, 255.2029, 255.2028, 255.2029, 
    255.2029, 255.2029, 255.203, 255.2031, 255.2032, 255.2032, 255.2031, 
    255.2029, 255.2029, 255.2028, 255.2028, 255.2026, 255.2027, 255.2023, 
    255.2024, 255.2021, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2022, 255.2023, 255.2026, 255.2025, 255.2029, 255.203, 255.2032, 
    255.2032, 255.2032, 255.2032, 255.2031, 255.203, 255.2029, 255.2028, 
    255.2028, 255.2026, 255.2025, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2021, 255.2021, 255.2021, 255.2023, 255.2021, 255.2023, 255.2023, 
    255.2028, 255.2029, 255.203, 255.2031, 255.2032, 255.2031, 255.2032, 
    255.2031, 255.203, 255.203, 255.2028, 255.2029, 255.2025, 255.2027, 
    255.2022, 255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.203, 255.2031, 255.2031, 255.2032, 255.2031, 255.2031, 255.203, 
    255.2029, 255.2029, 255.2028, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2023, 255.2023, 255.202, 255.2022, 255.2019, 
    255.2019, 255.2021, 255.2019, 255.203, 255.203, 255.2032, 255.2031, 
    255.2032, 255.2031, 255.2031, 255.2029, 255.2029, 255.2028, 255.2027, 
    255.2027, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2022, 
    255.2022, 255.2021, 255.2021, 255.2022, 255.2019, 255.202, 255.2019, 
    255.202, 255.203, 255.203, 255.203, 255.203, 255.203, 255.2028, 255.2028, 
    255.2026, 255.2027, 255.2025, 255.2026, 255.2026, 255.2025, 255.2026, 
    255.2023, 255.2025, 255.2022, 255.2024, 255.2021, 255.2022, 255.2021, 
    255.2021, 255.202, 255.2019, 255.2019, 255.2018, 255.2029, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2025, 255.2024, 
    255.2023, 255.2025, 255.2024, 255.2028, 255.2027, 255.2028, 255.2029, 
    255.2025, 255.2027, 255.2023, 255.2024, 255.2021, 255.2022, 255.2019, 
    255.2018, 255.2016, 255.2015, 255.2028, 255.2029, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2024, 255.2024, 255.2023, 255.2022, 255.2024, 
    255.2022, 255.2027, 255.2025, 255.2029, 255.2028, 255.2027, 255.2027, 
    255.2025, 255.2025, 255.2023, 255.2024, 255.2018, 255.2021, 255.2013, 
    255.2015, 255.2029, 255.2028, 255.2026, 255.2027, 255.2024, 255.2023, 
    255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.2021, 255.2024, 
    255.2023, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 255.2024, 
    255.2024, 255.2023, 255.2022, 255.2024, 255.2018, 255.2022, 255.2027, 
    255.2026, 255.2026, 255.2027, 255.2023, 255.2025, 255.2021, 255.2022, 
    255.2021, 255.2021, 255.2022, 255.2023, 255.2023, 255.2025, 255.2026, 
    255.2027, 255.2026, 255.2025, 255.2023, 255.2022, 255.2022, 255.2021, 
    255.2024, 255.2023, 255.2023, 255.2022, 255.2025, 255.2023, 255.2026, 
    255.2025, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2023, 
    255.2024, 255.2025, 255.2025, 255.2025, 255.2026, 255.2025, 255.2025, 
    255.2023, 255.2022, 255.2021, 255.202, 255.2019, 255.202, 255.2018, 
    255.202, 255.2016, 255.2022, 255.202, 255.2025, 255.2024, 255.2023, 
    255.2021, 255.2022, 255.2021, 255.2024, 255.2025, 255.2026, 255.2026, 
    255.2026, 255.2026, 255.2025, 255.2025, 255.2023, 255.2024, 255.2022, 
    255.2021, 255.2018, 255.2016, 255.2014, 255.2014, 255.2013, 255.2013 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  253.6898, 253.6917, 253.6913, 253.6929, 253.692, 253.693, 253.6902, 
    253.6918, 253.6908, 253.69, 253.6958, 253.6929, 253.6988, 253.697, 
    253.7016, 253.6985, 253.7023, 253.7016, 253.7037, 253.7031, 253.7058, 
    253.704, 253.7072, 253.7054, 253.7057, 253.7039, 253.6935, 253.6954, 
    253.6934, 253.6937, 253.6936, 253.692, 253.6913, 253.6897, 253.69, 
    253.6911, 253.6938, 253.6929, 253.6952, 253.6952, 253.6977, 253.6966, 
    253.7008, 253.6996, 253.7031, 253.7023, 253.7031, 253.7028, 253.7031, 
    253.7018, 253.7023, 253.7012, 253.6968, 253.6981, 253.6942, 253.6918, 
    253.6903, 253.6892, 253.6893, 253.6896, 253.6911, 253.6926, 253.6937, 
    253.6944, 253.6952, 253.6973, 253.6985, 253.701, 253.7006, 253.7014, 
    253.7022, 253.7034, 253.7032, 253.7038, 253.7014, 253.703, 253.7004, 
    253.7011, 253.6952, 253.6932, 253.6922, 253.6914, 253.6895, 253.6908, 
    253.6903, 253.6916, 253.6924, 253.692, 253.6945, 253.6935, 253.6985, 
    253.6964, 253.7021, 253.7007, 253.7024, 253.7015, 253.703, 253.7017, 
    253.704, 253.7045, 253.7041, 253.7055, 253.7016, 253.7031, 253.692, 
    253.692, 253.6923, 253.691, 253.6909, 253.6897, 253.6908, 253.6912, 
    253.6924, 253.6931, 253.6938, 253.6953, 253.6969, 253.6991, 253.7008, 
    253.7019, 253.7012, 253.7018, 253.7012, 253.7009, 253.7043, 253.7023, 
    253.7053, 253.7051, 253.7038, 253.7051, 253.6921, 253.6917, 253.6904, 
    253.6914, 253.6895, 253.6906, 253.6912, 253.6935, 253.694, 253.6945, 
    253.6954, 253.6966, 253.6987, 253.7005, 253.7022, 253.7021, 253.7021, 
    253.7025, 253.7016, 253.7027, 253.7028, 253.7024, 253.7051, 253.7043, 
    253.7051, 253.7046, 253.6918, 253.6925, 253.6921, 253.6927, 253.6923, 
    253.6943, 253.6949, 253.6977, 253.6966, 253.6984, 253.6968, 253.6971, 
    253.6984, 253.6969, 253.7004, 253.698, 253.7025, 253.7, 253.7027, 
    253.7022, 253.703, 253.7037, 253.7045, 253.7061, 253.7058, 253.7071, 
    253.6934, 253.6942, 253.6942, 253.695, 253.6956, 253.697, 253.6992, 
    253.6984, 253.6999, 253.7002, 253.6979, 253.6993, 253.6948, 253.6955, 
    253.6951, 253.6935, 253.6986, 253.6959, 253.7008, 253.6994, 253.7036, 
    253.7015, 253.7056, 253.7072, 253.709, 253.7108, 253.6947, 253.6941, 
    253.6951, 253.6965, 253.6978, 253.6995, 253.6997, 253.7, 253.7008, 
    253.7015, 253.7001, 253.7017, 253.6956, 253.6988, 253.6939, 253.6953, 
    253.6964, 253.696, 253.6983, 253.6989, 253.7011, 253.7, 253.7068, 
    253.7038, 253.7123, 253.7099, 253.6939, 253.6947, 253.6973, 253.696, 
    253.6996, 253.7005, 253.7012, 253.7021, 253.7022, 253.7027, 253.7019, 
    253.7027, 253.6995, 253.7009, 253.697, 253.6979, 253.6975, 253.697, 
    253.6985, 253.7001, 253.7001, 253.7006, 253.702, 253.6996, 253.7071, 
    253.7024, 253.6955, 253.6969, 253.6971, 253.6966, 253.7004, 253.699, 
    253.7027, 253.7017, 253.7034, 253.7025, 253.7024, 253.7014, 253.7007, 
    253.6991, 253.6977, 253.6967, 253.6969, 253.6981, 253.7002, 253.7022, 
    253.7018, 253.7032, 253.6993, 253.701, 253.7003, 253.702, 253.6984, 
    253.7013, 253.6976, 253.698, 253.699, 253.701, 253.7016, 253.702, 
    253.7018, 253.7002, 253.7, 253.699, 253.6987, 253.6979, 253.6972, 
    253.6978, 253.6984, 253.7003, 253.7019, 253.7037, 253.7041, 253.7061, 
    253.7044, 253.7072, 253.7048, 253.7089, 253.7016, 253.7048, 253.699, 
    253.6997, 253.7008, 253.7033, 253.702, 253.7036, 253.7, 253.6981, 
    253.6976, 253.6967, 253.6977, 253.6976, 253.6985, 253.6982, 253.7003, 
    253.6992, 253.7024, 253.7036, 253.707, 253.709, 253.7111, 253.7121, 
    253.7124, 253.7125,
  255.2211, 255.2229, 255.2225, 255.2239, 255.2231, 255.2241, 255.2215, 
    255.2229, 255.222, 255.2213, 255.2266, 255.224, 255.2295, 255.2278, 
    255.2321, 255.2292, 255.2327, 255.232, 255.2341, 255.2335, 255.236, 
    255.2343, 255.2374, 255.2356, 255.2359, 255.2343, 255.2245, 255.2263, 
    255.2244, 255.2247, 255.2246, 255.2232, 255.2224, 255.221, 255.2212, 
    255.2223, 255.2248, 255.224, 255.2261, 255.2261, 255.2284, 255.2274, 
    255.2313, 255.2302, 255.2335, 255.2327, 255.2335, 255.2332, 255.2335, 
    255.2322, 255.2328, 255.2317, 255.2275, 255.2288, 255.2251, 255.2229, 
    255.2215, 255.2205, 255.2206, 255.2209, 255.2223, 255.2237, 255.2247, 
    255.2254, 255.2261, 255.228, 255.2291, 255.2316, 255.2311, 255.2319, 
    255.2326, 255.2338, 255.2336, 255.2341, 255.2319, 255.2333, 255.2309, 
    255.2316, 255.2261, 255.2242, 255.2233, 255.2226, 255.2207, 255.222, 
    255.2215, 255.2227, 255.2235, 255.2231, 255.2254, 255.2245, 255.2292, 
    255.2272, 255.2325, 255.2312, 255.2328, 255.232, 255.2334, 255.2321, 
    255.2343, 255.2348, 255.2345, 255.2357, 255.2321, 255.2334, 255.2231, 
    255.2231, 255.2234, 255.2222, 255.2221, 255.221, 255.222, 255.2224, 
    255.2235, 255.2242, 255.2248, 255.2261, 255.2276, 255.2298, 255.2313, 
    255.2323, 255.2317, 255.2323, 255.2316, 255.2314, 255.2346, 255.2328, 
    255.2355, 255.2354, 255.2341, 255.2354, 255.2232, 255.2228, 255.2216, 
    255.2226, 255.2208, 255.2218, 255.2223, 255.2245, 255.225, 255.2254, 
    255.2263, 255.2274, 255.2294, 255.231, 255.2326, 255.2325, 255.2326, 
    255.2329, 255.232, 255.233, 255.2332, 255.2328, 255.2354, 255.2346, 
    255.2354, 255.2349, 255.2229, 255.2235, 255.2232, 255.2238, 255.2234, 
    255.2252, 255.2258, 255.2284, 255.2274, 255.2291, 255.2276, 255.2278, 
    255.2291, 255.2276, 255.2309, 255.2287, 255.2329, 255.2306, 255.2331, 
    255.2326, 255.2334, 255.234, 255.2348, 255.2363, 255.236, 255.2372, 
    255.2244, 255.2252, 255.2251, 255.2259, 255.2265, 255.2278, 255.2298, 
    255.2291, 255.2305, 255.2308, 255.2286, 255.2299, 255.2257, 255.2263, 
    255.226, 255.2245, 255.2292, 255.2268, 255.2313, 255.23, 255.2339, 
    255.2319, 255.2358, 255.2374, 255.239, 255.2407, 255.2256, 255.2251, 
    255.226, 255.2273, 255.2285, 255.2301, 255.2303, 255.2305, 255.2313, 
    255.232, 255.2306, 255.2321, 255.2265, 255.2294, 255.2249, 255.2262, 
    255.2272, 255.2268, 255.229, 255.2295, 255.2316, 255.2305, 255.237, 
    255.2341, 255.2421, 255.2399, 255.2249, 255.2256, 255.228, 255.2269, 
    255.2302, 255.231, 255.2317, 255.2325, 255.2326, 255.2331, 255.2323, 
    255.2331, 255.2301, 255.2314, 255.2278, 255.2286, 255.2282, 255.2278, 
    255.2292, 255.2306, 255.2307, 255.2312, 255.2324, 255.2302, 255.2373, 
    255.2328, 255.2264, 255.2277, 255.2279, 255.2274, 255.2309, 255.2296, 
    255.2331, 255.2322, 255.2337, 255.233, 255.2328, 255.2319, 255.2312, 
    255.2297, 255.2284, 255.2275, 255.2277, 255.2288, 255.2307, 255.2326, 
    255.2322, 255.2336, 255.2299, 255.2315, 255.2309, 255.2324, 255.229, 
    255.2318, 255.2283, 255.2286, 255.2296, 255.2315, 255.232, 255.2325, 
    255.2322, 255.2308, 255.2306, 255.2296, 255.2293, 255.2286, 255.228, 
    255.2285, 255.2291, 255.2308, 255.2323, 255.234, 255.2344, 255.2363, 
    255.2347, 255.2373, 255.235, 255.239, 255.232, 255.235, 255.2297, 
    255.2303, 255.2313, 255.2337, 255.2324, 255.2339, 255.2306, 255.2288, 
    255.2284, 255.2275, 255.2284, 255.2283, 255.2291, 255.2289, 255.2309, 
    255.2298, 255.2328, 255.2339, 255.2371, 255.239, 255.241, 255.2419, 
    255.2422, 255.2423,
  257.287, 257.2885, 257.2882, 257.2893, 257.2887, 257.2894, 257.2874, 
    257.2885, 257.2878, 257.2872, 257.2915, 257.2894, 257.2938, 257.2924, 
    257.2959, 257.2936, 257.2964, 257.2959, 257.2975, 257.2971, 257.2991, 
    257.2978, 257.3003, 257.2988, 257.299, 257.2977, 257.2898, 257.2912, 
    257.2897, 257.2899, 257.2899, 257.2887, 257.2881, 257.287, 257.2872, 
    257.288, 257.29, 257.2894, 257.2911, 257.291, 257.293, 257.2921, 
    257.2953, 257.2944, 257.2971, 257.2964, 257.2971, 257.2969, 257.2971, 
    257.2961, 257.2965, 257.2956, 257.2922, 257.2932, 257.2903, 257.2885, 
    257.2874, 257.2866, 257.2867, 257.2869, 257.288, 257.2891, 257.2899, 
    257.2905, 257.291, 257.2926, 257.2935, 257.2955, 257.2952, 257.2957, 
    257.2964, 257.2973, 257.2971, 257.2976, 257.2957, 257.297, 257.295, 
    257.2955, 257.2911, 257.2896, 257.2888, 257.2882, 257.2868, 257.2878, 
    257.2874, 257.2884, 257.2889, 257.2887, 257.2905, 257.2898, 257.2936, 
    257.2919, 257.2963, 257.2952, 257.2965, 257.2959, 257.297, 257.296, 
    257.2978, 257.2981, 257.2979, 257.2989, 257.2959, 257.2971, 257.2886, 
    257.2887, 257.2889, 257.2879, 257.2878, 257.287, 257.2878, 257.2881, 
    257.289, 257.2895, 257.29, 257.2911, 257.2923, 257.294, 257.2953, 
    257.2961, 257.2956, 257.2961, 257.2956, 257.2953, 257.298, 257.2965, 
    257.2987, 257.2986, 257.2976, 257.2986, 257.2887, 257.2885, 257.2875, 
    257.2882, 257.2869, 257.2876, 257.2881, 257.2898, 257.2902, 257.2905, 
    257.2912, 257.2921, 257.2937, 257.2951, 257.2964, 257.2963, 257.2963, 
    257.2966, 257.2959, 257.2967, 257.2968, 257.2965, 257.2986, 257.298, 
    257.2986, 257.2982, 257.2885, 257.289, 257.2888, 257.2892, 257.2889, 
    257.2904, 257.2908, 257.293, 257.2921, 257.2935, 257.2923, 257.2925, 
    257.2935, 257.2923, 257.295, 257.2932, 257.2966, 257.2947, 257.2967, 
    257.2964, 257.297, 257.2975, 257.2982, 257.2994, 257.2991, 257.3001, 
    257.2897, 257.2903, 257.2903, 257.2909, 257.2914, 257.2924, 257.2941, 
    257.2935, 257.2946, 257.2949, 257.2931, 257.2942, 257.2907, 257.2913, 
    257.291, 257.2898, 257.2936, 257.2916, 257.2953, 257.2943, 257.2974, 
    257.2958, 257.299, 257.3003, 257.3016, 257.303, 257.2907, 257.2903, 
    257.291, 257.292, 257.293, 257.2943, 257.2944, 257.2947, 257.2953, 
    257.2958, 257.2947, 257.296, 257.2914, 257.2938, 257.2901, 257.2912, 
    257.292, 257.2916, 257.2934, 257.2939, 257.2955, 257.2947, 257.2999, 
    257.2976, 257.3042, 257.3023, 257.2901, 257.2907, 257.2926, 257.2917, 
    257.2944, 257.295, 257.2956, 257.2963, 257.2964, 257.2968, 257.2961, 
    257.2968, 257.2943, 257.2954, 257.2924, 257.2931, 257.2928, 257.2924, 
    257.2936, 257.2948, 257.2948, 257.2952, 257.2962, 257.2944, 257.3002, 
    257.2966, 257.2913, 257.2924, 257.2925, 257.2921, 257.295, 257.2939, 
    257.2968, 257.296, 257.2973, 257.2966, 257.2965, 257.2957, 257.2953, 
    257.294, 257.293, 257.2922, 257.2924, 257.2932, 257.2948, 257.2964, 
    257.296, 257.2972, 257.2942, 257.2954, 257.295, 257.2962, 257.2935, 
    257.2957, 257.2929, 257.2932, 257.2939, 257.2955, 257.2959, 257.2963, 
    257.296, 257.2949, 257.2947, 257.2939, 257.2937, 257.2931, 257.2926, 
    257.293, 257.2935, 257.2949, 257.2961, 257.2975, 257.2979, 257.2994, 
    257.2981, 257.3002, 257.2984, 257.3016, 257.2959, 257.2983, 257.294, 
    257.2944, 257.2953, 257.2972, 257.2962, 257.2975, 257.2947, 257.2932, 
    257.2929, 257.2922, 257.2929, 257.2929, 257.2935, 257.2933, 257.295, 
    257.2941, 257.2965, 257.2975, 257.3, 257.3016, 257.3033, 257.304, 
    257.3042, 257.3043,
  259.794, 259.7949, 259.7947, 259.7953, 259.795, 259.7954, 259.7942, 
    259.7949, 259.7944, 259.7941, 259.7966, 259.7954, 259.798, 259.7972, 
    259.7993, 259.7979, 259.7996, 259.7993, 259.8002, 259.8, 259.8012, 
    259.8004, 259.8019, 259.801, 259.8011, 259.8004, 259.7957, 259.7965, 
    259.7956, 259.7957, 259.7957, 259.795, 259.7946, 259.794, 259.7941, 
    259.7946, 259.7958, 259.7954, 259.7964, 259.7964, 259.7975, 259.797, 
    259.7989, 259.7984, 259.8, 259.7996, 259.8, 259.7998, 259.8, 259.7993, 
    259.7996, 259.7991, 259.7971, 259.7976, 259.7959, 259.7949, 259.7942, 
    259.7938, 259.7938, 259.7939, 259.7946, 259.7952, 259.7957, 259.7961, 
    259.7964, 259.7973, 259.7978, 259.799, 259.7988, 259.7992, 259.7995, 
    259.8001, 259.8, 259.8003, 259.7992, 259.7999, 259.7987, 259.799, 
    259.7964, 259.7955, 259.795, 259.7947, 259.7939, 259.7945, 259.7942, 
    259.7948, 259.7951, 259.795, 259.7961, 259.7956, 259.7979, 259.7969, 
    259.7995, 259.7989, 259.7996, 259.7992, 259.7999, 259.7993, 259.8004, 
    259.8006, 259.8004, 259.8011, 259.7993, 259.7999, 259.795, 259.795, 
    259.7951, 259.7945, 259.7945, 259.794, 259.7944, 259.7946, 259.7952, 
    259.7955, 259.7957, 259.7964, 259.7971, 259.7981, 259.7989, 259.7994, 
    259.7991, 259.7993, 259.799, 259.7989, 259.8005, 259.7996, 259.801, 
    259.8009, 259.8003, 259.8009, 259.795, 259.7948, 259.7943, 259.7947, 
    259.7939, 259.7943, 259.7946, 259.7956, 259.7959, 259.7961, 259.7965, 
    259.797, 259.7979, 259.7988, 259.7995, 259.7995, 259.7995, 259.7997, 
    259.7993, 259.7997, 259.7998, 259.7996, 259.8009, 259.8005, 259.8009, 
    259.8007, 259.7949, 259.7952, 259.795, 259.7953, 259.7951, 259.796, 
    259.7962, 259.7975, 259.797, 259.7978, 259.7971, 259.7972, 259.7978, 
    259.7971, 259.7987, 259.7976, 259.7997, 259.7986, 259.7997, 259.7995, 
    259.7999, 259.8002, 259.8006, 259.8014, 259.8012, 259.8018, 259.7956, 
    259.7959, 259.7959, 259.7963, 259.7966, 259.7972, 259.7982, 259.7978, 
    259.7985, 259.7986, 259.7976, 259.7982, 259.7962, 259.7965, 259.7963, 
    259.7956, 259.7979, 259.7967, 259.7989, 259.7982, 259.8002, 259.7992, 
    259.8011, 259.8019, 259.8027, 259.8036, 259.7961, 259.7959, 259.7964, 
    259.7969, 259.7975, 259.7983, 259.7984, 259.7985, 259.7989, 259.7992, 
    259.7986, 259.7993, 259.7966, 259.798, 259.7958, 259.7964, 259.7969, 
    259.7967, 259.7978, 259.798, 259.799, 259.7985, 259.8017, 259.8003, 
    259.8043, 259.8032, 259.7958, 259.7961, 259.7973, 259.7968, 259.7983, 
    259.7987, 259.7991, 259.7995, 259.7995, 259.7998, 259.7994, 259.7998, 
    259.7983, 259.799, 259.7972, 259.7976, 259.7974, 259.7972, 259.7979, 
    259.7986, 259.7986, 259.7988, 259.7994, 259.7984, 259.8018, 259.7997, 
    259.7965, 259.7971, 259.7972, 259.797, 259.7987, 259.7981, 259.7998, 
    259.7993, 259.8001, 259.7997, 259.7997, 259.7992, 259.7989, 259.7981, 
    259.7975, 259.797, 259.7971, 259.7977, 259.7986, 259.7995, 259.7993, 
    259.8, 259.7982, 259.799, 259.7987, 259.7994, 259.7978, 259.7992, 
    259.7975, 259.7976, 259.7981, 259.799, 259.7992, 259.7995, 259.7993, 
    259.7986, 259.7985, 259.7981, 259.7979, 259.7976, 259.7973, 259.7975, 
    259.7978, 259.7986, 259.7994, 259.8002, 259.8004, 259.8014, 259.8006, 
    259.8018, 259.8007, 259.8027, 259.7993, 259.8007, 259.7981, 259.7984, 
    259.7989, 259.8001, 259.7994, 259.8002, 259.7985, 259.7977, 259.7975, 
    259.7971, 259.7975, 259.7975, 259.7979, 259.7977, 259.7987, 259.7982, 
    259.7996, 259.8002, 259.8018, 259.8027, 259.8037, 259.8042, 259.8043, 
    259.8044,
  262.0097, 262.0099, 262.0099, 262.0101, 262.01, 262.0101, 262.0098, 
    262.0099, 262.0098, 262.0097, 262.0104, 262.0101, 262.0108, 262.0106, 
    262.0111, 262.0107, 262.0112, 262.0111, 262.0114, 262.0113, 262.0117, 
    262.0114, 262.0119, 262.0116, 262.0117, 262.0114, 262.0101, 262.0103, 
    262.0101, 262.0102, 262.0101, 262.01, 262.0099, 262.0097, 262.0097, 
    262.0099, 262.0102, 262.0101, 262.0103, 262.0103, 262.0106, 262.0105, 
    262.011, 262.0109, 262.0113, 262.0112, 262.0113, 262.0113, 262.0113, 
    262.0111, 262.0112, 262.0111, 262.0105, 262.0107, 262.0102, 262.0099, 
    262.0098, 262.0096, 262.0097, 262.0097, 262.0099, 262.01, 262.0102, 
    262.0103, 262.0103, 262.0106, 262.0107, 262.011, 262.011, 262.0111, 
    262.0112, 262.0114, 262.0113, 262.0114, 262.0111, 262.0113, 262.011, 
    262.011, 262.0103, 262.0101, 262.01, 262.0099, 262.0097, 262.0098, 
    262.0098, 262.0099, 262.01, 262.0099, 262.0103, 262.0101, 262.0107, 
    262.0105, 262.0112, 262.011, 262.0112, 262.0111, 262.0113, 262.0111, 
    262.0114, 262.0115, 262.0114, 262.0116, 262.0111, 262.0113, 262.0099, 
    262.01, 262.01, 262.0099, 262.0098, 262.0097, 262.0098, 262.0099, 262.01, 
    262.0101, 262.0102, 262.0103, 262.0105, 262.0108, 262.011, 262.0112, 
    262.0111, 262.0111, 262.0111, 262.011, 262.0115, 262.0112, 262.0116, 
    262.0116, 262.0114, 262.0116, 262.01, 262.0099, 262.0098, 262.0099, 
    262.0097, 262.0098, 262.0099, 262.0101, 262.0102, 262.0103, 262.0103, 
    262.0105, 262.0107, 262.011, 262.0112, 262.0112, 262.0112, 262.0112, 
    262.0111, 262.0113, 262.0113, 262.0112, 262.0116, 262.0115, 262.0116, 
    262.0115, 262.0099, 262.01, 262.01, 262.01, 262.01, 262.0102, 262.0103, 
    262.0106, 262.0105, 262.0107, 262.0105, 262.0106, 262.0107, 262.0105, 
    262.011, 262.0107, 262.0112, 262.0109, 262.0113, 262.0112, 262.0113, 
    262.0114, 262.0115, 262.0117, 262.0117, 262.0119, 262.0101, 262.0102, 
    262.0102, 262.0103, 262.0104, 262.0106, 262.0108, 262.0107, 262.0109, 
    262.011, 262.0107, 262.0108, 262.0103, 262.0104, 262.0103, 262.0101, 
    262.0107, 262.0104, 262.011, 262.0108, 262.0114, 262.0111, 262.0117, 
    262.0119, 262.0121, 262.0124, 262.0103, 262.0102, 262.0103, 262.0105, 
    262.0107, 262.0109, 262.0109, 262.0109, 262.011, 262.0111, 262.0109, 
    262.0111, 262.0104, 262.0108, 262.0102, 262.0103, 262.0105, 262.0104, 
    262.0107, 262.0108, 262.011, 262.0109, 262.0118, 262.0114, 262.0126, 
    262.0123, 262.0102, 262.0103, 262.0106, 262.0104, 262.0109, 262.011, 
    262.0111, 262.0112, 262.0112, 262.0113, 262.0112, 262.0113, 262.0109, 
    262.011, 262.0106, 262.0107, 262.0106, 262.0106, 262.0107, 262.0109, 
    262.0109, 262.011, 262.0112, 262.0109, 262.0119, 262.0112, 262.0104, 
    262.0105, 262.0106, 262.0105, 262.011, 262.0108, 262.0113, 262.0111, 
    262.0114, 262.0112, 262.0112, 262.0111, 262.011, 262.0108, 262.0106, 
    262.0105, 262.0105, 262.0107, 262.0109, 262.0112, 262.0111, 262.0113, 
    262.0108, 262.011, 262.011, 262.0112, 262.0107, 262.0111, 262.0106, 
    262.0107, 262.0108, 262.011, 262.0111, 262.0112, 262.0111, 262.011, 
    262.0109, 262.0108, 262.0107, 262.0107, 262.0106, 262.0107, 262.0107, 
    262.011, 262.0112, 262.0114, 262.0114, 262.0117, 262.0115, 262.0119, 
    262.0115, 262.0121, 262.0111, 262.0115, 262.0108, 262.0109, 262.011, 
    262.0114, 262.0112, 262.0114, 262.0109, 262.0107, 262.0106, 262.0105, 
    262.0106, 262.0106, 262.0107, 262.0107, 262.011, 262.0108, 262.0112, 
    262.0114, 262.0118, 262.0121, 262.0125, 262.0126, 262.0126, 262.0126,
  262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985,
  263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.1129, 263.1252, 263.1229, 263.1328, 263.1273, 263.1338, 263.1154, 
    263.1257, 263.1191, 263.114, 263.1519, 263.1332, 263.1713, 263.1594, 
    263.1892, 263.1694, 263.1932, 263.1887, 263.2022, 263.1984, 263.2156, 
    263.204, 263.2245, 263.2129, 263.2147, 263.2036, 263.137, 263.1495, 
    263.1363, 263.1381, 263.1373, 263.1274, 263.1224, 263.112, 263.1139, 
    263.1215, 263.1389, 263.133, 263.1478, 263.1475, 263.1638, 263.1564, 
    263.1839, 263.1761, 263.1985, 263.193, 263.1983, 263.1967, 263.1983, 
    263.1901, 263.1936, 263.1863, 263.1578, 263.1662, 263.1411, 263.1259, 
    263.1159, 263.1087, 263.1097, 263.1116, 263.1216, 263.1309, 263.138, 
    263.1428, 263.1474, 263.1614, 263.1689, 263.1855, 263.1825, 263.1876, 
    263.1924, 263.2004, 263.1991, 263.2026, 263.1874, 263.1975, 263.1808, 
    263.1854, 263.1486, 263.1346, 263.1285, 263.1233, 263.1105, 263.1193, 
    263.1158, 263.1242, 263.1294, 263.1268, 263.1429, 263.1367, 263.1693, 
    263.1553, 263.1918, 263.1831, 263.1939, 263.1884, 263.1978, 263.1894, 
    263.2039, 263.2071, 263.2049, 263.2133, 263.1889, 263.1983, 263.1267, 
    263.1272, 263.1292, 263.1204, 263.1199, 263.1119, 263.119, 263.122, 
    263.1297, 263.1343, 263.1386, 263.148, 263.1585, 263.1732, 263.1837, 
    263.1907, 263.1864, 263.1902, 263.1859, 263.184, 263.2059, 263.1936, 
    263.212, 263.211, 263.2027, 263.2112, 263.1275, 263.125, 263.1165, 
    263.1232, 263.1111, 263.1178, 263.1217, 263.1367, 263.1401, 263.1431, 
    263.1491, 263.1568, 263.1703, 263.182, 263.1927, 263.1919, 263.1922, 
    263.1945, 263.1887, 263.1955, 263.1966, 263.1936, 263.2109, 263.206, 
    263.211, 263.2078, 263.1258, 263.1299, 263.1277, 263.1319, 263.1289, 
    263.142, 263.1459, 263.1641, 263.1567, 263.1685, 263.1579, 263.1598, 
    263.1689, 263.1585, 263.1813, 263.1658, 263.1946, 263.1791, 263.1956, 
    263.1926, 263.1975, 263.2019, 263.2074, 263.2175, 263.2151, 263.2236, 
    263.1361, 263.1414, 263.1409, 263.1465, 263.1506, 263.1595, 263.1737, 
    263.1683, 263.1781, 263.1801, 263.1652, 263.1743, 263.1449, 263.1497, 
    263.1469, 263.1365, 263.1695, 263.1526, 263.1838, 263.1747, 263.2012, 
    263.1881, 263.2138, 263.2247, 263.2351, 263.247, 263.1443, 263.1407, 
    263.1471, 263.156, 263.1643, 263.1753, 263.1764, 263.1784, 263.1837, 
    263.1882, 263.1791, 263.1893, 263.1507, 263.171, 263.1393, 263.1488, 
    263.1555, 263.1526, 263.1677, 263.1713, 263.1857, 263.1783, 263.222, 
    263.2028, 263.2562, 263.2413, 263.1394, 263.1443, 263.1611, 263.1531, 
    263.176, 263.1816, 263.1862, 263.192, 263.1926, 263.196, 263.1904, 
    263.1958, 263.1753, 263.1845, 263.1592, 263.1654, 263.1625, 263.1594, 
    263.169, 263.1792, 263.1795, 263.1827, 263.1918, 263.1761, 263.2245, 
    263.1947, 263.1496, 263.1588, 263.1602, 263.1566, 263.1811, 263.1722, 
    263.196, 263.1896, 263.2, 263.1948, 263.1941, 263.1874, 263.1832, 
    263.1726, 263.164, 263.1571, 263.1587, 263.1662, 263.1798, 263.1927, 
    263.1899, 263.1992, 263.1743, 263.1848, 263.1808, 263.1913, 263.1682, 
    263.1878, 263.1631, 263.1653, 263.172, 263.1855, 263.1885, 263.1917, 
    263.1897, 263.1802, 263.1786, 263.1719, 263.17, 263.1648, 263.1606, 
    263.1645, 263.1685, 263.1802, 263.1907, 263.2019, 263.2047, 263.2177, 
    263.2071, 263.2246, 263.2096, 263.2356, 263.189, 263.2093, 263.1723, 
    263.1764, 263.1836, 263.2001, 263.1913, 263.2016, 263.1786, 263.1665, 
    263.1634, 263.1575, 263.1635, 263.163, 263.1687, 263.1669, 263.1806, 
    263.1732, 263.194, 263.2015, 263.2227, 263.2356, 263.2488, 263.2546, 
    263.2563, 263.2571 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9098, 253.9106, 253.9105, 253.9111, 253.9108, 253.9112, 253.91, 
    253.9107, 253.9102, 253.9099, 253.9124, 253.9112, 253.9138, 253.913, 
    253.9151, 253.9137, 253.9153, 253.915, 253.916, 253.9157, 253.9169, 
    253.9161, 253.9175, 253.9167, 253.9168, 253.9161, 253.9115, 253.9123, 
    253.9114, 253.9115, 253.9115, 253.9108, 253.9104, 253.9097, 253.9099, 
    253.9104, 253.9116, 253.9112, 253.9122, 253.9122, 253.9133, 253.9128, 
    253.9147, 253.9142, 253.9157, 253.9153, 253.9157, 253.9156, 253.9157, 
    253.9151, 253.9154, 253.9149, 253.9129, 253.9135, 253.9117, 253.9107, 
    253.91, 253.9095, 253.9096, 253.9097, 253.9104, 253.911, 253.9115, 
    253.9118, 253.9122, 253.9131, 253.9137, 253.9148, 253.9146, 253.9149, 
    253.9153, 253.9158, 253.9158, 253.916, 253.9149, 253.9156, 253.9145, 
    253.9148, 253.9122, 253.9113, 253.9108, 253.9105, 253.9096, 253.9102, 
    253.91, 253.9106, 253.9109, 253.9108, 253.9119, 253.9114, 253.9137, 
    253.9127, 253.9153, 253.9146, 253.9154, 253.915, 253.9157, 253.9151, 
    253.9161, 253.9163, 253.9162, 253.9168, 253.9151, 253.9157, 253.9107, 
    253.9108, 253.9109, 253.9103, 253.9103, 253.9097, 253.9102, 253.9104, 
    253.9109, 253.9113, 253.9116, 253.9122, 253.9129, 253.914, 253.9147, 
    253.9152, 253.9149, 253.9151, 253.9148, 253.9147, 253.9162, 253.9154, 
    253.9167, 253.9166, 253.916, 253.9166, 253.9108, 253.9106, 253.91, 
    253.9105, 253.9097, 253.9101, 253.9104, 253.9114, 253.9117, 253.9119, 
    253.9123, 253.9128, 253.9138, 253.9146, 253.9153, 253.9153, 253.9153, 
    253.9154, 253.915, 253.9155, 253.9156, 253.9154, 253.9166, 253.9162, 
    253.9166, 253.9164, 253.9107, 253.911, 253.9108, 253.9111, 253.9109, 
    253.9118, 253.912, 253.9133, 253.9128, 253.9136, 253.9129, 253.913, 
    253.9136, 253.9129, 253.9145, 253.9134, 253.9155, 253.9144, 253.9155, 
    253.9153, 253.9156, 253.916, 253.9164, 253.9171, 253.9169, 253.9175, 
    253.9114, 253.9117, 253.9117, 253.9121, 253.9124, 253.913, 253.914, 
    253.9136, 253.9143, 253.9144, 253.9134, 253.914, 253.912, 253.9123, 
    253.9121, 253.9114, 253.9137, 253.9125, 253.9147, 253.9141, 253.9159, 
    253.915, 253.9168, 253.9175, 253.9183, 253.9191, 253.912, 253.9117, 
    253.9122, 253.9128, 253.9133, 253.9141, 253.9142, 253.9143, 253.9147, 
    253.915, 253.9144, 253.9151, 253.9124, 253.9138, 253.9116, 253.9123, 
    253.9127, 253.9125, 253.9136, 253.9138, 253.9148, 253.9143, 253.9174, 
    253.916, 253.9198, 253.9187, 253.9116, 253.912, 253.9131, 253.9126, 
    253.9142, 253.9145, 253.9149, 253.9153, 253.9153, 253.9155, 253.9152, 
    253.9155, 253.9141, 253.9147, 253.913, 253.9134, 253.9132, 253.913, 
    253.9137, 253.9144, 253.9144, 253.9146, 253.9152, 253.9142, 253.9175, 
    253.9154, 253.9123, 253.9129, 253.9131, 253.9128, 253.9145, 253.9139, 
    253.9155, 253.9151, 253.9158, 253.9155, 253.9154, 253.9149, 253.9147, 
    253.9139, 253.9133, 253.9129, 253.913, 253.9135, 253.9144, 253.9153, 
    253.9151, 253.9158, 253.914, 253.9148, 253.9145, 253.9152, 253.9136, 
    253.9149, 253.9133, 253.9134, 253.9139, 253.9148, 253.915, 253.9152, 
    253.9151, 253.9144, 253.9143, 253.9139, 253.9137, 253.9134, 253.9131, 
    253.9134, 253.9136, 253.9144, 253.9152, 253.916, 253.9162, 253.917, 
    253.9163, 253.9175, 253.9164, 253.9183, 253.915, 253.9164, 253.9139, 
    253.9142, 253.9147, 253.9158, 253.9152, 253.9159, 253.9143, 253.9135, 
    253.9133, 253.9129, 253.9133, 253.9133, 253.9137, 253.9135, 253.9145, 
    253.914, 253.9154, 253.9159, 253.9174, 253.9183, 253.9193, 253.9197, 
    253.9198, 253.9199 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1456411, 0.1456402, 0.1456404, 0.1456397, 0.1456401, 0.1456396, 
    0.1456409, 0.1456402, 0.1456406, 0.145641, 0.1456385, 0.1456397, 
    0.1456373, 0.145638, 0.1456362, 0.1456374, 0.145636, 0.1456362, 
    0.1456355, 0.1456357, 0.1456349, 0.1456354, 0.1456345, 0.145635, 
    0.1456349, 0.1456355, 0.1456394, 0.1456386, 0.1456395, 0.1456393, 
    0.1456394, 0.1456401, 0.1456404, 0.1456411, 0.145641, 0.1456405, 
    0.1456393, 0.1456397, 0.1456387, 0.1456387, 0.1456377, 0.1456382, 
    0.1456365, 0.145637, 0.1456357, 0.145636, 0.1456357, 0.1456358, 
    0.1456357, 0.1456362, 0.145636, 0.1456364, 0.1456381, 0.1456376, 
    0.1456391, 0.1456402, 0.1456409, 0.1456414, 0.1456413, 0.1456412, 
    0.1456405, 0.1456398, 0.1456393, 0.145639, 0.1456387, 0.1456379, 
    0.1456374, 0.1456364, 0.1456366, 0.1456363, 0.145636, 0.1456356, 
    0.1456357, 0.1456355, 0.1456363, 0.1456358, 0.1456367, 0.1456364, 
    0.1456387, 0.1456396, 0.14564, 0.1456403, 0.1456412, 0.1456406, 
    0.1456409, 0.1456403, 0.1456399, 0.1456401, 0.145639, 0.1456394, 
    0.1456374, 0.1456382, 0.1456361, 0.1456365, 0.145636, 0.1456362, 
    0.1456358, 0.1456362, 0.1456354, 0.1456353, 0.1456354, 0.145635, 
    0.1456362, 0.1456357, 0.1456401, 0.1456401, 0.1456399, 0.1456405, 
    0.1456406, 0.1456411, 0.1456406, 0.1456404, 0.1456399, 0.1456396, 
    0.1456393, 0.1456387, 0.145638, 0.1456372, 0.1456365, 0.1456361, 
    0.1456364, 0.1456362, 0.1456364, 0.1456365, 0.1456353, 0.145636, 
    0.145635, 0.1456351, 0.1456355, 0.1456351, 0.1456401, 0.1456402, 
    0.1456408, 0.1456403, 0.1456412, 0.1456407, 0.1456404, 0.1456394, 
    0.1456392, 0.145639, 0.1456386, 0.1456381, 0.1456373, 0.1456366, 
    0.145636, 0.1456361, 0.1456361, 0.1456359, 0.1456362, 0.1456359, 
    0.1456358, 0.145636, 0.1456351, 0.1456353, 0.1456351, 0.1456352, 
    0.1456402, 0.1456399, 0.14564, 0.1456397, 0.14564, 0.1456391, 0.1456388, 
    0.1456377, 0.1456381, 0.1456374, 0.1456381, 0.145638, 0.1456374, 
    0.145638, 0.1456366, 0.1456376, 0.1456359, 0.1456368, 0.1456359, 
    0.145636, 0.1456358, 0.1456355, 0.1456353, 0.1456348, 0.1456349, 
    0.1456345, 0.1456395, 0.1456391, 0.1456392, 0.1456388, 0.1456385, 
    0.145638, 0.1456371, 0.1456374, 0.1456369, 0.1456368, 0.1456376, 
    0.1456371, 0.1456389, 0.1456386, 0.1456388, 0.1456394, 0.1456374, 
    0.1456384, 0.1456365, 0.1456371, 0.1456356, 0.1456363, 0.1456349, 
    0.1456345, 0.145634, 0.1456336, 0.1456389, 0.1456392, 0.1456387, 
    0.1456382, 0.1456377, 0.145637, 0.145637, 0.1456368, 0.1456365, 
    0.1456363, 0.1456368, 0.1456362, 0.1456385, 0.1456373, 0.1456393, 
    0.1456386, 0.1456382, 0.1456384, 0.1456375, 0.1456373, 0.1456364, 
    0.1456369, 0.1456346, 0.1456355, 0.1456332, 0.1456338, 0.1456393, 
    0.1456389, 0.1456379, 0.1456384, 0.145637, 0.1456366, 0.1456364, 
    0.1456361, 0.145636, 0.1456358, 0.1456361, 0.1456359, 0.145637, 
    0.1456365, 0.145638, 0.1456376, 0.1456378, 0.145638, 0.1456374, 
    0.1456368, 0.1456368, 0.1456366, 0.1456361, 0.145637, 0.1456345, 
    0.1456359, 0.1456386, 0.145638, 0.1456379, 0.1456382, 0.1456367, 
    0.1456372, 0.1456358, 0.1456362, 0.1456356, 0.1456359, 0.1456359, 
    0.1456363, 0.1456365, 0.1456372, 0.1456377, 0.1456381, 0.145638, 
    0.1456376, 0.1456368, 0.145636, 0.1456362, 0.1456357, 0.1456371, 
    0.1456365, 0.1456367, 0.1456361, 0.1456374, 0.1456363, 0.1456378, 
    0.1456376, 0.1456372, 0.1456364, 0.1456362, 0.1456361, 0.1456362, 
    0.1456367, 0.1456368, 0.1456372, 0.1456373, 0.1456376, 0.1456379, 
    0.1456377, 0.1456374, 0.1456367, 0.1456361, 0.1456355, 0.1456354, 
    0.1456348, 0.1456353, 0.1456345, 0.1456351, 0.145634, 0.1456362, 
    0.1456352, 0.1456372, 0.145637, 0.1456365, 0.1456356, 0.1456361, 
    0.1456356, 0.1456368, 0.1456375, 0.1456377, 0.1456381, 0.1456377, 
    0.1456378, 0.1456374, 0.1456375, 0.1456367, 0.1456371, 0.1456359, 
    0.1456356, 0.1456345, 0.145634, 0.1456335, 0.1456333, 0.1456332, 0.1456332,
  0.1512731, 0.1512778, 0.1512769, 0.1512807, 0.1512786, 0.1512811, 
    0.1512741, 0.151278, 0.1512755, 0.1512736, 0.151288, 0.1512809, 
    0.1512957, 0.1512911, 0.1513027, 0.1512949, 0.1513043, 0.1513026, 
    0.1513081, 0.1513065, 0.1513134, 0.1513088, 0.1513171, 0.1513123, 
    0.1513131, 0.1513086, 0.1512824, 0.151287, 0.1512821, 0.1512827, 
    0.1512825, 0.1512786, 0.1512767, 0.1512728, 0.1512735, 0.1512764, 
    0.1512831, 0.1512808, 0.1512866, 0.1512865, 0.1512928, 0.1512899, 
    0.1513007, 0.1512977, 0.1513066, 0.1513043, 0.1513065, 0.1513058, 
    0.1513065, 0.1513031, 0.1513046, 0.1513017, 0.1512904, 0.1512937, 
    0.151284, 0.151278, 0.1512742, 0.1512715, 0.1512719, 0.1512726, 
    0.1512764, 0.15128, 0.1512828, 0.1512846, 0.1512864, 0.1512917, 
    0.1512947, 0.1513013, 0.1513001, 0.1513021, 0.1513041, 0.1513073, 
    0.1513068, 0.1513082, 0.1513021, 0.1513061, 0.1512995, 0.1513013, 
    0.1512866, 0.1512814, 0.151279, 0.1512771, 0.1512722, 0.1512756, 
    0.1512742, 0.1512775, 0.1512795, 0.1512785, 0.1512847, 0.1512823, 
    0.1512949, 0.1512894, 0.1513039, 0.1513004, 0.1513047, 0.1513025, 
    0.1513062, 0.1513029, 0.1513087, 0.15131, 0.1513091, 0.1513125, 
    0.1513027, 0.1513064, 0.1512784, 0.1512786, 0.1512794, 0.151276, 
    0.1512758, 0.1512728, 0.1512755, 0.1512766, 0.1512796, 0.1512813, 
    0.151283, 0.1512866, 0.1512907, 0.1512964, 0.1513006, 0.1513034, 
    0.1513017, 0.1513032, 0.1513015, 0.1513007, 0.1513095, 0.1513046, 
    0.1513121, 0.1513117, 0.1513082, 0.1513117, 0.1512787, 0.1512778, 
    0.1512745, 0.1512771, 0.1512724, 0.151275, 0.1512765, 0.1512822, 
    0.1512836, 0.1512847, 0.1512871, 0.1512901, 0.1512953, 0.1512999, 
    0.1513042, 0.1513039, 0.151304, 0.1513049, 0.1513026, 0.1513053, 
    0.1513058, 0.1513046, 0.1513116, 0.1513096, 0.1513116, 0.1513103, 
    0.1512781, 0.1512797, 0.1512788, 0.1512804, 0.1512793, 0.1512842, 
    0.1512858, 0.1512928, 0.15129, 0.1512946, 0.1512905, 0.1512912, 
    0.1512946, 0.1512907, 0.1512996, 0.1512935, 0.151305, 0.1512987, 
    0.1513054, 0.1513042, 0.1513062, 0.1513079, 0.1513101, 0.1513142, 
    0.1513133, 0.1513168, 0.151282, 0.151284, 0.1512839, 0.1512861, 
    0.1512876, 0.1512911, 0.1512967, 0.1512946, 0.1512984, 0.1512992, 
    0.1512934, 0.1512969, 0.1512854, 0.1512872, 0.1512862, 0.1512821, 
    0.151295, 0.1512884, 0.1513007, 0.1512971, 0.1513076, 0.1513023, 
    0.1513128, 0.1513171, 0.1513215, 0.1513264, 0.1512852, 0.1512838, 
    0.1512863, 0.1512897, 0.151293, 0.1512973, 0.1512978, 0.1512986, 
    0.1513007, 0.1513024, 0.1512988, 0.1513029, 0.1512875, 0.1512956, 
    0.1512832, 0.1512869, 0.1512895, 0.1512884, 0.1512944, 0.1512958, 
    0.1513014, 0.1512985, 0.151316, 0.1513082, 0.1513303, 0.151324, 
    0.1512833, 0.1512852, 0.1512917, 0.1512886, 0.1512976, 0.1512998, 
    0.1513016, 0.1513039, 0.1513042, 0.1513055, 0.1513033, 0.1513055, 
    0.1512973, 0.1513009, 0.151291, 0.1512934, 0.1512923, 0.1512911, 
    0.1512949, 0.1512988, 0.151299, 0.1513002, 0.1513036, 0.1512976, 
    0.1513169, 0.1513048, 0.1512873, 0.1512908, 0.1512914, 0.15129, 
    0.1512996, 0.1512961, 0.1513055, 0.151303, 0.1513072, 0.1513051, 
    0.1513048, 0.1513021, 0.1513004, 0.1512962, 0.1512929, 0.1512902, 
    0.1512908, 0.1512937, 0.1512991, 0.1513042, 0.151303, 0.1513069, 
    0.1512969, 0.151301, 0.1512994, 0.1513036, 0.1512945, 0.151302, 
    0.1512926, 0.1512934, 0.151296, 0.1513012, 0.1513025, 0.1513038, 
    0.151303, 0.1512992, 0.1512986, 0.151296, 0.1512952, 0.1512932, 
    0.1512915, 0.1512931, 0.1512946, 0.1512993, 0.1513034, 0.1513079, 
    0.1513091, 0.1513142, 0.1513099, 0.1513169, 0.1513108, 0.1513215, 
    0.1513026, 0.1513108, 0.1512962, 0.1512978, 0.1513005, 0.1513071, 
    0.1513036, 0.1513077, 0.1512986, 0.1512938, 0.1512927, 0.1512904, 
    0.1512927, 0.1512925, 0.1512948, 0.1512941, 0.1512994, 0.1512965, 
    0.1513047, 0.1513077, 0.1513164, 0.1513217, 0.1513272, 0.1513296, 
    0.1513304, 0.1513307,
  0.1611241, 0.1611301, 0.1611289, 0.1611337, 0.1611311, 0.1611342, 
    0.1611253, 0.1611303, 0.1611271, 0.1611246, 0.161143, 0.1611339, 
    0.1611529, 0.161147, 0.1611619, 0.1611519, 0.161164, 0.1611618, 
    0.1611688, 0.1611668, 0.1611757, 0.1611697, 0.1611805, 0.1611743, 
    0.1611752, 0.1611695, 0.1611359, 0.1611418, 0.1611355, 0.1611363, 
    0.161136, 0.1611311, 0.1611286, 0.1611236, 0.1611246, 0.1611282, 
    0.1611367, 0.1611339, 0.1611412, 0.1611411, 0.1611492, 0.1611455, 
    0.1611593, 0.1611554, 0.1611669, 0.161164, 0.1611667, 0.1611659, 
    0.1611667, 0.1611625, 0.1611643, 0.1611606, 0.1611462, 0.1611504, 
    0.1611379, 0.1611303, 0.1611255, 0.1611221, 0.1611225, 0.1611235, 
    0.1611283, 0.1611329, 0.1611364, 0.1611387, 0.161141, 0.1611478, 
    0.1611516, 0.1611601, 0.1611586, 0.1611611, 0.1611637, 0.1611678, 
    0.1611671, 0.161169, 0.1611611, 0.1611663, 0.1611578, 0.1611601, 
    0.1611413, 0.1611347, 0.1611316, 0.1611291, 0.1611229, 0.1611272, 
    0.1611255, 0.1611296, 0.1611321, 0.1611309, 0.1611388, 0.1611357, 
    0.1611519, 0.1611449, 0.1611634, 0.1611589, 0.1611645, 0.1611616, 
    0.1611664, 0.1611621, 0.1611697, 0.1611713, 0.1611702, 0.1611746, 
    0.1611619, 0.1611667, 0.1611308, 0.161131, 0.161132, 0.1611277, 
    0.1611275, 0.1611236, 0.1611271, 0.1611285, 0.1611323, 0.1611345, 
    0.1611366, 0.1611413, 0.1611465, 0.1611538, 0.1611592, 0.1611628, 
    0.1611606, 0.1611626, 0.1611604, 0.1611594, 0.1611706, 0.1611643, 
    0.1611739, 0.1611734, 0.161169, 0.1611734, 0.1611312, 0.16113, 0.1611258, 
    0.1611291, 0.1611232, 0.1611265, 0.1611283, 0.1611357, 0.1611374, 
    0.1611389, 0.1611419, 0.1611457, 0.1611524, 0.1611583, 0.1611638, 
    0.1611634, 0.1611636, 0.1611648, 0.1611618, 0.1611653, 0.1611658, 
    0.1611643, 0.1611733, 0.1611708, 0.1611734, 0.1611717, 0.1611304, 
    0.1611324, 0.1611313, 0.1611333, 0.1611319, 0.1611383, 0.1611402, 
    0.1611492, 0.1611456, 0.1611515, 0.1611462, 0.1611471, 0.1611516, 
    0.1611465, 0.1611579, 0.1611501, 0.1611648, 0.1611568, 0.1611653, 
    0.1611638, 0.1611663, 0.1611686, 0.1611715, 0.1611767, 0.1611755, 
    0.16118, 0.1611354, 0.161138, 0.1611378, 0.1611406, 0.1611426, 0.161147, 
    0.1611541, 0.1611515, 0.1611564, 0.1611574, 0.1611499, 0.1611544, 
    0.1611398, 0.1611421, 0.1611407, 0.1611356, 0.161152, 0.1611435, 
    0.1611593, 0.1611547, 0.1611682, 0.1611614, 0.1611748, 0.1611805, 
    0.1611861, 0.1611924, 0.1611395, 0.1611377, 0.1611409, 0.1611452, 
    0.1611494, 0.1611549, 0.1611555, 0.1611566, 0.1611593, 0.1611615, 
    0.1611568, 0.1611621, 0.1611425, 0.1611528, 0.161137, 0.1611416, 
    0.161145, 0.1611436, 0.1611512, 0.161153, 0.1611602, 0.1611565, 0.161179, 
    0.161169, 0.1611974, 0.1611893, 0.1611371, 0.1611395, 0.1611478, 
    0.1611438, 0.1611553, 0.1611582, 0.1611605, 0.1611634, 0.1611638, 
    0.1611655, 0.1611627, 0.1611654, 0.161155, 0.1611596, 0.1611469, 
    0.1611499, 0.1611486, 0.161147, 0.1611518, 0.1611569, 0.1611571, 
    0.1611587, 0.161163, 0.1611554, 0.1611801, 0.1611646, 0.1611421, 
    0.1611466, 0.1611474, 0.1611456, 0.1611579, 0.1611534, 0.1611655, 
    0.1611622, 0.1611676, 0.1611649, 0.1611645, 0.1611611, 0.161159, 
    0.1611536, 0.1611492, 0.1611459, 0.1611467, 0.1611504, 0.1611572, 
    0.1611638, 0.1611623, 0.1611672, 0.1611545, 0.1611598, 0.1611577, 
    0.1611631, 0.1611514, 0.1611611, 0.1611489, 0.16115, 0.1611533, 0.16116, 
    0.1611617, 0.1611633, 0.1611623, 0.1611574, 0.1611566, 0.1611533, 
    0.1611523, 0.1611497, 0.1611476, 0.1611495, 0.1611515, 0.1611574, 
    0.1611627, 0.1611686, 0.1611701, 0.1611767, 0.1611712, 0.1611802, 
    0.1611723, 0.1611861, 0.1611618, 0.1611723, 0.1611535, 0.1611555, 
    0.1611591, 0.1611676, 0.1611631, 0.1611684, 0.1611566, 0.1611505, 
    0.161149, 0.1611461, 0.1611491, 0.1611488, 0.1611517, 0.1611508, 
    0.1611577, 0.161154, 0.1611645, 0.1611684, 0.1611795, 0.1611863, 
    0.1611934, 0.1611966, 0.1611975, 0.1611979,
  0.175334, 0.1753385, 0.1753377, 0.1753413, 0.1753393, 0.1753417, 0.175335, 
    0.1753387, 0.1753363, 0.1753345, 0.1753483, 0.1753415, 0.1753558, 
    0.1753513, 0.1753628, 0.1753551, 0.1753644, 0.1753627, 0.1753681, 
    0.1753666, 0.1753735, 0.1753689, 0.1753772, 0.1753724, 0.1753731, 
    0.1753687, 0.1753429, 0.1753474, 0.1753426, 0.1753433, 0.175343, 
    0.1753393, 0.1753374, 0.1753338, 0.1753344, 0.1753372, 0.1753436, 
    0.1753414, 0.175347, 0.1753468, 0.175353, 0.1753502, 0.1753608, 
    0.1753578, 0.1753667, 0.1753644, 0.1753665, 0.1753659, 0.1753665, 
    0.1753632, 0.1753646, 0.1753618, 0.1753507, 0.1753539, 0.1753444, 
    0.1753387, 0.1753351, 0.1753326, 0.1753329, 0.1753336, 0.1753372, 
    0.1753407, 0.1753433, 0.1753451, 0.1753468, 0.175352, 0.1753549, 
    0.1753614, 0.1753603, 0.1753622, 0.1753642, 0.1753674, 0.1753669, 
    0.1753683, 0.1753622, 0.1753662, 0.1753596, 0.1753614, 0.175347, 
    0.175342, 0.1753397, 0.1753378, 0.1753332, 0.1753364, 0.1753351, 
    0.1753382, 0.1753401, 0.1753392, 0.1753451, 0.1753428, 0.1753551, 
    0.1753497, 0.1753639, 0.1753605, 0.1753648, 0.1753626, 0.1753663, 
    0.175363, 0.1753688, 0.1753701, 0.1753692, 0.1753726, 0.1753628, 
    0.1753665, 0.1753391, 0.1753393, 0.17534, 0.1753368, 0.1753366, 
    0.1753337, 0.1753363, 0.1753374, 0.1753403, 0.1753419, 0.1753435, 
    0.175347, 0.1753509, 0.1753566, 0.1753607, 0.1753635, 0.1753618, 
    0.1753633, 0.1753616, 0.1753609, 0.1753696, 0.1753646, 0.1753721, 
    0.1753717, 0.1753683, 0.1753718, 0.1753394, 0.1753385, 0.1753354, 
    0.1753378, 0.1753334, 0.1753358, 0.1753372, 0.1753428, 0.1753441, 
    0.1753452, 0.1753475, 0.1753504, 0.1753555, 0.1753601, 0.1753643, 
    0.175364, 0.1753641, 0.175365, 0.1753627, 0.1753654, 0.1753658, 
    0.1753647, 0.1753717, 0.1753697, 0.1753717, 0.1753704, 0.1753388, 
    0.1753403, 0.1753395, 0.175341, 0.1753399, 0.1753447, 0.1753462, 
    0.1753531, 0.1753503, 0.1753548, 0.1753508, 0.1753515, 0.1753549, 
    0.175351, 0.1753597, 0.1753537, 0.1753651, 0.1753588, 0.1753654, 
    0.1753643, 0.1753662, 0.175368, 0.1753702, 0.1753743, 0.1753734, 
    0.1753769, 0.1753426, 0.1753445, 0.1753444, 0.1753465, 0.175348, 
    0.1753514, 0.1753568, 0.1753548, 0.1753586, 0.1753593, 0.1753536, 
    0.175357, 0.1753459, 0.1753476, 0.1753466, 0.1753427, 0.1753552, 
    0.1753487, 0.1753608, 0.1753572, 0.1753677, 0.1753624, 0.1753728, 
    0.1753773, 0.1753817, 0.1753867, 0.1753456, 0.1753443, 0.1753467, 
    0.17535, 0.1753532, 0.1753574, 0.1753579, 0.1753587, 0.1753608, 
    0.1753625, 0.1753589, 0.175363, 0.1753479, 0.1753558, 0.1753438, 
    0.1753473, 0.1753498, 0.1753488, 0.1753546, 0.1753559, 0.1753615, 
    0.1753586, 0.1753761, 0.1753683, 0.1753906, 0.1753842, 0.1753438, 
    0.1753456, 0.175352, 0.175349, 0.1753577, 0.1753599, 0.1753617, 0.175364, 
    0.1753643, 0.1753656, 0.1753634, 0.1753656, 0.1753574, 0.1753611, 
    0.1753513, 0.1753536, 0.1753526, 0.1753514, 0.175355, 0.1753589, 
    0.1753591, 0.1753603, 0.1753637, 0.1753578, 0.175377, 0.1753649, 
    0.1753476, 0.1753511, 0.1753516, 0.1753503, 0.1753597, 0.1753563, 
    0.1753656, 0.1753631, 0.1753672, 0.1753651, 0.1753648, 0.1753622, 
    0.1753605, 0.1753564, 0.1753531, 0.1753505, 0.1753511, 0.1753539, 
    0.1753592, 0.1753643, 0.1753631, 0.1753669, 0.1753571, 0.1753611, 
    0.1753595, 0.1753637, 0.1753547, 0.1753621, 0.1753528, 0.1753536, 
    0.1753562, 0.1753614, 0.1753626, 0.1753639, 0.1753631, 0.1753593, 
    0.1753587, 0.1753561, 0.1753554, 0.1753535, 0.1753518, 0.1753533, 
    0.1753548, 0.1753594, 0.1753635, 0.175368, 0.1753691, 0.1753743, 0.17537, 
    0.1753771, 0.1753709, 0.1753817, 0.1753627, 0.1753709, 0.1753563, 
    0.1753579, 0.1753606, 0.1753672, 0.1753637, 0.1753678, 0.1753587, 
    0.175354, 0.1753529, 0.1753507, 0.1753529, 0.1753528, 0.1753549, 
    0.1753542, 0.1753595, 0.1753567, 0.1753648, 0.1753678, 0.1753765, 
    0.1753818, 0.1753875, 0.17539, 0.1753907, 0.175391,
  0.1899463, 0.1899477, 0.1899474, 0.1899485, 0.1899479, 0.1899486, 
    0.1899466, 0.1899477, 0.189947, 0.1899464, 0.1899507, 0.1899486, 
    0.1899532, 0.1899517, 0.1899556, 0.189953, 0.1899561, 0.1899555, 
    0.1899574, 0.1899568, 0.1899593, 0.1899576, 0.1899606, 0.1899589, 
    0.1899591, 0.1899576, 0.189949, 0.1899505, 0.1899489, 0.1899491, 
    0.1899491, 0.1899479, 0.1899473, 0.1899462, 0.1899464, 0.1899472, 
    0.1899492, 0.1899486, 0.1899503, 0.1899503, 0.1899523, 0.1899514, 
    0.1899549, 0.1899539, 0.1899569, 0.1899561, 0.1899568, 0.1899566, 
    0.1899568, 0.1899557, 0.1899562, 0.1899552, 0.1899515, 0.1899526, 
    0.1899495, 0.1899477, 0.1899466, 0.1899458, 0.189946, 0.1899462, 
    0.1899472, 0.1899483, 0.1899492, 0.1899497, 0.1899503, 0.1899519, 
    0.1899529, 0.1899551, 0.1899547, 0.1899554, 0.189956, 0.1899571, 
    0.1899569, 0.1899574, 0.1899554, 0.1899567, 0.1899545, 0.1899551, 
    0.1899503, 0.1899488, 0.189948, 0.1899475, 0.189946, 0.189947, 0.1899466, 
    0.1899476, 0.1899482, 0.1899479, 0.1899497, 0.189949, 0.189953, 
    0.1899512, 0.1899559, 0.1899548, 0.1899562, 0.1899555, 0.1899568, 
    0.1899556, 0.1899576, 0.1899581, 0.1899578, 0.189959, 0.1899555, 
    0.1899568, 0.1899479, 0.1899479, 0.1899481, 0.1899471, 0.1899471, 
    0.1899462, 0.189947, 0.1899473, 0.1899482, 0.1899487, 0.1899492, 
    0.1899503, 0.1899516, 0.1899535, 0.1899548, 0.1899558, 0.1899552, 
    0.1899557, 0.1899552, 0.1899549, 0.1899579, 0.1899562, 0.1899588, 
    0.1899586, 0.1899574, 0.1899587, 0.1899479, 0.1899477, 0.1899467, 
    0.1899475, 0.1899461, 0.1899468, 0.1899473, 0.189949, 0.1899494, 
    0.1899498, 0.1899505, 0.1899514, 0.1899531, 0.1899546, 0.1899561, 
    0.189956, 0.189956, 0.1899563, 0.1899555, 0.1899564, 0.1899566, 
    0.1899562, 0.1899586, 0.1899579, 0.1899586, 0.1899582, 0.1899478, 
    0.1899482, 0.189948, 0.1899484, 0.1899481, 0.1899496, 0.1899501, 
    0.1899523, 0.1899514, 0.1899529, 0.1899515, 0.1899518, 0.1899529, 
    0.1899516, 0.1899545, 0.1899525, 0.1899563, 0.1899542, 0.1899565, 
    0.1899561, 0.1899567, 0.1899573, 0.1899581, 0.1899596, 0.1899592, 
    0.1899605, 0.1899489, 0.1899495, 0.1899495, 0.1899502, 0.1899506, 
    0.1899517, 0.1899535, 0.1899529, 0.1899541, 0.1899544, 0.1899525, 
    0.1899536, 0.18995, 0.1899505, 0.1899502, 0.189949, 0.189953, 0.1899509, 
    0.1899549, 0.1899537, 0.1899572, 0.1899554, 0.189959, 0.1899606, 
    0.1899622, 0.189964, 0.1899499, 0.1899495, 0.1899502, 0.1899513, 
    0.1899523, 0.1899537, 0.1899539, 0.1899542, 0.1899549, 0.1899555, 
    0.1899542, 0.1899556, 0.1899506, 0.1899532, 0.1899493, 0.1899504, 
    0.1899512, 0.1899509, 0.1899528, 0.1899532, 0.1899551, 0.1899541, 
    0.1899602, 0.1899574, 0.1899655, 0.1899631, 0.1899493, 0.1899499, 
    0.1899519, 0.189951, 0.1899538, 0.1899546, 0.1899552, 0.1899559, 
    0.1899561, 0.1899565, 0.1899558, 0.1899565, 0.1899537, 0.189955, 
    0.1899517, 0.1899525, 0.1899521, 0.1899517, 0.189953, 0.1899542, 
    0.1899543, 0.1899547, 0.1899558, 0.1899539, 0.1899605, 0.1899563, 
    0.1899505, 0.1899516, 0.1899518, 0.1899514, 0.1899545, 0.1899533, 
    0.1899565, 0.1899556, 0.1899571, 0.1899564, 0.1899562, 0.1899554, 
    0.1899548, 0.1899534, 0.1899523, 0.1899515, 0.1899517, 0.1899526, 
    0.1899543, 0.1899561, 0.1899557, 0.189957, 0.1899536, 0.189955, 
    0.1899544, 0.1899559, 0.1899528, 0.1899553, 0.1899522, 0.1899525, 
    0.1899533, 0.1899551, 0.1899555, 0.1899559, 0.1899557, 0.1899544, 
    0.1899542, 0.1899533, 0.1899531, 0.1899524, 0.1899519, 0.1899524, 
    0.1899529, 0.1899544, 0.1899558, 0.1899573, 0.1899577, 0.1899596, 
    0.189958, 0.1899605, 0.1899583, 0.1899622, 0.1899555, 0.1899583, 
    0.1899534, 0.1899539, 0.1899548, 0.1899571, 0.1899559, 0.1899573, 
    0.1899542, 0.1899526, 0.1899522, 0.1899515, 0.1899523, 0.1899522, 
    0.1899529, 0.1899527, 0.1899544, 0.1899535, 0.1899562, 0.1899573, 
    0.1899603, 0.1899623, 0.1899643, 0.1899652, 0.1899655, 0.1899657,
  0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973189, 0.1973189, 0.197319, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973188, 0.1973188, 
    0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 
    0.1973188, 0.1973188, 0.1973189, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973188, 0.1973189, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 
    0.1973189, 0.197319, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.197319, 0.1973191, 0.1973192, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.197319, 0.1973189, 0.1973192, 0.1973191, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.197319, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973189, 0.197319, 0.1973189, 0.1973191, 
    0.1973188, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973189, 0.1973189, 0.197319, 0.1973191, 0.1973192, 0.1973192, 
    0.1973192, 0.1973193,
  0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 
    0.1984797, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 
    0.1984799, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984798, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984796, 
    0.1984796, 0.1984796,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  5.611711, 5.611763, 5.611753, 5.611795, 5.611772, 5.611799, 5.611722, 
    5.611765, 5.611738, 5.611716, 5.611874, 5.611797, 5.611958, 5.611908, 
    5.612037, 5.61195, 5.612055, 5.612035, 5.612096, 5.612079, 5.612154, 
    5.612104, 5.612195, 5.612143, 5.612151, 5.612103, 5.611814, 5.611864, 
    5.61181, 5.611817, 5.611814, 5.611773, 5.61175, 5.611707, 5.611715, 
    5.611747, 5.611821, 5.611797, 5.61186, 5.611858, 5.611928, 5.611896, 
    5.612014, 5.61198, 5.61208, 5.612055, 5.612079, 5.612072, 5.612079, 
    5.612041, 5.612058, 5.612025, 5.611902, 5.611937, 5.611831, 5.611764, 
    5.611723, 5.611693, 5.611698, 5.611705, 5.611747, 5.611788, 5.611818, 
    5.611838, 5.611858, 5.611915, 5.611948, 5.61202, 5.612008, 5.61203, 
    5.612052, 5.612088, 5.612082, 5.612098, 5.61203, 5.612075, 5.612, 
    5.612021, 5.611859, 5.611804, 5.611776, 5.611755, 5.611701, 5.611738, 
    5.611723, 5.611759, 5.611782, 5.611771, 5.611839, 5.611812, 5.611949, 
    5.611891, 5.61205, 5.61201, 5.612059, 5.612035, 5.612076, 5.612039, 
    5.612104, 5.612117, 5.612108, 5.612145, 5.612037, 5.612078, 5.61177, 
    5.611772, 5.611781, 5.611742, 5.611741, 5.611707, 5.611737, 5.61175, 
    5.611783, 5.611802, 5.61182, 5.61186, 5.611904, 5.611967, 5.612013, 
    5.612045, 5.612026, 5.612042, 5.612023, 5.612015, 5.612112, 5.612057, 
    5.61214, 5.612136, 5.612098, 5.612136, 5.611773, 5.611763, 5.611726, 
    5.611755, 5.611703, 5.611732, 5.611748, 5.611812, 5.611827, 5.611839, 
    5.611866, 5.611898, 5.611955, 5.612005, 5.612054, 5.61205, 5.612051, 
    5.612062, 5.612036, 5.612066, 5.612071, 5.612058, 5.612135, 5.612113, 
    5.612135, 5.612122, 5.611766, 5.611784, 5.611774, 5.611792, 5.611779, 
    5.611834, 5.61185, 5.611928, 5.611897, 5.611947, 5.611902, 5.61191, 
    5.611947, 5.611905, 5.612001, 5.611934, 5.612062, 5.61199, 5.612067, 
    5.612053, 5.612075, 5.612094, 5.612119, 5.612164, 5.612154, 5.612191, 
    5.61181, 5.611832, 5.611831, 5.611854, 5.611871, 5.611909, 5.611969, 
    5.611947, 5.611989, 5.611997, 5.611934, 5.611971, 5.611847, 5.611866, 
    5.611856, 5.611811, 5.611951, 5.611879, 5.612013, 5.611974, 5.612092, 
    5.612032, 5.612148, 5.612195, 5.612242, 5.612293, 5.611845, 5.61183, 
    5.611857, 5.611894, 5.611929, 5.611976, 5.611981, 5.611989, 5.612013, 
    5.612034, 5.611991, 5.612039, 5.611869, 5.611958, 5.611823, 5.611863, 
    5.611892, 5.61188, 5.611944, 5.611959, 5.612021, 5.611989, 5.612182, 
    5.612097, 5.612335, 5.612268, 5.611824, 5.611845, 5.611916, 5.611882, 
    5.611979, 5.612003, 5.612025, 5.61205, 5.612053, 5.612068, 5.612044, 
    5.612068, 5.611976, 5.612017, 5.611908, 5.611934, 5.611922, 5.611909, 
    5.61195, 5.611992, 5.611994, 5.612008, 5.612045, 5.61198, 5.612191, 
    5.612059, 5.611867, 5.611905, 5.611912, 5.611897, 5.612, 5.611963, 
    5.612068, 5.61204, 5.612086, 5.612063, 5.61206, 5.61203, 5.612011, 
    5.611965, 5.611928, 5.611899, 5.611906, 5.611938, 5.611995, 5.612053, 
    5.61204, 5.612083, 5.611972, 5.612018, 5.611999, 5.612047, 5.611946, 
    5.612028, 5.611925, 5.611934, 5.611962, 5.61202, 5.612035, 5.612049, 
    5.612041, 5.611996, 5.61199, 5.611962, 5.611953, 5.611932, 5.611914, 
    5.61193, 5.611947, 5.611997, 5.612044, 5.612094, 5.612107, 5.612163, 
    5.612116, 5.612191, 5.612125, 5.612241, 5.612035, 5.612125, 5.611964, 
    5.611981, 5.612011, 5.612085, 5.612047, 5.612092, 5.61199, 5.611938, 
    5.611926, 5.611901, 5.611927, 5.611925, 5.611949, 5.611941, 5.611999, 
    5.611968, 5.612059, 5.612092, 5.612186, 5.612243, 5.612302, 5.612328, 
    5.612336, 5.612339 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  5.912984e-15, 5.911852e-15, 5.912067e-15, 5.911167e-15, 5.911658e-15, 
    5.911075e-15, 5.912745e-15, 5.911816e-15, 5.912403e-15, 5.912869e-15, 
    5.909452e-15, 5.911124e-15, 5.907629e-15, 5.908707e-15, 5.905975e-15, 
    5.907809e-15, 5.905602e-15, 5.906006e-15, 5.904738e-15, 5.9051e-15, 
    5.903526e-15, 5.904571e-15, 5.902678e-15, 5.903764e-15, 5.903602e-15, 
    5.904609e-15, 5.910767e-15, 5.909667e-15, 5.910837e-15, 5.910679e-15, 
    5.910745e-15, 5.911656e-15, 5.912129e-15, 5.913056e-15, 5.912884e-15, 
    5.912195e-15, 5.910607e-15, 5.911132e-15, 5.90977e-15, 5.9098e-15, 
    5.908301e-15, 5.908977e-15, 5.906447e-15, 5.90716e-15, 5.905085e-15, 
    5.905609e-15, 5.905113e-15, 5.90526e-15, 5.905111e-15, 5.905878e-15, 
    5.905551e-15, 5.90622e-15, 5.908855e-15, 5.908086e-15, 5.910392e-15, 
    5.911814e-15, 5.912708e-15, 5.913359e-15, 5.913267e-15, 5.913096e-15, 
    5.912191e-15, 5.911324e-15, 5.910669e-15, 5.910235e-15, 5.909805e-15, 
    5.908559e-15, 5.907854e-15, 5.906313e-15, 5.906572e-15, 5.906119e-15, 
    5.90566e-15, 5.904915e-15, 5.905035e-15, 5.904711e-15, 5.906118e-15, 
    5.905189e-15, 5.906726e-15, 5.906307e-15, 5.90976e-15, 5.910987e-15, 
    5.911571e-15, 5.912029e-15, 5.913198e-15, 5.912394e-15, 5.912713e-15, 
    5.91194e-15, 5.91146e-15, 5.911695e-15, 5.910223e-15, 5.910797e-15, 
    5.907813e-15, 5.909096e-15, 5.905714e-15, 5.906518e-15, 5.905518e-15, 
    5.906024e-15, 5.905163e-15, 5.905938e-15, 5.904585e-15, 5.904299e-15, 
    5.904496e-15, 5.903715e-15, 5.905983e-15, 5.905119e-15, 5.911704e-15, 
    5.911667e-15, 5.911482e-15, 5.912295e-15, 5.912341e-15, 5.913064e-15, 
    5.912414e-15, 5.912143e-15, 5.911426e-15, 5.911017e-15, 5.910623e-15, 
    5.909756e-15, 5.908802e-15, 5.907449e-15, 5.906466e-15, 5.905813e-15, 
    5.906209e-15, 5.90586e-15, 5.906253e-15, 5.906434e-15, 5.904411e-15, 
    5.905552e-15, 5.903828e-15, 5.90392e-15, 5.904706e-15, 5.90391e-15, 
    5.911639e-15, 5.911859e-15, 5.912646e-15, 5.91203e-15, 5.913143e-15, 
    5.912528e-15, 5.912181e-15, 5.910801e-15, 5.910481e-15, 5.910207e-15, 
    5.909649e-15, 5.908943e-15, 5.90771e-15, 5.906627e-15, 5.90563e-15, 
    5.905702e-15, 5.905677e-15, 5.905462e-15, 5.906005e-15, 5.905373e-15, 
    5.905274e-15, 5.905543e-15, 5.903934e-15, 5.904392e-15, 5.903923e-15, 
    5.904219e-15, 5.911785e-15, 5.911412e-15, 5.911615e-15, 5.911238e-15, 
    5.911509e-15, 5.910324e-15, 5.909969e-15, 5.90829e-15, 5.908961e-15, 
    5.907874e-15, 5.908845e-15, 5.908677e-15, 5.907869e-15, 5.908787e-15, 
    5.9067e-15, 5.908142e-15, 5.905454e-15, 5.906919e-15, 5.905364e-15, 
    5.905635e-15, 5.90518e-15, 5.90478e-15, 5.904264e-15, 5.903335e-15, 
    5.903547e-15, 5.902759e-15, 5.91085e-15, 5.910373e-15, 5.910402e-15, 
    5.909894e-15, 5.909521e-15, 5.908698e-15, 5.907395e-15, 5.90788e-15, 
    5.906975e-15, 5.906798e-15, 5.908165e-15, 5.907339e-15, 5.910044e-15, 
    5.909621e-15, 5.909863e-15, 5.91082e-15, 5.907787e-15, 5.90935e-15, 
    5.906453e-15, 5.907295e-15, 5.904839e-15, 5.906072e-15, 5.903667e-15, 
    5.902677e-15, 5.901684e-15, 5.900598e-15, 5.910099e-15, 5.910424e-15, 
    5.909829e-15, 5.909033e-15, 5.908256e-15, 5.907247e-15, 5.907136e-15, 
    5.906951e-15, 5.906454e-15, 5.906045e-15, 5.906905e-15, 5.905941e-15, 
    5.909549e-15, 5.907646e-15, 5.910559e-15, 5.909699e-15, 5.909074e-15, 
    5.909334e-15, 5.907932e-15, 5.907607e-15, 5.906291e-15, 5.906964e-15, 
    5.902932e-15, 5.904714e-15, 5.899729e-15, 5.901127e-15, 5.91054e-15, 
    5.910093e-15, 5.908558e-15, 5.909286e-15, 5.907172e-15, 5.906658e-15, 
    5.906229e-15, 5.905704e-15, 5.905637e-15, 5.905325e-15, 5.905839e-15, 
    5.90534e-15, 5.907244e-15, 5.90639e-15, 5.908717e-15, 5.908158e-15, 
    5.908411e-15, 5.908698e-15, 5.907813e-15, 5.906896e-15, 5.906854e-15, 
    5.906563e-15, 5.905784e-15, 5.907163e-15, 5.902743e-15, 5.905505e-15, 
    5.909607e-15, 5.908776e-15, 5.908632e-15, 5.908958e-15, 5.906711e-15, 
    5.907527e-15, 5.905329e-15, 5.905917e-15, 5.904948e-15, 5.905432e-15, 
    5.905504e-15, 5.90612e-15, 5.90651e-15, 5.907494e-15, 5.908288e-15, 
    5.908908e-15, 5.908762e-15, 5.908081e-15, 5.906834e-15, 5.905641e-15, 
    5.905905e-15, 5.905022e-15, 5.907326e-15, 5.906369e-15, 5.906746e-15, 
    5.905761e-15, 5.907898e-15, 5.906143e-15, 5.908355e-15, 5.908156e-15, 
    5.907543e-15, 5.906319e-15, 5.906016e-15, 5.905733e-15, 5.905903e-15, 
    5.906798e-15, 5.906935e-15, 5.907553e-15, 5.907734e-15, 5.908198e-15, 
    5.908592e-15, 5.908237e-15, 5.907869e-15, 5.906789e-15, 5.905829e-15, 
    5.904778e-15, 5.904512e-15, 5.90334e-15, 5.904323e-15, 5.902731e-15, 
    5.904128e-15, 5.901689e-15, 5.906009e-15, 5.904127e-15, 5.907508e-15, 
    5.907137e-15, 5.90649e-15, 5.904965e-15, 5.905765e-15, 5.904819e-15, 
    5.906939e-15, 5.908068e-15, 5.908333e-15, 5.908874e-15, 5.908321e-15, 
    5.908365e-15, 5.907838e-15, 5.908007e-15, 5.906753e-15, 5.907425e-15, 
    5.905511e-15, 5.904821e-15, 5.902849e-15, 5.901658e-15, 5.900413e-15, 
    5.899875e-15, 5.89971e-15, 5.899642e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  7.064673, 7.091394, 7.086197, 7.107788, 7.095809, 7.109952, 7.07009, 
    7.092452, 7.078174, 7.067084, 7.149392, 7.108754, 7.191628, 7.1657, 
    7.230989, 7.18758, 7.23977, 7.22975, 7.259978, 7.251309, 7.290048, 
    7.263982, 7.310216, 7.283824, 7.287942, 7.263121, 7.117015, 7.144345, 
    7.115375, 7.119316, 7.11755, 7.096052, 7.085228, 7.062644, 7.066742, 
    7.083337, 7.121089, 7.108265, 7.140369, 7.139648, 7.175253, 7.159182, 
    7.219244, 7.202137, 7.251671, 7.239187, 7.251081, 7.247475, 7.251129, 
    7.232827, 7.240663, 7.224579, 7.162187, 7.180475, 7.126032, 7.092965, 
    7.071068, 7.055552, 7.057744, 7.061921, 7.083434, 7.103719, 7.119205, 
    7.129473, 7.139545, 7.170063, 7.186289, 7.2227, 7.216131, 7.227273, 
    7.237947, 7.255877, 7.252925, 7.260831, 7.226987, 7.249462, 7.212389, 
    7.222512, 7.142235, 7.111725, 7.098618, 7.087194, 7.059428, 7.078591, 
    7.071031, 7.089037, 7.100491, 7.094826, 7.129752, 7.116222, 7.187251, 
    7.156634, 7.236701, 7.21748, 7.241315, 7.229147, 7.250002, 7.231231, 
    7.263779, 7.270875, 7.266024, 7.284689, 7.230191, 7.251077, 7.094665, 
    7.095588, 7.099896, 7.080974, 7.07982, 7.062529, 7.077917, 7.084474, 
    7.101158, 7.111033, 7.120434, 7.140852, 7.163658, 7.195657, 7.218724, 
    7.234216, 7.224717, 7.233102, 7.223727, 7.219338, 7.268212, 7.240733, 
    7.282002, 7.279716, 7.261017, 7.279973, 7.096237, 7.090923, 7.072484, 
    7.086911, 7.060648, 7.075334, 7.083786, 7.116497, 7.123699, 7.130273, 
    7.143284, 7.160004, 7.189404, 7.21507, 7.23857, 7.236847, 7.237453, 
    7.242705, 7.229694, 7.244843, 7.247383, 7.240736, 7.279409, 7.268345, 
    7.279667, 7.272462, 7.092652, 7.101599, 7.096762, 7.105856, 7.099445, 
    7.127896, 7.136333, 7.175931, 7.159672, 7.185576, 7.162303, 7.16642, 
    7.186401, 7.163563, 7.213644, 7.179642, 7.242909, 7.208827, 7.245048, 
    7.238468, 7.24937, 7.259139, 7.271452, 7.2942, 7.28893, 7.307993, 
    7.114957, 7.126531, 7.125532, 7.137533, 7.146417, 7.165713, 7.196737, 
    7.185061, 7.206518, 7.210828, 7.178241, 7.198226, 7.134208, 7.144511, 
    7.138382, 7.11587, 7.187738, 7.150835, 7.219104, 7.199028, 7.257744, 
    7.228487, 7.286027, 7.310709, 7.334038, 7.361323, 7.132795, 7.125009, 
    7.138964, 7.15829, 7.176286, 7.200249, 7.20271, 7.207205, 7.218869, 
    7.228683, 7.208618, 7.231146, 7.146883, 7.190952, 7.122044, 7.142735, 
    7.157154, 7.150836, 7.183731, 7.191497, 7.223123, 7.206766, 7.304603, 
    7.26119, 7.38218, 7.34821, 7.122276, 7.132773, 7.169347, 7.151928, 
    7.201857, 7.214184, 7.224225, 7.237062, 7.238455, 7.246072, 7.233593, 
    7.245582, 7.200301, 7.22051, 7.165171, 7.178604, 7.172424, 7.165645, 
    7.186584, 7.20893, 7.209424, 7.216599, 7.236819, 7.20206, 7.310193, 
    7.24324, 7.144219, 7.164455, 7.167368, 7.159518, 7.212946, 7.19355, 
    7.245888, 7.231717, 7.254951, 7.243397, 7.241698, 7.226885, 7.217671, 
    7.194435, 7.175577, 7.160658, 7.164126, 7.180522, 7.210303, 7.238575, 
    7.232373, 7.253184, 7.198227, 7.221224, 7.212324, 7.235551, 7.184748, 
    7.227947, 7.173734, 7.178477, 7.193165, 7.222775, 7.229362, 7.236372, 
    7.232049, 7.211063, 7.207636, 7.192811, 7.188715, 7.177445, 7.168118, 
    7.176636, 7.185586, 7.211078, 7.234103, 7.259275, 7.265452, 7.294931, 
    7.270906, 7.310564, 7.276806, 7.335334, 7.230479, 7.275845, 7.193839, 
    7.202643, 7.218572, 7.25524, 7.235442, 7.258607, 7.207503, 7.181081, 
    7.174275, 7.161562, 7.174566, 7.173509, 7.185968, 7.181963, 7.211926, 
    7.19582, 7.241651, 7.258429, 7.305988, 7.335251, 7.365155, 7.378378, 
    7.382408, 7.384092 ;

 WIND =
  5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  0.0002557225, 0.0002556716, 0.0002556813, 0.0002556407, 0.0002556629, 
    0.0002556366, 0.0002557118, 0.0002556699, 0.0002556964, 0.0002557174, 
    0.0002555633, 0.0002556388, 0.0002554814, 0.00025553, 0.0002554069, 
    0.0002554895, 0.0002553901, 0.0002554084, 0.0002553513, 0.0002553676, 
    0.0002552965, 0.0002553437, 0.0002552582, 0.0002553073, 0.0002552999, 
    0.0002553455, 0.0002556227, 0.000255573, 0.0002556259, 0.0002556187, 
    0.0002556217, 0.0002556627, 0.000255684, 0.0002557258, 0.000255718, 
    0.000255687, 0.0002556155, 0.0002556391, 0.0002555778, 0.0002555792, 
    0.0002555117, 0.0002555421, 0.0002554283, 0.0002554604, 0.0002553669, 
    0.0002553905, 0.0002553682, 0.0002553748, 0.0002553681, 0.0002554027, 
    0.0002553879, 0.0002554181, 0.0002555366, 0.000255502, 0.0002556058, 
    0.0002556698, 0.0002557101, 0.0002557394, 0.0002557353, 0.0002557276, 
    0.0002556868, 0.0002556478, 0.0002556183, 0.0002555988, 0.0002555794, 
    0.0002555232, 0.0002554915, 0.0002554222, 0.0002554339, 0.0002554135, 
    0.0002553928, 0.0002553592, 0.0002553646, 0.00025535, 0.0002554134, 
    0.0002553716, 0.0002554408, 0.0002554219, 0.0002555772, 0.0002556326, 
    0.0002556588, 0.0002556795, 0.0002557322, 0.000255696, 0.0002557103, 
    0.0002556755, 0.0002556539, 0.0002556645, 0.0002555983, 0.0002556241, 
    0.0002554897, 0.0002555475, 0.0002553952, 0.0002554315, 0.0002553864, 
    0.0002554092, 0.0002553704, 0.0002554053, 0.0002553443, 0.0002553314, 
    0.0002553403, 0.0002553051, 0.0002554074, 0.0002553684, 0.0002556649, 
    0.0002556632, 0.0002556549, 0.0002556915, 0.0002556935, 0.0002557262, 
    0.0002556969, 0.0002556846, 0.0002556524, 0.000255634, 0.0002556162, 
    0.0002555772, 0.0002555342, 0.0002554733, 0.0002554292, 0.0002553997, 
    0.0002554176, 0.0002554018, 0.0002554195, 0.0002554277, 0.0002553365, 
    0.0002553879, 0.0002553102, 0.0002553144, 0.0002553498, 0.0002553139, 
    0.000255662, 0.0002556719, 0.0002557073, 0.0002556796, 0.0002557297, 
    0.000255702, 0.0002556863, 0.0002556242, 0.0002556099, 0.0002555975, 
    0.0002555724, 0.0002555406, 0.0002554851, 0.0002554363, 0.0002553915, 
    0.0002553947, 0.0002553936, 0.0002553839, 0.0002554083, 0.0002553799, 
    0.0002553754, 0.0002553876, 0.000255315, 0.0002553356, 0.0002553145, 
    0.0002553279, 0.0002556686, 0.0002556518, 0.0002556609, 0.0002556439, 
    0.0002556561, 0.0002556027, 0.0002555867, 0.0002555112, 0.0002555414, 
    0.0002554925, 0.0002555362, 0.0002555286, 0.0002554921, 0.0002555336, 
    0.0002554396, 0.0002555044, 0.0002553835, 0.0002554494, 0.0002553795, 
    0.0002553917, 0.0002553712, 0.0002553531, 0.0002553299, 0.0002552879, 
    0.0002552975, 0.0002552619, 0.0002556265, 0.000255605, 0.0002556063, 
    0.0002555834, 0.0002555666, 0.0002555296, 0.0002554709, 0.0002554928, 
    0.000255452, 0.000255444, 0.0002555056, 0.0002554683, 0.0002555902, 
    0.000255571, 0.000255582, 0.0002556251, 0.0002554885, 0.0002555589, 
    0.0002554285, 0.0002554664, 0.0002553558, 0.0002554113, 0.0002553029, 
    0.0002552581, 0.0002552134, 0.0002551642, 0.0002555926, 0.0002556073, 
    0.0002555805, 0.0002555446, 0.0002555097, 0.0002554642, 0.0002554593, 
    0.0002554509, 0.0002554286, 0.0002554102, 0.0002554488, 0.0002554055, 
    0.0002555677, 0.0002554822, 0.0002556134, 0.0002555746, 0.0002555465, 
    0.0002555582, 0.0002554951, 0.0002554805, 0.0002554212, 0.0002554515, 
    0.0002552697, 0.0002553501, 0.000255125, 0.0002551881, 0.0002556125, 
    0.0002555924, 0.0002555232, 0.000255556, 0.0002554609, 0.0002554378, 
    0.0002554185, 0.0002553948, 0.0002553918, 0.0002553777, 0.0002554009, 
    0.0002553784, 0.0002554641, 0.0002554257, 0.0002555305, 0.0002555053, 
    0.0002555166, 0.0002555296, 0.0002554898, 0.0002554484, 0.0002554466, 
    0.0002554335, 0.0002553982, 0.0002554605, 0.000255261, 0.0002553857, 
    0.0002555705, 0.0002555331, 0.0002555266, 0.0002555413, 0.0002554401, 
    0.0002554769, 0.0002553779, 0.0002554044, 0.0002553607, 0.0002553825, 
    0.0002553858, 0.0002554136, 0.0002554311, 0.0002554753, 0.0002555111, 
    0.000255539, 0.0002555325, 0.0002555018, 0.0002554456, 0.0002553919, 
    0.0002554038, 0.0002553641, 0.0002554678, 0.0002554248, 0.0002554417, 
    0.0002553973, 0.0002554936, 0.0002554144, 0.0002555141, 0.0002555052, 
    0.0002554776, 0.0002554224, 0.0002554089, 0.0002553961, 0.0002554038, 
    0.000255444, 0.0002554502, 0.000255478, 0.0002554861, 0.0002555071, 
    0.0002555249, 0.0002555088, 0.0002554922, 0.0002554437, 0.0002554004, 
    0.000255353, 0.0002553411, 0.000255288, 0.0002553324, 0.0002552605, 
    0.0002553236, 0.0002552135, 0.0002554085, 0.0002553236, 0.000255476, 
    0.0002554593, 0.0002554302, 0.0002553614, 0.0002553976, 0.0002553549, 
    0.0002554504, 0.0002555012, 0.0002555132, 0.0002555375, 0.0002555126, 
    0.0002555146, 0.0002554909, 0.0002554985, 0.000255442, 0.0002554723, 
    0.0002553861, 0.0002553549, 0.000255266, 0.0002552121, 0.0002551559, 
    0.0002551316, 0.0002551241, 0.000255121 ;

 W_SCALAR =
  0.6261148, 0.627772, 0.62745, 0.6287856, 0.6280448, 0.6289191, 0.6264508, 
    0.6278378, 0.6269525, 0.626264, 0.6313739, 0.6288451, 0.6339946, 
    0.6323858, 0.6364231, 0.6337445, 0.6369624, 0.6363456, 0.6382005, 
    0.6376694, 0.6400391, 0.6384455, 0.6412655, 0.6396586, 0.6399102, 
    0.6383929, 0.6293542, 0.6310594, 0.6292531, 0.6294965, 0.6293873, 
    0.6280602, 0.627391, 0.6259879, 0.6262427, 0.6272731, 0.6296058, 
    0.6288143, 0.6308079, 0.6307629, 0.6329789, 0.6319802, 0.6356989, 
    0.6346431, 0.6376916, 0.6369256, 0.6376556, 0.6374343, 0.6376585, 
    0.636535, 0.6370165, 0.6360273, 0.6321673, 0.633303, 0.629913, 0.6278706, 
    0.6265118, 0.6255469, 0.6256833, 0.6259434, 0.6272792, 0.6285336, 
    0.6294889, 0.6301275, 0.6307564, 0.6326588, 0.633664, 0.6359124, 
    0.6355067, 0.6361938, 0.6368494, 0.6379496, 0.6377686, 0.6382532, 
    0.6361755, 0.6375567, 0.6352757, 0.6359, 0.630928, 0.6290279, 0.62822, 
    0.6275119, 0.6257882, 0.6269789, 0.6265096, 0.6276255, 0.6283342, 
    0.6279837, 0.630145, 0.6293051, 0.6337236, 0.6318223, 0.6367729, 0.63559, 
    0.6370563, 0.6363083, 0.6375897, 0.6364365, 0.6384333, 0.6388679, 
    0.638571, 0.6397107, 0.6363725, 0.6376557, 0.6279739, 0.6280311, 
    0.6282973, 0.6271266, 0.6270549, 0.625981, 0.6269366, 0.6273434, 
    0.6283752, 0.6289852, 0.6295649, 0.6308383, 0.6322592, 0.6342434, 
    0.6356667, 0.63662, 0.6360355, 0.6365516, 0.6359747, 0.6357042, 
    0.6387051, 0.637021, 0.6395468, 0.6394072, 0.6382647, 0.6394229, 
    0.6280712, 0.6277422, 0.6265996, 0.6274939, 0.625864, 0.6267766, 
    0.6273012, 0.6293229, 0.6297665, 0.6301779, 0.6309899, 0.6320313, 
    0.6338563, 0.6354419, 0.6368875, 0.6367816, 0.6368189, 0.6371417, 
    0.636342, 0.6372729, 0.6374292, 0.6370207, 0.6393885, 0.6387125, 
    0.6394042, 0.6389641, 0.6278492, 0.6284026, 0.6281036, 0.6286659, 
    0.6282698, 0.6300302, 0.6305575, 0.6330219, 0.6320109, 0.6336194, 
    0.6321743, 0.6324306, 0.6336721, 0.6322524, 0.6353546, 0.6332525, 
    0.6371542, 0.6350583, 0.6372855, 0.6368812, 0.6375504, 0.6381494, 
    0.6389025, 0.640291, 0.6399696, 0.6411298, 0.6292272, 0.6299443, 
    0.629881, 0.630631, 0.6311855, 0.6323861, 0.6343096, 0.6335866, 
    0.6349136, 0.6351798, 0.6331637, 0.6344021, 0.6304239, 0.6310676, 
    0.6306843, 0.6292838, 0.6337535, 0.6314616, 0.6356903, 0.6344512, 
    0.6380641, 0.6362687, 0.6397927, 0.6412964, 0.6427092, 0.6443588, 
    0.6303353, 0.6298483, 0.6307201, 0.6319257, 0.6330429, 0.6345268, 
    0.6346784, 0.6349562, 0.6356754, 0.6362798, 0.6350442, 0.6364312, 
    0.6312171, 0.6339521, 0.6296642, 0.6309571, 0.6318546, 0.6314608, 
    0.6335039, 0.633985, 0.6359382, 0.6349289, 0.6409255, 0.6382761, 
    0.6456128, 0.6435673, 0.6296781, 0.6303336, 0.6326126, 0.6315288, 
    0.6346257, 0.6353869, 0.6360052, 0.6367954, 0.6368806, 0.6373485, 
    0.6365817, 0.6373182, 0.6345299, 0.6357767, 0.6323522, 0.6331866, 
    0.6328028, 0.6323817, 0.6336808, 0.6350636, 0.635093, 0.6355361, 
    0.6367843, 0.6346382, 0.6412675, 0.6371781, 0.631048, 0.6323094, 
    0.6324891, 0.6320008, 0.6353106, 0.6341124, 0.6373371, 0.6364663, 
    0.6378927, 0.6371841, 0.6370798, 0.6361691, 0.6356018, 0.6341674, 
    0.632999, 0.6320716, 0.6322873, 0.6333058, 0.6351482, 0.6368884, 
    0.6365075, 0.6377843, 0.6344014, 0.6358212, 0.6352727, 0.6367022, 
    0.6335675, 0.6362381, 0.632884, 0.6331784, 0.6340886, 0.6359175, 
    0.6363215, 0.6367531, 0.6364867, 0.6351948, 0.634983, 0.6340664, 
    0.6338133, 0.6331143, 0.6325353, 0.6330644, 0.6336197, 0.6351953, 
    0.6366136, 0.638158, 0.6385356, 0.6403375, 0.6388711, 0.6412902, 
    0.6392343, 0.6427908, 0.6363924, 0.6391734, 0.6341299, 0.6346742, 
    0.6356583, 0.6379119, 0.6366956, 0.6381178, 0.6349747, 0.633341, 
    0.6329178, 0.6321281, 0.6329358, 0.6328701, 0.6336426, 0.6333944, 
    0.6352476, 0.6342525, 0.6370773, 0.6381066, 0.6410084, 0.6427839, 
    0.6445881, 0.6453838, 0.6456259, 0.6457272,
  0.5467909, 0.548835, 0.5484377, 0.5500853, 0.5491714, 0.5502501, 0.5472054, 
    0.5489162, 0.5478241, 0.5469749, 0.5532789, 0.5501587, 0.5565134, 
    0.5545277, 0.5595115, 0.5562047, 0.5601775, 0.5594159, 0.5617064, 
    0.5610505, 0.5639775, 0.5620091, 0.5654924, 0.5635074, 0.5638182, 
    0.5619441, 0.5507868, 0.5528908, 0.5506622, 0.5509623, 0.5508276, 
    0.5491904, 0.5483649, 0.5466344, 0.5469487, 0.5482196, 0.5510973, 
    0.5501208, 0.5525804, 0.5525249, 0.5552596, 0.5540271, 0.5586174, 
    0.5573139, 0.5610779, 0.5601321, 0.5610335, 0.5607602, 0.5610371, 
    0.5596497, 0.5602443, 0.5590229, 0.554258, 0.5556598, 0.5514762, 
    0.5489565, 0.5472805, 0.5460905, 0.5462587, 0.5465795, 0.548227, 
    0.5497745, 0.550953, 0.5517409, 0.5525169, 0.5548645, 0.5561054, 
    0.558881, 0.5583802, 0.5592284, 0.560038, 0.5613967, 0.5611731, 
    0.5617715, 0.5592058, 0.5609115, 0.5580949, 0.5588657, 0.5527286, 
    0.5503842, 0.5493875, 0.5485141, 0.5463881, 0.5478566, 0.5472779, 
    0.5486543, 0.5495284, 0.549096, 0.5517624, 0.5507263, 0.5561789, 
    0.5538322, 0.5599436, 0.558483, 0.5602934, 0.5593698, 0.5609521, 
    0.5595281, 0.5619941, 0.5625306, 0.562164, 0.5635718, 0.5594491, 
    0.5610336, 0.549084, 0.5491545, 0.5494829, 0.5480388, 0.5479504, 
    0.5466259, 0.5478045, 0.5483062, 0.549579, 0.5503316, 0.5510467, 
    0.552618, 0.5543715, 0.5568205, 0.5585777, 0.5597547, 0.559033, 
    0.5596702, 0.5589579, 0.558624, 0.5623296, 0.5602499, 0.5633693, 
    0.5631968, 0.5617857, 0.5632163, 0.549204, 0.5487982, 0.5473888, 
    0.5484918, 0.5464815, 0.5476072, 0.5482541, 0.5507481, 0.5512955, 
    0.5518031, 0.552805, 0.5540902, 0.5563427, 0.5583001, 0.560085, 
    0.5599543, 0.5600003, 0.5603989, 0.5594115, 0.5605609, 0.5607539, 
    0.5602496, 0.5631738, 0.5623388, 0.5631932, 0.5626496, 0.5489301, 
    0.5496128, 0.5492439, 0.5499375, 0.549449, 0.5516208, 0.5522714, 
    0.5553128, 0.554065, 0.5560502, 0.5542667, 0.5545829, 0.5561153, 
    0.5543631, 0.5581924, 0.5555974, 0.5604144, 0.5578266, 0.5605764, 
    0.5600773, 0.5609036, 0.5616434, 0.5625735, 0.5642887, 0.5638916, 
    0.5653248, 0.5506301, 0.5515149, 0.5514368, 0.5523622, 0.5530463, 
    0.5545281, 0.5569023, 0.5560098, 0.5576478, 0.5579765, 0.5554878, 
    0.5570164, 0.5521066, 0.5529009, 0.5524279, 0.5506999, 0.5562158, 
    0.5533872, 0.5586067, 0.5570769, 0.561538, 0.559321, 0.563673, 0.5655306, 
    0.5672763, 0.5693149, 0.5519974, 0.5513964, 0.5524722, 0.5539598, 
    0.5553386, 0.5571703, 0.5573575, 0.5577005, 0.5585884, 0.5593346, 
    0.5578091, 0.5595216, 0.5530853, 0.556461, 0.5511693, 0.5527645, 
    0.5538721, 0.5533862, 0.5559078, 0.5565016, 0.5589129, 0.5576667, 
    0.5650725, 0.5617998, 0.5708649, 0.5683366, 0.5511864, 0.5519952, 
    0.5548077, 0.55347, 0.5572925, 0.5582322, 0.5589957, 0.5599713, 
    0.5600765, 0.5606543, 0.5597074, 0.5606169, 0.5571742, 0.5587134, 
    0.5544862, 0.5555161, 0.5550423, 0.5545226, 0.5561261, 0.5578331, 
    0.5578694, 0.5584164, 0.5599575, 0.5573079, 0.5654948, 0.5604437, 
    0.5528768, 0.5544333, 0.5546553, 0.5540525, 0.558138, 0.5566588, 
    0.5606402, 0.5595649, 0.5613263, 0.5604513, 0.5603225, 0.559198, 
    0.5584975, 0.5567267, 0.5552845, 0.55414, 0.5544061, 0.5556632, 
    0.5579374, 0.5600861, 0.5596157, 0.5611925, 0.5570156, 0.5587683, 
    0.5580912, 0.5598563, 0.5559862, 0.5592831, 0.5551426, 0.5555059, 
    0.5566294, 0.5588874, 0.5593861, 0.559919, 0.5595902, 0.5579951, 
    0.5577335, 0.5566021, 0.5562897, 0.5554268, 0.5547122, 0.5553652, 
    0.5560507, 0.5579957, 0.5597468, 0.561654, 0.5621203, 0.564346, 
    0.5625347, 0.565523, 0.5629832, 0.567377, 0.5594736, 0.562908, 0.5566804, 
    0.5573523, 0.5585672, 0.56135, 0.559848, 0.5616044, 0.5577233, 0.5557066, 
    0.5551842, 0.5542096, 0.5552065, 0.5551254, 0.5560789, 0.5557725, 
    0.5580602, 0.5568317, 0.5603194, 0.5615904, 0.5651748, 0.5673686, 
    0.5695983, 0.5705819, 0.5708812, 0.5710062,
  0.5141823, 0.5164323, 0.515995, 0.5178089, 0.5168027, 0.5179903, 0.5146385, 
    0.5165216, 0.5153195, 0.5143847, 0.521326, 0.5178897, 0.52489, 0.5227019, 
    0.5281949, 0.5245497, 0.5289292, 0.5280896, 0.5306154, 0.529892, 
    0.5331206, 0.5309492, 0.5347923, 0.5326021, 0.532945, 0.5308776, 
    0.5185813, 0.5208985, 0.5184441, 0.5187746, 0.5186262, 0.5168235, 
    0.5159149, 0.5140101, 0.514356, 0.5157548, 0.5189232, 0.5178479, 
    0.5205567, 0.5204955, 0.5235084, 0.5221503, 0.5272092, 0.5257723, 
    0.5299222, 0.5288792, 0.5298733, 0.5295719, 0.5298772, 0.5283473, 
    0.5290029, 0.5276563, 0.5224048, 0.5239493, 0.5193405, 0.516566, 
    0.5147212, 0.5134115, 0.5135967, 0.5139497, 0.515763, 0.5174666, 
    0.5187643, 0.519632, 0.5204868, 0.523073, 0.5244403, 0.5274998, 
    0.5269477, 0.5278828, 0.5287754, 0.5302737, 0.5300272, 0.5306872, 
    0.5278579, 0.5297386, 0.5266332, 0.5274829, 0.5207199, 0.518138, 
    0.5170406, 0.5160791, 0.513739, 0.5153552, 0.5147182, 0.5162333, 
    0.5171957, 0.5167197, 0.5196558, 0.5185147, 0.5245213, 0.5219356, 
    0.5286713, 0.527061, 0.5290571, 0.5280387, 0.5297835, 0.5282132, 
    0.5309327, 0.5315245, 0.5311201, 0.5326731, 0.5281262, 0.5298734, 
    0.5167064, 0.5167841, 0.5171456, 0.5155559, 0.5154586, 0.5140007, 
    0.5152978, 0.5158501, 0.5172514, 0.5180801, 0.5188676, 0.5205981, 
    0.5225298, 0.5252284, 0.5271654, 0.5284631, 0.5276674, 0.5283699, 
    0.5275846, 0.5272164, 0.5313028, 0.5290091, 0.5324497, 0.5322595, 
    0.5307029, 0.5322809, 0.5168386, 0.5163918, 0.5148403, 0.5160546, 
    0.5138418, 0.5150807, 0.5157929, 0.5185387, 0.5191414, 0.5197005, 
    0.5208041, 0.5222199, 0.5247018, 0.5268593, 0.5288273, 0.5286831, 
    0.5287339, 0.5291734, 0.5280847, 0.5293521, 0.5295649, 0.5290087, 
    0.532234, 0.5313129, 0.5322554, 0.5316557, 0.516537, 0.5172886, 
    0.5168825, 0.5176462, 0.5171083, 0.5194997, 0.5202163, 0.5235668, 
    0.5221921, 0.5243795, 0.5224143, 0.5227627, 0.5244512, 0.5225205, 
    0.5267406, 0.5238805, 0.5291905, 0.5263373, 0.5293692, 0.5288188, 
    0.52973, 0.5305459, 0.5315718, 0.533464, 0.5330259, 0.5346074, 0.5184087, 
    0.5193831, 0.5192971, 0.5203164, 0.5210699, 0.5227023, 0.5253186, 
    0.524335, 0.5261403, 0.5265027, 0.5237598, 0.5254443, 0.5200348, 
    0.5209097, 0.5203887, 0.5184857, 0.5245619, 0.5214453, 0.5271974, 
    0.5255111, 0.5304296, 0.5279849, 0.5327848, 0.5348344, 0.5367613, 
    0.539012, 0.5199145, 0.5192527, 0.5204375, 0.5220762, 0.5235954, 
    0.525614, 0.5258204, 0.5261984, 0.5271772, 0.5279999, 0.5263181, 
    0.5282061, 0.5211129, 0.5248322, 0.5190026, 0.5207595, 0.5219796, 
    0.5214443, 0.5242226, 0.524877, 0.527535, 0.5261612, 0.5343289, 
    0.5307184, 0.5407239, 0.5379319, 0.5190214, 0.5199122, 0.5230103, 
    0.5215366, 0.5257487, 0.5267845, 0.5276262, 0.5287019, 0.5288179, 
    0.5294551, 0.5284109, 0.5294138, 0.5256183, 0.5273151, 0.5226561, 
    0.523791, 0.5232689, 0.5226963, 0.5244632, 0.5263446, 0.5263845, 
    0.5269876, 0.5286866, 0.5257657, 0.534795, 0.5292228, 0.5208831, 
    0.5225978, 0.5228423, 0.5221784, 0.5266807, 0.5250502, 0.5294395, 
    0.5282539, 0.5301961, 0.5292312, 0.5290892, 0.5278493, 0.527077, 
    0.5251251, 0.5235357, 0.5222747, 0.5225679, 0.523953, 0.5264596, 
    0.5288286, 0.5283098, 0.5300485, 0.5254434, 0.5273756, 0.526629, 
    0.5285751, 0.5243089, 0.527943, 0.5233794, 0.5237797, 0.5250179, 
    0.5275068, 0.5280567, 0.5286442, 0.5282816, 0.5265232, 0.5262348, 
    0.5249877, 0.5246434, 0.5236925, 0.5229052, 0.5236247, 0.52438, 
    0.5265238, 0.5284544, 0.5305575, 0.5310718, 0.5335273, 0.531529, 
    0.534826, 0.5320237, 0.5368724, 0.5281531, 0.5319408, 0.5250741, 
    0.5258147, 0.5271538, 0.5302223, 0.5285659, 0.5305029, 0.5262235, 
    0.5240009, 0.5234252, 0.5223514, 0.5234498, 0.5233604, 0.5244111, 
    0.5240735, 0.5265949, 0.5252408, 0.5290857, 0.5304875, 0.5344418, 
    0.5368631, 0.539325, 0.5404113, 0.5407418, 0.54088,
  0.507082, 0.5094726, 0.5090079, 0.5109358, 0.5098663, 0.5111287, 0.5075666, 
    0.5095676, 0.5082902, 0.5072972, 0.5146762, 0.5110217, 0.5184694, 
    0.5161402, 0.5219896, 0.5181071, 0.5227723, 0.5218774, 0.5245696, 
    0.5237985, 0.5272414, 0.5249255, 0.5290251, 0.5266883, 0.527054, 
    0.5248492, 0.5117571, 0.5142214, 0.5116111, 0.5119625, 0.5118048, 
    0.5098885, 0.5089228, 0.5068991, 0.5072665, 0.5087527, 0.5121205, 
    0.5109773, 0.5138578, 0.5137928, 0.5169986, 0.5155533, 0.5209395, 
    0.5194089, 0.5238306, 0.5227189, 0.5237784, 0.5234572, 0.5237826, 
    0.5221521, 0.5228508, 0.5214157, 0.515824, 0.5174679, 0.5125643, 
    0.5096148, 0.5076545, 0.5062633, 0.50646, 0.506835, 0.5087614, 0.510572, 
    0.5119516, 0.5128743, 0.5137834, 0.5165351, 0.5179906, 0.521249, 
    0.5206609, 0.521657, 0.5226083, 0.5242054, 0.5239425, 0.5246461, 
    0.5216306, 0.5236349, 0.5203258, 0.5212311, 0.5140314, 0.5112857, 
    0.5101191, 0.5090972, 0.5066112, 0.5083281, 0.5076514, 0.5092612, 
    0.510284, 0.5097781, 0.5128996, 0.5116862, 0.5180768, 0.5153248, 
    0.5224974, 0.5207816, 0.5229085, 0.5218232, 0.5236828, 0.5220092, 
    0.5249079, 0.525539, 0.5251077, 0.526764, 0.5219164, 0.5237786, 0.509764, 
    0.5098465, 0.5102308, 0.5085413, 0.5084379, 0.5068891, 0.5082672, 
    0.508854, 0.5103432, 0.5112241, 0.5120614, 0.5139019, 0.5159571, 
    0.5188298, 0.5208928, 0.5222754, 0.5214276, 0.5221761, 0.5213394, 
    0.5209472, 0.5253026, 0.5228573, 0.5265257, 0.5263228, 0.5246629, 
    0.5263457, 0.5099044, 0.5094296, 0.5077811, 0.5090712, 0.5067204, 
    0.5080364, 0.5087932, 0.5117117, 0.5123526, 0.5129471, 0.514121, 
    0.5156273, 0.5182691, 0.5205668, 0.5226636, 0.5225099, 0.5225641, 
    0.5230325, 0.5218722, 0.5232229, 0.5234497, 0.522857, 0.5262956, 
    0.5253134, 0.5263185, 0.5256789, 0.5095839, 0.5103828, 0.5099511, 
    0.5107629, 0.5101911, 0.5127336, 0.5134957, 0.5170608, 0.5155977, 
    0.5179259, 0.5158342, 0.5162049, 0.5180022, 0.5159472, 0.5204403, 
    0.5173947, 0.5230507, 0.5200107, 0.5232412, 0.5226545, 0.5236257, 
    0.5244955, 0.5255894, 0.5276077, 0.5271404, 0.5288278, 0.5115736, 
    0.5126095, 0.5125182, 0.5136021, 0.5144038, 0.5161406, 0.5189258, 
    0.5178785, 0.5198009, 0.5201868, 0.5172662, 0.5190597, 0.5133027, 
    0.5142333, 0.5136791, 0.5116554, 0.5181201, 0.5148032, 0.520927, 
    0.5191308, 0.5243715, 0.5217658, 0.5268831, 0.5290701, 0.531127, 
    0.5335308, 0.5131748, 0.5124709, 0.513731, 0.5154744, 0.5170912, 
    0.5192404, 0.5194601, 0.5198628, 0.5209053, 0.5217819, 0.5199902, 
    0.5220016, 0.5144494, 0.5184079, 0.5122049, 0.5140735, 0.5153716, 
    0.514802, 0.5177588, 0.5184556, 0.5212865, 0.5198231, 0.5285305, 
    0.5246794, 0.5353601, 0.532377, 0.512225, 0.5131723, 0.5164685, 
    0.5149003, 0.5193838, 0.5204871, 0.5213837, 0.52253, 0.5226536, 
    0.5233327, 0.5222199, 0.5232886, 0.519245, 0.5210522, 0.5160915, 
    0.5172994, 0.5167437, 0.5161343, 0.518015, 0.5200185, 0.520061, 
    0.5207034, 0.5225136, 0.5194019, 0.5290279, 0.5230851, 0.5142051, 
    0.5160295, 0.5162897, 0.5155831, 0.5203764, 0.51864, 0.523316, 0.5220525, 
    0.5241226, 0.5230941, 0.5229427, 0.5216213, 0.5207987, 0.5187197, 
    0.5170277, 0.5156856, 0.5159976, 0.5174718, 0.5201409, 0.5226649, 
    0.5221121, 0.5239653, 0.5190588, 0.5211167, 0.5203214, 0.5223948, 
    0.5178508, 0.5217212, 0.5168613, 0.5172874, 0.5186055, 0.5212564, 
    0.5218424, 0.5224685, 0.5220821, 0.5202087, 0.5199016, 0.5185735, 
    0.5182068, 0.5171946, 0.5163566, 0.5171223, 0.5179265, 0.5202093, 
    0.5222661, 0.5245079, 0.5250563, 0.5276752, 0.5255437, 0.5290611, 
    0.5260714, 0.5312456, 0.5219451, 0.5259829, 0.5186654, 0.5194541, 
    0.5208805, 0.5241506, 0.5223851, 0.5244496, 0.5198895, 0.5175229, 
    0.5169101, 0.5157672, 0.5169362, 0.5168411, 0.5179596, 0.5176002, 
    0.5202851, 0.518843, 0.522939, 0.5244332, 0.5286511, 0.5312357, 
    0.5338653, 0.535026, 0.5353792, 0.5355269,
  0.5310288, 0.5334982, 0.5330179, 0.5350106, 0.533905, 0.5352101, 0.5315292, 
    0.5335963, 0.5322765, 0.5312509, 0.5388809, 0.5350995, 0.5428115, 
    0.5403972, 0.5464646, 0.5424359, 0.5472774, 0.546348, 0.5491452, 
    0.5483436, 0.5519241, 0.5495152, 0.5537811, 0.5513485, 0.5517291, 
    0.5494357, 0.5358599, 0.53841, 0.535709, 0.5360725, 0.5359093, 0.5339279, 
    0.53293, 0.5308399, 0.5312192, 0.5327542, 0.5362359, 0.5350536, 
    0.5380336, 0.5379663, 0.5412867, 0.5397893, 0.5453742, 0.543786, 
    0.548377, 0.547222, 0.5483229, 0.547989, 0.5483272, 0.5466332, 0.5473589, 
    0.5458686, 0.5400698, 0.5417732, 0.536695, 0.533645, 0.5316199, 
    0.5301836, 0.5303866, 0.5307737, 0.5327632, 0.5346345, 0.5360612, 
    0.5370158, 0.5379566, 0.5408065, 0.5423151, 0.5456956, 0.5450851, 
    0.5461192, 0.5471071, 0.5487666, 0.5484933, 0.5492247, 0.5460917, 
    0.5481737, 0.5447374, 0.545677, 0.5382133, 0.5353725, 0.5341663, 
    0.5331103, 0.5305427, 0.5323157, 0.5316167, 0.5332797, 0.5343368, 
    0.5338139, 0.5370419, 0.5357866, 0.5424045, 0.5395526, 0.5469918, 
    0.5452104, 0.547419, 0.5462918, 0.5482234, 0.5464849, 0.5494968, 
    0.5501531, 0.5497046, 0.5514273, 0.5463886, 0.5483229, 0.5337992, 
    0.5338845, 0.5342818, 0.5325359, 0.5324291, 0.5308296, 0.5322527, 
    0.532859, 0.534398, 0.5353088, 0.5361747, 0.5380793, 0.5402075, 
    0.5431852, 0.5453258, 0.5467614, 0.545881, 0.5466582, 0.5457894, 
    0.5453822, 0.5499072, 0.5473658, 0.5511795, 0.5509683, 0.5492421, 
    0.5509921, 0.5339444, 0.5334537, 0.5317506, 0.5330834, 0.5306554, 
    0.5320144, 0.5327961, 0.5358131, 0.536476, 0.5370911, 0.5383061, 
    0.5398659, 0.5426038, 0.5449874, 0.5471645, 0.5470049, 0.5470611, 
    0.5475478, 0.5463426, 0.5477456, 0.5479812, 0.5473654, 0.55094, 
    0.5499184, 0.5509638, 0.5502986, 0.5336131, 0.5344389, 0.5339927, 
    0.5348319, 0.5342407, 0.5368702, 0.5376589, 0.5413513, 0.5398353, 
    0.542248, 0.5400802, 0.5404643, 0.5423271, 0.5401973, 0.5448561, 
    0.5416973, 0.5475667, 0.5444103, 0.5477645, 0.5471551, 0.5481641, 
    0.5490681, 0.5502055, 0.5523053, 0.551819, 0.5535756, 0.5356702, 
    0.5367419, 0.5366473, 0.537769, 0.5385988, 0.5403978, 0.5432849, 
    0.5421989, 0.5441927, 0.5445932, 0.5415641, 0.5434238, 0.5374591, 
    0.5384223, 0.5378487, 0.5357548, 0.5424494, 0.5390124, 0.5453612, 
    0.5434975, 0.5489392, 0.5462322, 0.5515513, 0.5538279, 0.555971, 
    0.5584781, 0.5373267, 0.5365984, 0.5379024, 0.5397075, 0.5413827, 
    0.5436112, 0.5438392, 0.5442569, 0.5453388, 0.5462488, 0.5443891, 
    0.546477, 0.5386461, 0.5427478, 0.5363232, 0.5382569, 0.539601, 
    0.5390112, 0.5420747, 0.5427972, 0.5457345, 0.5442157, 0.553266, 
    0.5492593, 0.5603875, 0.5572744, 0.536344, 0.5373241, 0.5407374, 
    0.5391129, 0.5437599, 0.5449046, 0.5458354, 0.5470257, 0.5471541, 
    0.5478596, 0.5467037, 0.5478138, 0.5436159, 0.5454913, 0.5403469, 
    0.5415985, 0.5410226, 0.5403911, 0.5423404, 0.5444184, 0.5444626, 
    0.5451292, 0.5470088, 0.5437787, 0.553784, 0.5476024, 0.5383931, 
    0.5402825, 0.5405522, 0.5398202, 0.5447899, 0.5429885, 0.5478423, 
    0.5465299, 0.5486805, 0.5476117, 0.5474545, 0.5460821, 0.5452281, 
    0.5430712, 0.5413169, 0.5399263, 0.5402496, 0.5417773, 0.5445455, 
    0.5471659, 0.5465918, 0.548517, 0.5434228, 0.5455582, 0.5447328, 
    0.5468853, 0.5421701, 0.5461859, 0.5411444, 0.5415861, 0.5429527, 
    0.5457033, 0.5463117, 0.5469618, 0.5465606, 0.5446157, 0.5442971, 
    0.5429195, 0.5425393, 0.54149, 0.5406215, 0.541415, 0.5422486, 0.5446165, 
    0.5467517, 0.549081, 0.5496511, 0.5523756, 0.550158, 0.5538185, 
    0.5507067, 0.5560948, 0.5464183, 0.5506147, 0.5430148, 0.5438328, 
    0.545313, 0.5487095, 0.5468752, 0.5490204, 0.5442846, 0.5418302, 
    0.541195, 0.5400109, 0.5412221, 0.5411236, 0.5422829, 0.5419103, 
    0.5446951, 0.543199, 0.5474506, 0.5490034, 0.5533916, 0.5560843, 
    0.558827, 0.5600387, 0.5604075, 0.5605618,
  0.535215, 0.5380583, 0.537505, 0.5398022, 0.5385273, 0.5400323, 0.5357908, 
    0.5381714, 0.5366511, 0.5354705, 0.5442734, 0.5399048, 0.5488272, 
    0.5460286, 0.5530714, 0.5483914, 0.5540173, 0.5529358, 0.5561932, 
    0.555259, 0.5594366, 0.5566247, 0.5616078, 0.5587642, 0.5592087, 
    0.5565321, 0.5407823, 0.5437287, 0.5406081, 0.5410277, 0.5408393, 
    0.5385537, 0.5374036, 0.5349978, 0.5354341, 0.5372012, 0.5412164, 
    0.5398518, 0.5432935, 0.5432156, 0.5470591, 0.5453246, 0.5518034, 
    0.5499582, 0.555298, 0.5539528, 0.5552348, 0.5548459, 0.5552399, 
    0.5532677, 0.5541123, 0.5523782, 0.5456493, 0.5476229, 0.5417466, 
    0.5382276, 0.5358952, 0.5342429, 0.5344764, 0.5349216, 0.5372116, 
    0.5393683, 0.5410146, 0.5421172, 0.5432045, 0.5465026, 0.5482513, 
    0.552177, 0.5514672, 0.5526696, 0.5538191, 0.5557519, 0.5554335, 
    0.5562859, 0.5526377, 0.5550611, 0.5510632, 0.5521553, 0.5435013, 
    0.5402197, 0.5388285, 0.5376113, 0.5346559, 0.5366962, 0.5358915, 
    0.5378065, 0.539025, 0.5384222, 0.5421473, 0.5406978, 0.548355, 
    0.5450506, 0.5536849, 0.5516129, 0.5541821, 0.5528703, 0.555119, 
    0.553095, 0.5566033, 0.5573688, 0.5568456, 0.5588562, 0.5529829, 
    0.555235, 0.5384053, 0.5385036, 0.5389616, 0.5369498, 0.5368267, 
    0.5349858, 0.5366237, 0.5373218, 0.5390956, 0.5401462, 0.5411457, 
    0.5433463, 0.5458089, 0.5492609, 0.5517471, 0.5534167, 0.5523925, 
    0.5532967, 0.5522861, 0.5518126, 0.5570819, 0.5541202, 0.5585667, 
    0.5583202, 0.5563062, 0.558348, 0.5385727, 0.538007, 0.5360457, 
    0.5375804, 0.5347855, 0.5363493, 0.5372494, 0.5407283, 0.5414937, 
    0.5422042, 0.5436085, 0.5454133, 0.5485862, 0.5513538, 0.5538859, 
    0.5537002, 0.5537656, 0.5543321, 0.5529295, 0.5545625, 0.5548369, 
    0.5541198, 0.5582872, 0.557095, 0.558315, 0.5575385, 0.5381908, 
    0.5391428, 0.5386283, 0.539596, 0.5389143, 0.5419489, 0.5428603, 
    0.5471339, 0.5453779, 0.5481735, 0.5456614, 0.5461062, 0.5482653, 
    0.545797, 0.5512012, 0.5475349, 0.5543541, 0.5506833, 0.5545846, 
    0.553875, 0.55505, 0.5561034, 0.55743, 0.559882, 0.5593137, 0.5613673, 
    0.5405633, 0.5418007, 0.5416915, 0.5429876, 0.5439471, 0.5460292, 
    0.5493765, 0.5481166, 0.5504305, 0.5508956, 0.5473805, 0.5495377, 
    0.5426294, 0.543743, 0.5430797, 0.540661, 0.5484071, 0.5444255, 
    0.5517883, 0.5496233, 0.5559531, 0.552801, 0.559001, 0.5616626, 
    0.5641724, 0.5671141, 0.5424764, 0.541635, 0.5431418, 0.54523, 0.5471703, 
    0.5497553, 0.5500199, 0.550505, 0.5517622, 0.5528204, 0.5506586, 
    0.5530857, 0.5440018, 0.5487532, 0.5413172, 0.5435517, 0.5451067, 
    0.5444241, 0.5479726, 0.5488106, 0.5522222, 0.5504572, 0.5610052, 
    0.5563263, 0.5693585, 0.5657009, 0.5413412, 0.5424734, 0.5464225, 
    0.5445418, 0.5499279, 0.5512576, 0.5523396, 0.5537243, 0.5538738, 
    0.5546952, 0.5533496, 0.554642, 0.5497608, 0.5519395, 0.5459703, 
    0.5474204, 0.546753, 0.5460215, 0.5482807, 0.5506927, 0.5507439, 
    0.5515186, 0.5537046, 0.5499498, 0.5616112, 0.5543957, 0.5437092, 
    0.5458958, 0.546208, 0.5453604, 0.5511243, 0.5490325, 0.5546752, 
    0.5531473, 0.5556517, 0.5544065, 0.5542235, 0.5526266, 0.5516335, 
    0.5491284, 0.547094, 0.5454832, 0.5458576, 0.5476277, 0.5508403, 
    0.5538875, 0.5532194, 0.5554611, 0.5495365, 0.5520173, 0.5510579, 
    0.553561, 0.5480832, 0.5527471, 0.5468942, 0.5474061, 0.548991, 0.552186, 
    0.5528935, 0.5536501, 0.5531831, 0.5509219, 0.5505518, 0.5489524, 
    0.5485114, 0.5472946, 0.5462883, 0.5472078, 0.5481742, 0.5509228, 
    0.5534055, 0.5561185, 0.5567833, 0.5599641, 0.5573745, 0.5616516, 
    0.5580149, 0.5643175, 0.5530175, 0.5579075, 0.5490631, 0.5500126, 
    0.5517322, 0.5556855, 0.5535492, 0.5560478, 0.5505372, 0.547689, 
    0.5469528, 0.5455812, 0.5469842, 0.54687, 0.548214, 0.5477819, 0.5510141, 
    0.5492768, 0.554219, 0.5560279, 0.561152, 0.5643053, 0.567524, 0.5689483, 
    0.5693821, 0.5695636,
  0.5840928, 0.5875039, 0.586839, 0.5896026, 0.5880677, 0.5898799, 0.5847825, 
    0.5876399, 0.585814, 0.5843988, 0.5950066, 0.5897262, 0.6005461, 
    0.5971375, 0.6057424, 0.6000144, 0.606905, 0.6055759, 0.6095858, 
    0.6084337, 0.6135982, 0.6101183, 0.6162958, 0.6127648, 0.6133156, 
    0.610004, 0.5907843, 0.5943465, 0.5905741, 0.5910804, 0.5908531, 
    0.5880995, 0.5867173, 0.5838327, 0.5843552, 0.5864743, 0.5913082, 
    0.5896623, 0.5938194, 0.5937251, 0.598391, 0.5962822, 0.6041865, 
    0.6019276, 0.6084818, 0.6068256, 0.6084039, 0.6079248, 0.6084102, 
    0.6059834, 0.6070218, 0.6048915, 0.5966766, 0.5990776, 0.5919484, 
    0.5877073, 0.5849076, 0.5829297, 0.5832089, 0.5837415, 0.5864867, 
    0.58908, 0.5910646, 0.5923963, 0.5937116, 0.5977138, 0.5998436, 
    0.6046446, 0.6037745, 0.605249, 0.6066612, 0.6090413, 0.6086487, 
    0.6097001, 0.6052099, 0.6081898, 0.6032797, 0.6046181, 0.594071, 
    0.5901058, 0.5884302, 0.5869668, 0.5834237, 0.5858681, 0.5849032, 
    0.5872012, 0.5886666, 0.5879413, 0.5924328, 0.5906823, 0.59997, 
    0.5959496, 0.6064963, 0.603953, 0.6071077, 0.6054955, 0.6082612, 
    0.6057714, 0.6100919, 0.6110377, 0.6103912, 0.6128787, 0.6056337, 
    0.608404, 0.5879211, 0.5880393, 0.5885903, 0.5861724, 0.5860248, 
    0.5838185, 0.5857811, 0.5866191, 0.5887516, 0.5900171, 0.5912229, 
    0.5938833, 0.5968704, 0.6010756, 0.6041175, 0.6061666, 0.6049091, 
    0.6060191, 0.6047784, 0.6041979, 0.6106832, 0.6070316, 0.6125202, 
    0.6122149, 0.6097252, 0.6122493, 0.5881223, 0.5874423, 0.585088, 
    0.5869296, 0.5835787, 0.585452, 0.5865321, 0.590719, 0.591643, 0.5925015, 
    0.5942009, 0.5963899, 0.600252, 0.6036355, 0.6067434, 0.606515, 
    0.6065955, 0.6072922, 0.6055682, 0.6075758, 0.6079137, 0.607031, 
    0.612174, 0.6106994, 0.6122084, 0.6112477, 0.5876632, 0.5888084, 
    0.5881893, 0.5893542, 0.5885333, 0.592193, 0.593295, 0.598482, 0.5963469, 
    0.5997487, 0.5966913, 0.5972319, 0.5998606, 0.596856, 0.6034486, 
    0.5989705, 0.6073194, 0.6028146, 0.607603, 0.6067299, 0.6081761, 
    0.6094749, 0.6111134, 0.614151, 0.6134459, 0.6159967, 0.59052, 0.5920138, 
    0.5918819, 0.5934491, 0.5946111, 0.5971382, 0.6012169, 0.5996793, 
    0.6025052, 0.6030745, 0.5987824, 0.6014137, 0.5930157, 0.5943638, 
    0.5935606, 0.5906379, 0.6000335, 0.5951911, 0.6041679, 0.6015183, 
    0.6092895, 0.6054103, 0.6130582, 0.616364, 0.6194943, 0.6231793, 
    0.5928306, 0.5918136, 0.5936357, 0.5961673, 0.5985264, 0.6016796, 
    0.6020032, 0.6025964, 0.604136, 0.6054341, 0.6027843, 0.60576, 0.5946774, 
    0.6004559, 0.5914299, 0.5941321, 0.5960177, 0.5951895, 0.5995038, 
    0.6005259, 0.6047001, 0.6025379, 0.6155463, 0.60975, 0.6260031, 
    0.6214069, 0.5914588, 0.592827, 0.5976165, 0.5953323, 0.6018906, 
    0.6035177, 0.604844, 0.6065448, 0.6067286, 0.6077392, 0.6060841, 
    0.6076736, 0.6016863, 0.6043533, 0.5970665, 0.5988309, 0.5980185, 
    0.5971288, 0.5998793, 0.6028261, 0.6028888, 0.6038374, 0.6065205, 
    0.6019173, 0.6163, 0.6073706, 0.5943229, 0.596976, 0.5973556, 0.5963256, 
    0.6033544, 0.6007968, 0.6077145, 0.6058357, 0.6089177, 0.6073838, 
    0.6071586, 0.6051962, 0.6039783, 0.6009138, 0.5984336, 0.5964749, 
    0.5969296, 0.5990835, 0.6030067, 0.6067454, 0.6059241, 0.6086828, 
    0.6014124, 0.6044487, 0.6032732, 0.6063439, 0.5996386, 0.6053442, 
    0.5981902, 0.5988135, 0.6007462, 0.6046556, 0.6055239, 0.6064534, 
    0.6058796, 0.6031066, 0.6026536, 0.600699, 0.6001608, 0.5986778, 
    0.5974532, 0.598572, 0.5997495, 0.6031076, 0.6061528, 0.6094934, 
    0.6103142, 0.6142529, 0.6110448, 0.6163503, 0.6118369, 0.6196756, 
    0.6056762, 0.611704, 0.6008341, 0.6019941, 0.6040993, 0.6089594, 
    0.6063294, 0.6094063, 0.6026358, 0.5991582, 0.5982617, 0.5965938, 
    0.5982998, 0.5981609, 0.5997981, 0.5992714, 0.6032195, 0.601095, 
    0.6071531, 0.6093818, 0.6157289, 0.6196603, 0.6236942, 0.6254861, 
    0.6260328, 0.6262615,
  0.662225, 0.6677868, 0.6666974, 0.6712427, 0.6687127, 0.6717014, 0.6633441, 
    0.6680099, 0.665023, 0.6627212, 0.680266, 0.671447, 0.6897113, 0.683875, 
    0.6987641, 0.6887957, 0.7008164, 0.698471, 0.7055875, 0.7035305, 
    0.7128335, 0.706542, 0.7177785, 0.7113178, 0.712319, 0.7063369, 
    0.6732004, 0.6791539, 0.6728516, 0.6736922, 0.6733146, 0.6687649, 
    0.6664983, 0.6618037, 0.6626505, 0.6661009, 0.674071, 0.6713414, 
    0.6782679, 0.6781096, 0.6860121, 0.6824228, 0.6960331, 0.6920994, 
    0.703616, 0.700676, 0.7034774, 0.7026249, 0.7034885, 0.6991888, 
    0.7010232, 0.6972683, 0.6830918, 0.6871873, 0.6751373, 0.6681207, 
    0.6635474, 0.6603436, 0.6607946, 0.6616561, 0.6661212, 0.6703797, 
    0.673666, 0.6758847, 0.6780869, 0.6848563, 0.6885019, 0.6968353, 
    0.695313, 0.6978962, 0.7003852, 0.704614, 0.7039136, 0.7057922, 
    0.6978274, 0.7030962, 0.6944495, 0.6967888, 0.6786906, 0.6720753, 
    0.6693089, 0.6669066, 0.6611418, 0.6651112, 0.6635403, 0.6672907, 
    0.6696983, 0.668505, 0.6759456, 0.673031, 0.6887194, 0.6818594, 
    0.7000937, 0.6956248, 0.7011753, 0.6983294, 0.7032232, 0.6988151, 
    0.7064945, 0.7081947, 0.7070318, 0.7115247, 0.6985728, 0.7034776, 
    0.6684718, 0.6686661, 0.6695726, 0.6656078, 0.6653668, 0.6617806, 
    0.6649694, 0.6663377, 0.6698383, 0.6719286, 0.6739291, 0.6783752, 
    0.6834211, 0.6906249, 0.6959124, 0.6995118, 0.6972992, 0.6992517, 
    0.6970699, 0.696053, 0.7075566, 0.7010404, 0.7108741, 0.7103208, 
    0.7058372, 0.7103831, 0.6688025, 0.6676857, 0.6638407, 0.6668457, 
    0.6613926, 0.6644331, 0.6661955, 0.6730921, 0.6746283, 0.6760604, 
    0.6789089, 0.6826055, 0.6892046, 0.6950702, 0.7005305, 0.7001269, 
    0.700269, 0.7015022, 0.6984574, 0.7020051, 0.7026052, 0.7010394, 
    0.7102469, 0.7075857, 0.7103091, 0.7085731, 0.6680483, 0.6699319, 
    0.6689126, 0.6708323, 0.6694788, 0.6755452, 0.6773883, 0.6861677, 
    0.6825324, 0.6883389, 0.6831169, 0.6840355, 0.6885312, 0.6833965, 
    0.6947441, 0.6870037, 0.7015502, 0.6936396, 0.7020534, 0.7005067, 
    0.7030718, 0.7053891, 0.708331, 0.7138419, 0.7125561, 0.7172271, 
    0.6727619, 0.6752464, 0.6750264, 0.6776465, 0.6795993, 0.6838762, 
    0.690869, 0.6882196, 0.6931018, 0.694092, 0.6866816, 0.6912094, 
    0.6769204, 0.679183, 0.6778335, 0.6729574, 0.6888286, 0.6805772, 
    0.6960006, 0.6913904, 0.7050576, 0.6981798, 0.7118508, 0.7179043, 
    0.7237218, 0.7306814, 0.6766106, 0.6749126, 0.6779595, 0.6822281, 
    0.6862437, 0.6916696, 0.6922303, 0.6932602, 0.6959448, 0.6982216, 
    0.6935871, 0.6987951, 0.679711, 0.6895557, 0.6742734, 0.6787932, 
    0.6819746, 0.6805744, 0.6879182, 0.6896763, 0.6969326, 0.6931586, 
    0.7163985, 0.7058816, 0.7360994, 0.7273186, 0.6743217, 0.6766046, 
    0.6846904, 0.6808155, 0.6920352, 0.6948647, 0.697185, 0.7001794, 
    0.7005042, 0.7022953, 0.6993663, 0.7021788, 0.6916813, 0.6963251, 
    0.6837544, 0.6867647, 0.6853759, 0.6838603, 0.6885634, 0.6936595, 
    0.6937687, 0.6954227, 0.7001365, 0.6920815, 0.7177864, 0.701641, 
    0.6791142, 0.6836005, 0.6842462, 0.6824965, 0.6945798, 0.6901435, 
    0.7022514, 0.6989284, 0.7043933, 0.7016647, 0.7012655, 0.6978033, 
    0.6956689, 0.6903456, 0.6860849, 0.6827495, 0.6835217, 0.6871973, 
    0.693974, 0.700534, 0.6990843, 0.7039743, 0.6912071, 0.6964921, 
    0.6944382, 0.6998247, 0.6881497, 0.6980636, 0.6856692, 0.6867349, 
    0.6900561, 0.6968546, 0.6983795, 0.700018, 0.6990057, 0.694148, 
    0.6933596, 0.6899748, 0.6890475, 0.6865025, 0.6844124, 0.6863216, 
    0.6883402, 0.6941498, 0.6994875, 0.7054223, 0.7068934, 0.7140279, 
    0.7082076, 0.7178791, 0.709637, 0.7240613, 0.6986476, 0.7093968, 
    0.690208, 0.6922146, 0.6958805, 0.7044677, 0.6997991, 0.7052664, 
    0.6933287, 0.6873253, 0.6857911, 0.6829513, 0.6858563, 0.6856189, 
    0.6884237, 0.6875194, 0.6943446, 0.6906585, 0.7012556, 0.7052225, 
    0.7167342, 0.7240328, 0.7316638, 0.7351018, 0.7361567, 0.736599,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01193812, 0.01193812, 0.01193812, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01893771, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01193812, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 0.01193812, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 0.01193812, 
    0.01193812, 0.01193812 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.353658e-11, 3.368474e-11, 3.365585e-11, 3.377543e-11, 3.370904e-11, 
    3.37873e-11, 3.356643e-11, 3.369039e-11, 3.36112e-11, 3.354962e-11, 
    3.400744e-11, 3.378049e-11, 3.424349e-11, 3.409844e-11, 3.446284e-11, 
    3.422082e-11, 3.451165e-11, 3.445576e-11, 3.462384e-11, 3.457562e-11, 
    3.479075e-11, 3.464599e-11, 3.490232e-11, 3.47561e-11, 3.477893e-11, 
    3.464105e-11, 3.382638e-11, 3.397943e-11, 3.381725e-11, 3.383907e-11, 
    3.382924e-11, 3.371027e-11, 3.365036e-11, 3.352495e-11, 3.354766e-11, 
    3.363974e-11, 3.384863e-11, 3.377762e-11, 3.395646e-11, 3.395243e-11, 
    3.415173e-11, 3.406181e-11, 3.439721e-11, 3.430176e-11, 3.457759e-11, 
    3.450812e-11, 3.457426e-11, 3.455414e-11, 3.457442e-11, 3.447263e-11, 
    3.451616e-11, 3.442662e-11, 3.407906e-11, 3.41813e-11, 3.387637e-11, 
    3.369325e-11, 3.357173e-11, 3.348559e-11, 3.349769e-11, 3.352092e-11, 
    3.364021e-11, 3.375245e-11, 3.383806e-11, 3.389531e-11, 3.395175e-11, 
    3.412284e-11, 3.421341e-11, 3.441643e-11, 3.437975e-11, 3.444182e-11, 
    3.450117e-11, 3.460084e-11, 3.458441e-11, 3.462831e-11, 3.444e-11, 
    3.45651e-11, 3.435858e-11, 3.441502e-11, 3.396745e-11, 3.379692e-11, 
    3.37245e-11, 3.366109e-11, 3.350703e-11, 3.361338e-11, 3.357141e-11, 
    3.367113e-11, 3.373454e-11, 3.370312e-11, 3.389684e-11, 3.382144e-11, 
    3.421873e-11, 3.404748e-11, 3.449429e-11, 3.438719e-11, 3.451986e-11, 
    3.445214e-11, 3.456813e-11, 3.446367e-11, 3.46446e-11, 3.468404e-11, 
    3.465701e-11, 3.476057e-11, 3.445767e-11, 3.457391e-11, 3.370244e-11, 
    3.370756e-11, 3.373136e-11, 3.362654e-11, 3.362012e-11, 3.352412e-11, 
    3.360945e-11, 3.364582e-11, 3.373813e-11, 3.379273e-11, 3.384466e-11, 
    3.3959e-11, 3.408673e-11, 3.426552e-11, 3.43941e-11, 3.44803e-11, 
    3.442739e-11, 3.447403e-11, 3.442181e-11, 3.43973e-11, 3.466916e-11, 
    3.451643e-11, 3.474557e-11, 3.473289e-11, 3.462908e-11, 3.473422e-11, 
    3.371109e-11, 3.368159e-11, 3.35794e-11, 3.36593e-11, 3.351361e-11, 
    3.359513e-11, 3.364197e-11, 3.382297e-11, 3.386273e-11, 3.389965e-11, 
    3.397255e-11, 3.406615e-11, 3.423056e-11, 3.437368e-11, 3.450449e-11, 
    3.449484e-11, 3.449821e-11, 3.452739e-11, 3.445496e-11, 3.453921e-11, 
    3.455332e-11, 3.451632e-11, 3.473109e-11, 3.466969e-11, 3.473248e-11, 
    3.469244e-11, 3.369112e-11, 3.374062e-11, 3.37138e-11, 3.376416e-11, 
    3.372861e-11, 3.388642e-11, 3.393372e-11, 3.415538e-11, 3.40643e-11, 
    3.42092e-11, 3.407895e-11, 3.410202e-11, 3.421382e-11, 3.408589e-11, 
    3.436567e-11, 3.417588e-11, 3.452849e-11, 3.433878e-11, 3.454031e-11, 
    3.450364e-11, 3.456423e-11, 3.461856e-11, 3.468684e-11, 3.481307e-11, 
    3.478375e-11, 3.488936e-11, 3.381447e-11, 3.387874e-11, 3.387306e-11, 
    3.394034e-11, 3.399011e-11, 3.409814e-11, 3.42715e-11, 3.420621e-11, 
    3.432594e-11, 3.435e-11, 3.416797e-11, 3.427967e-11, 3.392144e-11, 
    3.397921e-11, 3.394477e-11, 3.381902e-11, 3.422096e-11, 3.40145e-11, 
    3.439581e-11, 3.42838e-11, 3.461071e-11, 3.444803e-11, 3.476764e-11, 
    3.490448e-11, 3.503331e-11, 3.518397e-11, 3.391381e-11, 3.387004e-11, 
    3.394828e-11, 3.405665e-11, 3.415719e-11, 3.429105e-11, 3.43047e-11, 
    3.432974e-11, 3.439469e-11, 3.444937e-11, 3.433759e-11, 3.446298e-11, 
    3.399258e-11, 3.423888e-11, 3.385307e-11, 3.396915e-11, 3.404978e-11, 
    3.401438e-11, 3.419831e-11, 3.424165e-11, 3.441803e-11, 3.432683e-11, 
    3.48706e-11, 3.462978e-11, 3.529873e-11, 3.511154e-11, 3.385473e-11, 
    3.391352e-11, 3.41184e-11, 3.402087e-11, 3.429989e-11, 3.436865e-11, 
    3.442449e-11, 3.449602e-11, 3.450366e-11, 3.454606e-11, 3.447653e-11, 
    3.454325e-11, 3.429096e-11, 3.440362e-11, 3.409459e-11, 3.416969e-11, 
    3.41351e-11, 3.409712e-11, 3.421414e-11, 3.433896e-11, 3.434159e-11, 
    3.438155e-11, 3.449442e-11, 3.430038e-11, 3.490157e-11, 3.452998e-11, 
    3.397766e-11, 3.409104e-11, 3.41072e-11, 3.406325e-11, 3.436167e-11, 
    3.425346e-11, 3.454503e-11, 3.446611e-11, 3.45953e-11, 3.453108e-11, 
    3.452155e-11, 3.44391e-11, 3.438771e-11, 3.425815e-11, 3.415271e-11, 
    3.406922e-11, 3.408855e-11, 3.41803e-11, 3.43465e-11, 3.450394e-11, 
    3.446939e-11, 3.458504e-11, 3.427893e-11, 3.44072e-11, 3.435755e-11, 
    3.448688e-11, 3.420434e-11, 3.444553e-11, 3.414271e-11, 3.416918e-11, 
    3.425121e-11, 3.441643e-11, 3.445293e-11, 3.4492e-11, 3.446782e-11, 
    3.435098e-11, 3.433179e-11, 3.424899e-11, 3.42261e-11, 3.416309e-11, 
    3.411086e-11, 3.415852e-11, 3.42085e-11, 3.435075e-11, 3.447898e-11, 
    3.46189e-11, 3.465316e-11, 3.481683e-11, 3.468353e-11, 3.490347e-11, 
    3.47164e-11, 3.504027e-11, 3.445941e-11, 3.471161e-11, 3.425495e-11, 
    3.430404e-11, 3.439291e-11, 3.459695e-11, 3.448669e-11, 3.46156e-11, 
    3.433102e-11, 3.418352e-11, 3.414535e-11, 3.407424e-11, 3.414691e-11, 
    3.4141e-11, 3.421059e-11, 3.418815e-11, 3.435538e-11, 3.426551e-11, 
    3.452085e-11, 3.461417e-11, 3.487789e-11, 3.503972e-11, 3.520463e-11, 
    3.527743e-11, 3.52996e-11, 3.530884e-11,
  1.907281e-11, 1.921687e-11, 1.918883e-11, 1.930526e-11, 1.924065e-11, 
    1.931692e-11, 1.910199e-11, 1.92226e-11, 1.914557e-11, 1.908576e-11, 
    1.953192e-11, 1.931046e-11, 1.976297e-11, 1.9621e-11, 1.997833e-11, 
    1.974085e-11, 2.002633e-11, 1.997147e-11, 2.013679e-11, 2.008938e-11, 
    2.030135e-11, 2.015868e-11, 2.041155e-11, 2.026725e-11, 2.02898e-11, 
    2.015398e-11, 1.935496e-11, 1.95043e-11, 1.934612e-11, 1.936739e-11, 
    1.935785e-11, 1.924198e-11, 1.918368e-11, 1.906182e-11, 1.908392e-11, 
    1.917344e-11, 1.937695e-11, 1.930778e-11, 1.948229e-11, 1.947835e-11, 
    1.967328e-11, 1.95853e-11, 1.9914e-11, 1.982038e-11, 2.009135e-11, 
    2.002308e-11, 2.008814e-11, 2.006841e-11, 2.00884e-11, 1.99883e-11, 
    2.003117e-11, 1.994317e-11, 1.960177e-11, 1.970188e-11, 1.940384e-11, 
    1.922542e-11, 1.910727e-11, 1.902358e-11, 1.903541e-11, 1.905795e-11, 
    1.917396e-11, 1.928328e-11, 1.936674e-11, 1.942264e-11, 1.947778e-11, 
    1.964501e-11, 1.973375e-11, 1.993294e-11, 1.989695e-11, 1.995795e-11, 
    2.001629e-11, 2.011438e-11, 2.009823e-11, 2.014148e-11, 1.995634e-11, 
    2.007932e-11, 1.987645e-11, 1.993186e-11, 1.949276e-11, 1.932644e-11, 
    1.925589e-11, 1.919422e-11, 1.90445e-11, 1.914785e-11, 1.910708e-11, 
    1.920412e-11, 1.926588e-11, 1.923533e-11, 1.942417e-11, 1.935067e-11, 
    1.973901e-11, 1.957139e-11, 2.000949e-11, 1.990433e-11, 2.003472e-11, 
    1.996815e-11, 2.008226e-11, 1.997955e-11, 2.015759e-11, 2.019643e-11, 
    2.016988e-11, 2.027193e-11, 1.997386e-11, 2.008814e-11, 1.923447e-11, 
    1.923945e-11, 1.926267e-11, 1.91607e-11, 1.915447e-11, 1.906121e-11, 
    1.914418e-11, 1.917955e-11, 1.926946e-11, 1.932271e-11, 1.937338e-11, 
    1.948496e-11, 1.960985e-11, 1.978498e-11, 1.991114e-11, 1.999588e-11, 
    1.99439e-11, 1.998979e-11, 1.99385e-11, 1.991448e-11, 2.018187e-11, 
    2.003157e-11, 2.025724e-11, 2.024473e-11, 2.014251e-11, 2.024614e-11, 
    1.924295e-11, 1.921429e-11, 1.91149e-11, 1.919266e-11, 1.905107e-11, 
    1.913028e-11, 1.917587e-11, 1.93522e-11, 1.939103e-11, 1.942705e-11, 
    1.949827e-11, 1.95898e-11, 1.975075e-11, 1.989118e-11, 2.001969e-11, 
    2.001026e-11, 2.001358e-11, 2.004233e-11, 1.997115e-11, 2.005402e-11, 
    2.006794e-11, 2.003155e-11, 2.024306e-11, 2.018255e-11, 2.024447e-11, 
    2.020506e-11, 1.92236e-11, 1.927185e-11, 1.924577e-11, 1.929482e-11, 
    1.926026e-11, 1.941409e-11, 1.94603e-11, 1.967706e-11, 1.9588e-11, 
    1.972981e-11, 1.960239e-11, 1.962494e-11, 1.973444e-11, 1.960927e-11, 
    1.988342e-11, 1.96974e-11, 2.004344e-11, 1.985713e-11, 2.005514e-11, 
    2.001913e-11, 2.007876e-11, 2.013222e-11, 2.019955e-11, 2.032398e-11, 
    2.029514e-11, 2.039936e-11, 1.934385e-11, 1.940658e-11, 1.940106e-11, 
    1.946678e-11, 1.951543e-11, 1.962104e-11, 1.979086e-11, 1.972694e-11, 
    1.984434e-11, 1.986794e-11, 1.96896e-11, 1.979903e-11, 1.944861e-11, 
    1.950506e-11, 1.947144e-11, 1.93488e-11, 1.974166e-11, 1.953968e-11, 
    1.991323e-11, 1.980338e-11, 2.012459e-11, 1.996461e-11, 2.027927e-11, 
    2.041432e-11, 2.054171e-11, 2.069093e-11, 1.944085e-11, 1.939819e-11, 
    1.94746e-11, 1.958049e-11, 1.967893e-11, 1.981008e-11, 1.982351e-11, 
    1.984812e-11, 1.991192e-11, 1.996561e-11, 1.98559e-11, 1.997908e-11, 
    1.951816e-11, 1.975923e-11, 1.938207e-11, 1.949536e-11, 1.957424e-11, 
    1.953963e-11, 1.971964e-11, 1.976215e-11, 1.993524e-11, 1.98457e-11, 
    2.038095e-11, 2.014351e-11, 2.08048e-11, 2.061925e-11, 1.93833e-11, 
    1.94407e-11, 1.964099e-11, 1.95456e-11, 1.981884e-11, 1.98863e-11, 
    1.994121e-11, 2.001148e-11, 2.001907e-11, 2.006075e-11, 1.999247e-11, 
    2.005806e-11, 1.981035e-11, 1.992091e-11, 1.961806e-11, 1.969161e-11, 
    1.965776e-11, 1.962066e-11, 1.973526e-11, 1.985763e-11, 1.986025e-11, 
    1.989954e-11, 2.001041e-11, 1.981995e-11, 2.041166e-11, 2.004549e-11, 
    1.950338e-11, 1.961425e-11, 1.963011e-11, 1.958712e-11, 1.987954e-11, 
    1.977341e-11, 2.005974e-11, 1.998221e-11, 2.01093e-11, 2.004611e-11, 
    2.003682e-11, 1.995578e-11, 1.990538e-11, 1.977827e-11, 1.967506e-11, 
    1.959336e-11, 1.961234e-11, 1.970213e-11, 1.986512e-11, 2.001976e-11, 
    1.998585e-11, 2.009963e-11, 1.979898e-11, 1.992485e-11, 1.987617e-11, 
    2.000319e-11, 1.972524e-11, 1.996183e-11, 1.966493e-11, 1.969089e-11, 
    1.97713e-11, 1.993339e-11, 1.996932e-11, 2.000771e-11, 1.998402e-11, 
    1.986927e-11, 1.985049e-11, 1.976935e-11, 1.974696e-11, 1.968524e-11, 
    1.963419e-11, 1.968083e-11, 1.972985e-11, 1.986932e-11, 1.99953e-11, 
    2.013298e-11, 2.016673e-11, 2.032811e-11, 2.01967e-11, 2.041371e-11, 
    2.022914e-11, 2.054901e-11, 1.997558e-11, 2.022374e-11, 1.977496e-11, 
    1.982314e-11, 1.991037e-11, 2.011099e-11, 2.00026e-11, 2.012938e-11, 
    1.984976e-11, 1.970523e-11, 1.96679e-11, 1.959832e-11, 1.966949e-11, 
    1.96637e-11, 1.973188e-11, 1.970996e-11, 1.987395e-11, 1.97858e-11, 
    2.003658e-11, 2.012838e-11, 2.038843e-11, 2.054843e-11, 2.071176e-11, 
    2.0784e-11, 2.080601e-11, 2.081521e-11,
  1.783539e-11, 1.799306e-11, 1.796236e-11, 1.808986e-11, 1.801909e-11, 
    1.810264e-11, 1.786731e-11, 1.799933e-11, 1.791501e-11, 1.784957e-11, 
    1.833837e-11, 1.809556e-11, 1.859205e-11, 1.843613e-11, 1.882885e-11, 
    1.856774e-11, 1.888168e-11, 1.88213e-11, 1.90033e-11, 1.895108e-11, 
    1.918465e-11, 1.902742e-11, 1.93062e-11, 1.914705e-11, 1.917191e-11, 
    1.902224e-11, 1.814432e-11, 1.830806e-11, 1.813463e-11, 1.815794e-11, 
    1.814748e-11, 1.802055e-11, 1.795672e-11, 1.782337e-11, 1.784755e-11, 
    1.794551e-11, 1.816843e-11, 1.809263e-11, 1.828392e-11, 1.827959e-11, 
    1.849353e-11, 1.839694e-11, 1.875808e-11, 1.865514e-11, 1.895326e-11, 
    1.88781e-11, 1.894973e-11, 1.8928e-11, 1.895001e-11, 1.883983e-11, 
    1.8887e-11, 1.879017e-11, 1.841501e-11, 1.852494e-11, 1.81979e-11, 
    1.800242e-11, 1.787309e-11, 1.778156e-11, 1.779449e-11, 1.781914e-11, 
    1.794608e-11, 1.806578e-11, 1.815723e-11, 1.821851e-11, 1.827897e-11, 
    1.846249e-11, 1.855994e-11, 1.877892e-11, 1.873933e-11, 1.880643e-11, 
    1.887063e-11, 1.897862e-11, 1.896083e-11, 1.900847e-11, 1.880466e-11, 
    1.894001e-11, 1.871679e-11, 1.877773e-11, 1.829541e-11, 1.811306e-11, 
    1.803578e-11, 1.796826e-11, 1.780443e-11, 1.79175e-11, 1.787289e-11, 
    1.79791e-11, 1.804672e-11, 1.801326e-11, 1.822018e-11, 1.813962e-11, 
    1.856573e-11, 1.838168e-11, 1.886314e-11, 1.874745e-11, 1.889091e-11, 
    1.881765e-11, 1.894325e-11, 1.88302e-11, 1.902621e-11, 1.9069e-11, 
    1.903976e-11, 1.915221e-11, 1.882394e-11, 1.894973e-11, 1.801233e-11, 
    1.801778e-11, 1.80432e-11, 1.793156e-11, 1.792474e-11, 1.782271e-11, 
    1.791349e-11, 1.79522e-11, 1.805065e-11, 1.810898e-11, 1.816451e-11, 
    1.828685e-11, 1.842389e-11, 1.861624e-11, 1.875494e-11, 1.884816e-11, 
    1.879098e-11, 1.884146e-11, 1.878503e-11, 1.875861e-11, 1.905296e-11, 
    1.888744e-11, 1.913602e-11, 1.912223e-11, 1.90096e-11, 1.912378e-11, 
    1.802161e-11, 1.799023e-11, 1.788144e-11, 1.796655e-11, 1.781161e-11, 
    1.789827e-11, 1.794817e-11, 1.81413e-11, 1.818385e-11, 1.822334e-11, 
    1.830144e-11, 1.840188e-11, 1.857863e-11, 1.873299e-11, 1.887437e-11, 
    1.8864e-11, 1.886765e-11, 1.889929e-11, 1.882096e-11, 1.891216e-11, 
    1.892748e-11, 1.888743e-11, 1.912038e-11, 1.905371e-11, 1.912194e-11, 
    1.907851e-11, 1.800043e-11, 1.805326e-11, 1.80247e-11, 1.807842e-11, 
    1.804057e-11, 1.820913e-11, 1.82598e-11, 1.849768e-11, 1.83999e-11, 
    1.855562e-11, 1.841569e-11, 1.844045e-11, 1.85607e-11, 1.842324e-11, 
    1.872446e-11, 1.852002e-11, 1.890052e-11, 1.869555e-11, 1.891339e-11, 
    1.887376e-11, 1.89394e-11, 1.899827e-11, 1.907244e-11, 1.92096e-11, 
    1.91778e-11, 1.929275e-11, 1.813215e-11, 1.82009e-11, 1.819485e-11, 
    1.826691e-11, 1.832027e-11, 1.843617e-11, 1.86227e-11, 1.855246e-11, 
    1.868149e-11, 1.870743e-11, 1.851145e-11, 1.863168e-11, 1.824698e-11, 
    1.83089e-11, 1.827202e-11, 1.813757e-11, 1.856863e-11, 1.834688e-11, 
    1.875724e-11, 1.863646e-11, 1.898987e-11, 1.881376e-11, 1.916031e-11, 
    1.930925e-11, 1.944987e-11, 1.961472e-11, 1.823847e-11, 1.819171e-11, 
    1.827548e-11, 1.839165e-11, 1.849973e-11, 1.864382e-11, 1.865859e-11, 
    1.868564e-11, 1.875579e-11, 1.881486e-11, 1.869419e-11, 1.882968e-11, 
    1.832326e-11, 1.858794e-11, 1.817403e-11, 1.829825e-11, 1.83848e-11, 
    1.834682e-11, 1.854444e-11, 1.859115e-11, 1.878145e-11, 1.868298e-11, 
    1.927244e-11, 1.901071e-11, 1.974063e-11, 1.953551e-11, 1.817537e-11, 
    1.823831e-11, 1.845806e-11, 1.835337e-11, 1.865345e-11, 1.872763e-11, 
    1.878802e-11, 1.886533e-11, 1.887369e-11, 1.891957e-11, 1.884441e-11, 
    1.89166e-11, 1.864412e-11, 1.876568e-11, 1.843289e-11, 1.851366e-11, 
    1.847649e-11, 1.843575e-11, 1.856161e-11, 1.869609e-11, 1.869897e-11, 
    1.874218e-11, 1.886416e-11, 1.865467e-11, 1.930632e-11, 1.890277e-11, 
    1.830705e-11, 1.842872e-11, 1.844613e-11, 1.839894e-11, 1.872019e-11, 
    1.860352e-11, 1.891845e-11, 1.883312e-11, 1.897302e-11, 1.890345e-11, 
    1.889322e-11, 1.880404e-11, 1.874861e-11, 1.860886e-11, 1.849548e-11, 
    1.840578e-11, 1.842662e-11, 1.852521e-11, 1.870433e-11, 1.887445e-11, 
    1.883713e-11, 1.896238e-11, 1.863163e-11, 1.877002e-11, 1.871648e-11, 
    1.885622e-11, 1.85506e-11, 1.88107e-11, 1.848435e-11, 1.851287e-11, 
    1.86012e-11, 1.877942e-11, 1.881895e-11, 1.886119e-11, 1.883512e-11, 
    1.870889e-11, 1.868824e-11, 1.859906e-11, 1.857446e-11, 1.850666e-11, 
    1.845061e-11, 1.850182e-11, 1.855566e-11, 1.870894e-11, 1.884753e-11, 
    1.89991e-11, 1.903628e-11, 1.921415e-11, 1.90693e-11, 1.930857e-11, 
    1.910505e-11, 1.945793e-11, 1.882583e-11, 1.909909e-11, 1.860523e-11, 
    1.865818e-11, 1.87541e-11, 1.897488e-11, 1.885556e-11, 1.899514e-11, 
    1.868744e-11, 1.852861e-11, 1.848762e-11, 1.841123e-11, 1.848937e-11, 
    1.848301e-11, 1.85579e-11, 1.853382e-11, 1.871404e-11, 1.861714e-11, 
    1.889296e-11, 1.899404e-11, 1.928069e-11, 1.945728e-11, 1.963774e-11, 
    1.971762e-11, 1.974196e-11, 1.975214e-11,
  1.829493e-11, 1.846855e-11, 1.843474e-11, 1.857523e-11, 1.849723e-11, 
    1.858931e-11, 1.833006e-11, 1.847546e-11, 1.838258e-11, 1.831052e-11, 
    1.884933e-11, 1.858151e-11, 1.912946e-11, 1.895722e-11, 1.939129e-11, 
    1.910261e-11, 1.944975e-11, 1.938293e-11, 1.958437e-11, 1.952656e-11, 
    1.97853e-11, 1.961108e-11, 1.992006e-11, 1.974363e-11, 1.977118e-11, 
    1.960534e-11, 1.863525e-11, 1.881588e-11, 1.862458e-11, 1.865028e-11, 
    1.863874e-11, 1.849884e-11, 1.842853e-11, 1.828169e-11, 1.830831e-11, 
    1.841618e-11, 1.866184e-11, 1.857827e-11, 1.878922e-11, 1.878445e-11, 
    1.902061e-11, 1.891396e-11, 1.9313e-11, 1.919918e-11, 1.952897e-11, 
    1.944578e-11, 1.952506e-11, 1.9501e-11, 1.952537e-11, 1.940343e-11, 
    1.945563e-11, 1.93485e-11, 1.893391e-11, 1.905531e-11, 1.869433e-11, 
    1.847888e-11, 1.833643e-11, 1.823567e-11, 1.82499e-11, 1.827704e-11, 
    1.841681e-11, 1.854868e-11, 1.864949e-11, 1.871706e-11, 1.878376e-11, 
    1.898635e-11, 1.909399e-11, 1.933606e-11, 1.929226e-11, 1.936648e-11, 
    1.943751e-11, 1.955705e-11, 1.953735e-11, 1.95901e-11, 1.936452e-11, 
    1.95143e-11, 1.926734e-11, 1.933474e-11, 1.880192e-11, 1.86008e-11, 
    1.851563e-11, 1.844123e-11, 1.826084e-11, 1.838533e-11, 1.833621e-11, 
    1.845317e-11, 1.852768e-11, 1.849081e-11, 1.871891e-11, 1.863007e-11, 
    1.910037e-11, 1.889711e-11, 1.942922e-11, 1.930125e-11, 1.945996e-11, 
    1.937889e-11, 1.951789e-11, 1.939277e-11, 1.960975e-11, 1.965715e-11, 
    1.962475e-11, 1.974934e-11, 1.938585e-11, 1.952506e-11, 1.848978e-11, 
    1.849579e-11, 1.85238e-11, 1.840081e-11, 1.83933e-11, 1.828096e-11, 
    1.838091e-11, 1.842355e-11, 1.8532e-11, 1.85963e-11, 1.865752e-11, 
    1.879246e-11, 1.894371e-11, 1.915619e-11, 1.930953e-11, 1.941265e-11, 
    1.934939e-11, 1.940523e-11, 1.934281e-11, 1.931358e-11, 1.963938e-11, 
    1.945612e-11, 1.973139e-11, 1.971611e-11, 1.959135e-11, 1.971784e-11, 
    1.850001e-11, 1.846543e-11, 1.834562e-11, 1.843935e-11, 1.826875e-11, 
    1.836415e-11, 1.841911e-11, 1.863193e-11, 1.867884e-11, 1.87224e-11, 
    1.880856e-11, 1.891941e-11, 1.911462e-11, 1.928525e-11, 1.944165e-11, 
    1.943017e-11, 1.943421e-11, 1.946923e-11, 1.938255e-11, 1.948347e-11, 
    1.950044e-11, 1.94561e-11, 1.971407e-11, 1.96402e-11, 1.971579e-11, 
    1.966768e-11, 1.847667e-11, 1.853488e-11, 1.850342e-11, 1.856261e-11, 
    1.85209e-11, 1.870673e-11, 1.876262e-11, 1.90252e-11, 1.891722e-11, 
    1.90892e-11, 1.893466e-11, 1.8962e-11, 1.909483e-11, 1.894299e-11, 
    1.927583e-11, 1.904988e-11, 1.947059e-11, 1.924387e-11, 1.948484e-11, 
    1.944097e-11, 1.951362e-11, 1.95788e-11, 1.966095e-11, 1.981295e-11, 
    1.97777e-11, 1.990514e-11, 1.862184e-11, 1.869765e-11, 1.869097e-11, 
    1.877045e-11, 1.882934e-11, 1.895727e-11, 1.916332e-11, 1.908571e-11, 
    1.92283e-11, 1.925699e-11, 1.90404e-11, 1.917325e-11, 1.874847e-11, 
    1.881679e-11, 1.87761e-11, 1.862781e-11, 1.910358e-11, 1.88587e-11, 
    1.931207e-11, 1.917853e-11, 1.95695e-11, 1.93746e-11, 1.975831e-11, 
    1.992345e-11, 2.007945e-11, 2.026251e-11, 1.873909e-11, 1.86875e-11, 
    1.877991e-11, 1.890813e-11, 1.902746e-11, 1.918666e-11, 1.920299e-11, 
    1.92329e-11, 1.931047e-11, 1.937581e-11, 1.924236e-11, 1.93922e-11, 
    1.883266e-11, 1.912491e-11, 1.866802e-11, 1.880505e-11, 1.890056e-11, 
    1.885863e-11, 1.907685e-11, 1.912846e-11, 1.933886e-11, 1.922995e-11, 
    1.988263e-11, 1.959259e-11, 2.040242e-11, 2.017453e-11, 1.86695e-11, 
    1.873891e-11, 1.898145e-11, 1.886586e-11, 1.919731e-11, 1.927932e-11, 
    1.934611e-11, 1.943166e-11, 1.94409e-11, 1.949168e-11, 1.94085e-11, 
    1.948839e-11, 1.9187e-11, 1.932141e-11, 1.895365e-11, 1.904285e-11, 
    1.900179e-11, 1.89568e-11, 1.909581e-11, 1.924446e-11, 1.924764e-11, 
    1.929542e-11, 1.943038e-11, 1.919866e-11, 1.992022e-11, 1.947311e-11, 
    1.881474e-11, 1.894905e-11, 1.896826e-11, 1.891616e-11, 1.927109e-11, 
    1.914212e-11, 1.949044e-11, 1.939601e-11, 1.955085e-11, 1.947383e-11, 
    1.946251e-11, 1.936384e-11, 1.930252e-11, 1.914803e-11, 1.902276e-11, 
    1.892371e-11, 1.894672e-11, 1.90556e-11, 1.925357e-11, 1.944174e-11, 
    1.940044e-11, 1.953906e-11, 1.917319e-11, 1.93262e-11, 1.926699e-11, 
    1.942156e-11, 1.908365e-11, 1.937123e-11, 1.901047e-11, 1.904197e-11, 
    1.913957e-11, 1.933661e-11, 1.938032e-11, 1.942706e-11, 1.939822e-11, 
    1.92586e-11, 1.923578e-11, 1.913719e-11, 1.911002e-11, 1.903511e-11, 
    1.89732e-11, 1.902976e-11, 1.908925e-11, 1.925866e-11, 1.941195e-11, 
    1.957973e-11, 1.96209e-11, 1.981801e-11, 1.965748e-11, 1.992272e-11, 
    1.969712e-11, 2.008843e-11, 1.938795e-11, 1.96905e-11, 1.914401e-11, 
    1.920253e-11, 1.93086e-11, 1.955292e-11, 1.942083e-11, 1.957535e-11, 
    1.923488e-11, 1.905937e-11, 1.901408e-11, 1.892973e-11, 1.901601e-11, 
    1.900899e-11, 1.909171e-11, 1.906511e-11, 1.92643e-11, 1.915718e-11, 
    1.946223e-11, 1.957412e-11, 1.989177e-11, 2.00877e-11, 2.028808e-11, 
    2.037684e-11, 2.04039e-11, 2.041521e-11,
  1.973493e-11, 1.991887e-11, 1.988303e-11, 2.003195e-11, 1.994926e-11, 
    2.004689e-11, 1.977214e-11, 1.99262e-11, 1.982776e-11, 1.975144e-11, 
    2.032279e-11, 2.003861e-11, 2.062036e-11, 2.043734e-11, 2.089887e-11, 
    2.059183e-11, 2.096109e-11, 2.088996e-11, 2.110444e-11, 2.104287e-11, 
    2.131862e-11, 2.11329e-11, 2.146236e-11, 2.127417e-11, 2.130355e-11, 
    2.112679e-11, 2.00956e-11, 2.028729e-11, 2.008428e-11, 2.011154e-11, 
    2.009931e-11, 1.995097e-11, 1.987647e-11, 1.97209e-11, 1.974909e-11, 
    1.986337e-11, 2.012381e-11, 2.003517e-11, 2.025896e-11, 2.025389e-11, 
    2.050468e-11, 2.039138e-11, 2.081555e-11, 2.069448e-11, 2.104543e-11, 
    2.095685e-11, 2.104127e-11, 2.101565e-11, 2.10416e-11, 2.091178e-11, 
    2.096735e-11, 2.085331e-11, 2.041258e-11, 2.054155e-11, 2.015828e-11, 
    1.992983e-11, 1.977888e-11, 1.967217e-11, 1.968724e-11, 1.971598e-11, 
    1.986404e-11, 2.00038e-11, 2.01107e-11, 2.018239e-11, 2.025316e-11, 
    2.046829e-11, 2.058266e-11, 2.084008e-11, 2.079348e-11, 2.087246e-11, 
    2.094805e-11, 2.107534e-11, 2.105436e-11, 2.111055e-11, 2.087036e-11, 
    2.102982e-11, 2.076696e-11, 2.083867e-11, 2.027247e-11, 2.005906e-11, 
    1.996878e-11, 1.988992e-11, 1.969883e-11, 1.983068e-11, 1.977864e-11, 
    1.990256e-11, 1.998154e-11, 1.994245e-11, 2.018435e-11, 2.009011e-11, 
    2.058945e-11, 2.03735e-11, 2.093923e-11, 2.080304e-11, 2.097194e-11, 
    2.088565e-11, 2.103364e-11, 2.090043e-11, 2.113148e-11, 2.1182e-11, 
    2.114747e-11, 2.128025e-11, 2.089306e-11, 2.104127e-11, 1.994136e-11, 
    1.994773e-11, 1.997742e-11, 1.984709e-11, 1.983913e-11, 1.972013e-11, 
    1.982599e-11, 1.987117e-11, 1.998612e-11, 2.005429e-11, 2.011922e-11, 
    2.026239e-11, 2.042299e-11, 2.064877e-11, 2.081185e-11, 2.092158e-11, 
    2.085426e-11, 2.091369e-11, 2.084726e-11, 2.081616e-11, 2.116306e-11, 
    2.096787e-11, 2.126113e-11, 2.124484e-11, 2.111189e-11, 2.124667e-11, 
    1.99522e-11, 1.991555e-11, 1.978861e-11, 1.988791e-11, 1.970719e-11, 
    1.980824e-11, 1.986648e-11, 2.009209e-11, 2.014184e-11, 2.018805e-11, 
    2.027948e-11, 2.039717e-11, 2.060459e-11, 2.078603e-11, 2.095245e-11, 
    2.094023e-11, 2.094453e-11, 2.098182e-11, 2.088955e-11, 2.099699e-11, 
    2.101505e-11, 2.096784e-11, 2.124266e-11, 2.116393e-11, 2.124449e-11, 
    2.119321e-11, 1.992746e-11, 1.998917e-11, 1.995581e-11, 2.001858e-11, 
    1.997435e-11, 2.017144e-11, 2.023074e-11, 2.050956e-11, 2.039486e-11, 
    2.057757e-11, 2.041337e-11, 2.044241e-11, 2.058357e-11, 2.042222e-11, 
    2.077601e-11, 2.053579e-11, 2.098327e-11, 2.074202e-11, 2.099844e-11, 
    2.095173e-11, 2.102909e-11, 2.109852e-11, 2.118604e-11, 2.13481e-11, 
    2.13105e-11, 2.144643e-11, 2.008137e-11, 2.01618e-11, 2.01547e-11, 
    2.023904e-11, 2.030154e-11, 2.043738e-11, 2.065635e-11, 2.057385e-11, 
    2.072545e-11, 2.075596e-11, 2.05257e-11, 2.066691e-11, 2.021572e-11, 
    2.028823e-11, 2.024503e-11, 2.008772e-11, 2.059286e-11, 2.033272e-11, 
    2.081455e-11, 2.067252e-11, 2.108861e-11, 2.088109e-11, 2.128983e-11, 
    2.146598e-11, 2.16325e-11, 2.18281e-11, 2.020576e-11, 2.015102e-11, 
    2.024908e-11, 2.03852e-11, 2.051195e-11, 2.068117e-11, 2.069852e-11, 
    2.073033e-11, 2.081285e-11, 2.088237e-11, 2.074041e-11, 2.089982e-11, 
    2.030509e-11, 2.061552e-11, 2.013036e-11, 2.027577e-11, 2.037716e-11, 
    2.033264e-11, 2.056443e-11, 2.061928e-11, 2.084306e-11, 2.07272e-11, 
    2.142244e-11, 2.111321e-11, 2.197769e-11, 2.173408e-11, 2.013192e-11, 
    2.020556e-11, 2.046307e-11, 2.034032e-11, 2.069249e-11, 2.077972e-11, 
    2.085077e-11, 2.094182e-11, 2.095166e-11, 2.100572e-11, 2.091717e-11, 
    2.100222e-11, 2.068153e-11, 2.082449e-11, 2.043354e-11, 2.05283e-11, 
    2.048467e-11, 2.043688e-11, 2.058459e-11, 2.074264e-11, 2.074601e-11, 
    2.079684e-11, 2.09405e-11, 2.069392e-11, 2.146257e-11, 2.098599e-11, 
    2.028604e-11, 2.042866e-11, 2.044906e-11, 2.039372e-11, 2.077096e-11, 
    2.063382e-11, 2.10044e-11, 2.090387e-11, 2.106874e-11, 2.098672e-11, 
    2.097467e-11, 2.086963e-11, 2.080439e-11, 2.06401e-11, 2.050696e-11, 
    2.040174e-11, 2.042618e-11, 2.054186e-11, 2.075233e-11, 2.095256e-11, 
    2.09086e-11, 2.105618e-11, 2.066684e-11, 2.082959e-11, 2.076661e-11, 
    2.093107e-11, 2.057166e-11, 2.087754e-11, 2.04939e-11, 2.052737e-11, 
    2.06311e-11, 2.084067e-11, 2.088718e-11, 2.093693e-11, 2.090622e-11, 
    2.075768e-11, 2.07334e-11, 2.062857e-11, 2.059969e-11, 2.052008e-11, 
    2.045431e-11, 2.05144e-11, 2.057762e-11, 2.075774e-11, 2.092084e-11, 
    2.109951e-11, 2.114336e-11, 2.135351e-11, 2.118237e-11, 2.146524e-11, 
    2.122464e-11, 2.164212e-11, 2.089532e-11, 2.121756e-11, 2.063582e-11, 
    2.069804e-11, 2.081087e-11, 2.107096e-11, 2.09303e-11, 2.109484e-11, 
    2.073245e-11, 2.054587e-11, 2.049773e-11, 2.040813e-11, 2.049978e-11, 
    2.049232e-11, 2.058023e-11, 2.055195e-11, 2.076373e-11, 2.064982e-11, 
    2.097437e-11, 2.109354e-11, 2.143217e-11, 2.164132e-11, 2.185541e-11, 
    2.195033e-11, 2.197926e-11, 2.199137e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
